PK   '�X���@  H�     cirkitFile.json�]���8r�����_���e�.�nw����A���m�ܖO��#�y��L�)E�m˲d��س.�A�,������5_'���yU����^ϫ�䖩�����'۽O'���~���qr����/+��ӪZ�e�3�H^بd��d����E<�S.DZZ����݇鋻3�>ԙ�"O
GY�m$Y�#��4*+%�y���&��i�ZwI�h�ZwM랎�yl�$.xL�RDY��H�<ifR� ad32r�䆕����:�V�(�)�r����8�ei#3�:a��D�3"����xF�<#b�����֟����LX��*G�s��,"��ܨ2�e����]N�.'B��ˉ��D��1{��z>��̌r`�39I�Ȧ�E̘XX�2U4��ǌ=JlF{����Rc��0��Ǣ�04�̕��,(#������H$
�H�"���g"���J?t���̠3%�&H=T5�2���
�j�gF�c##'eI�M4���!B���0D�=<4Җ���s�e�@�HJ�DV�,҂W�y,���DR���(���\H���1|!���r�^��"�>�p��32e'�3��o�}��ZT5q�l�Oq�Cr�!�� \D.2�K���%�r��.��b����.xà���/�_�,�Y�0fi6&���b�C�.2Ea�<�y�0(�aP�à��P̔�Qޢ�,ǥ����.=v�&�,��M	��]�؝��`w�G ����
�p~��y�y�aS���Ŧ����#l:z�6�<�l�x^/ؔ��:¦o{.�Tl���QS���4�]S1:���EᢂpI�p�A��A��0��0�ea������0�`�,�Y�0(�aP���0(�aP�à��A1�b�<��E�S1:��F�bt.�N��\.���ѹ\���ѹ���"^Щ��E��N��\.j��ѹ\���ѹte�Tl�>7ۚ�ü�<�e�t�i^���jasW<@�VՅ�'�w�+��%��J1���G�et5>�3�O/Pj��e?22��P�i{��g�������c�ƙuJ�OYU#6�)�V�.ʁoRV724VrJHO:�v���Dk�T}/j�ŐC�!7���>&��p�t�>��4�u�g��� ����5@��t��Y��7>?��)ӗ!�7�%��h�TO}V���H@���sۺ�̗����s�\����ͼ�V.�5����t��(� ������?!������t&�
e��#��QPʨeT�2*F���Ҷ�Hb`�8�|�p�x-|ő$��
LN&��S��짦�{�(�E�� �G�]q챣��q	��5���H]�����UI�t��d�e�g@�c�.X�`��\�`�.a�p��e��Qϗ�f]��	�eN����N��Ѕ���5�����)_
=��>��k��a\��z�D�5?�^>o|��'�ۯ��XK�)�'e��yb橙'g������oy�����=���}�6��~cc�O����^�����c؎:`�߰>�h��q4�G0�t �l�xY����a�������K��2��] }�WЪڧ���uZ��Ԟ��YM�}�F0��g�]
ڧf���8Z���?�^�G+{�Z���]vhO���N+�=�<}��^�F��?��Ɵ[��-�7���C��\s�뵰];m�&~�$vM�I��i��5�Ӧdה�6�]�>mJwM�i��5#���!��-��־�_V�����������d>|mo���������bT��7�]�P3��	�j*x:c�I���߷�Mt^
�"2��`f�"2V�H�9��� r?���N'�6v�o���餪���n��lV����n�@w�虚J�>L��Y<c���$�Χ4�I՝�CS��bi?�&�F��{�ff�}�g���&n�,=Pr��1�ʴ�I��m[����U{-;���}ݹo�en8���kЀ6=��5���6$jf��aB�`�����L�\���z�kfJ�iY-
WO��O����On�'뿹&��L�'�S�q�T�7���%ZD*.�MK��k���բ�]���i�v�7v�9�y�hL�B�H;@t���2����w��"c&�/�����hR�!����b�4����.W���9S��2.A��A c`Ʃ���),BUJQnp�v���,~�@��.֮�$?<�E�s�K�Y�)DG�������Z�1KS~��l]Wͻ�[v�gt�Y�����R�2�Q��I
aAH1��E�v]i$�h��jbnb�Tp���Ǧ.�x��������~M��+�������-[�-u��gXt[�Wu�EQ��z��m� `rZ�n M3��E�b�2�
�;����	;�'�
+d1�(�5eQ.2x��)�*,-4HQ&C�:K ^��2/�"s���F�4�����(�`F�*����`��4�d�,���cP�yD�ۏ���ռ�Y�f�����z�����o`��/զ޶�x�GW��MS�ԛ�M����߷ퟖѢ���<��r�M�V�6�X|�2�J��[���c��4�N���>�x?��X*g`B���z��͛_�M1���l�f`$"���r�����!�A�'�ֲ�XU�\��w�*��B�(�	ئ�L�K��XQ[0�*w^���5��*&�b�Ⳙ'
ݝ��5tz�D���������uSϗ�����ٷN'�b�?��?���jwu7�9�B�Z?V��- �� �l֮�u��g��W��o�+��2y��Mi�fS���]��,o���8D��i�
��9��S�}���>LI��[�s *�l�	Q��Th� N1+5.nCm���pes��{P1�1��fpyF��#�_k��Ӈ�J�g��[G�-xg�8�:��2���!��Ln'IR^Z�n}^Vj����>�mճ���ẍ��κa��ʄ�FZ�����z�}���j㱺���~������{�o�v�m�y�]��⩁
LWR�_2̧��^-\�d.�O˃H��D�^�+��u��:��-���O�5����?��y`ٞX��6O��oޕ7o 6Y���Oۑ�HH9U�5��H��u�f65rf�~�2;�k�Te�X:��P�c��R�i�,j��� U�&�|g���aP�M��4aI�L�D�ԑ).M�0-#�@�g
G6O�AkVs��P5���B�6��^SL&;�����ہ,; �A|d|"�
KU�B/�!�O�>"�N1&����MY,�Ę)/�`8�J���B�إ�F�֠S۽&ƌͩ�6��C"��"v��k�y^��ʯ=�"nm\+��$�0����O�y�{&1���G7��i��Y�@J7?�:~��'l��7�����k�/��ݧ�����v���Uݦ��p��0h�n�ϗ����%��Ʋ8�
W�mY���/!E~'ݪ�/���yly}�������w�{��K�>�������mz���c�<�����)���˰OĤ��H�����~���:���t���U���P�x�j�M������kΦā�!�ڔ80�n����6俖
k~�)ǝ�����
�^e�Y�{�Tۍ�S*!f�	�c�@��j7u�ٕ�1��ח"A�;,���dW�� ��]	�6�: ��x��Ѓ#j#j�'�����F@Ѿ�	
ܡ5(pg��B4(�����̺3��hb�v{��qqJ�%����;O�Z�X`\!ݵ��M����I���Jo�� ��B_���;,�b��q�tD`�L&n�{Al{�넪=�t�*�+��������y	0��iǜD�j{�Ҕ�R�)Q��Myz����j�� S>-��;{D���`qJ5�H�Lgy8X�+pq�l�p�_���B�do[%G^Kut6�@���T�q�lu\>\�� {/�.N�5����0��F�:d�!�:�o�tL��`�
قY�E#}���D�G�B?���@���@Wd�Wb-�zQj{q���t�T������-����C��(`��C������E��o��S��CE5��=�����]��m\=����֣e�~���+~�ˍ]����6��=��GԪ����͟�:���)�ɷ�PK   �Xh��;�� �0 /   images/08e4a639-d7b6-43fd-85af-03d86c8bfac2.png̺gTS]�5�R�U��+�#Jo�;��j�j齆�{BGjh!"�$�� �};��s�1���<?NF�J�^�ּ�5����KM%��L�A ������R�
0�Ջ�~]��Wѻ
���|���l��v�~.t9�����
F޺nv�P+O[
�s;{Y[���yڧb��@�� ���|ӶQ~(�����v薼�v~�f9nIy�l�0��f̂$r?^���+��^�[�{�㣫W��T�Ҙ�>�9��"�1���4���7���s��k�X[�!�x���<:��ϴVo�b����U����A��/����ۋ���3����߃_�����`���%����-���%��iɂķ�#.�^	D!��"LY.������Z��3A1�ri����	�&1�`��w�g��{e
���kp�"���Bj��H���]ޗ������t��\2d�we*�1������ᨑ�y��ˆ���[?B�\��Oq����)��M�&��D��T#}����L{|�W2}�$k���z�\	�iKiT͈�V�o�k !��h����5ÈD�ǌ�q�ǕSË~lW�����p\�Ѕ�0d����Uq]���*�V��m9ޟ:�+C�^���'���E}�a��$��O��3�_,O{E�@	��\-QS�c��_=ur����4œ\�<��X)!?�-�V��dP��CQM4\�Ff�{� �=�xS��e\ӯ���WeJ˸�D���]�`��muݛ�H��?	�b�=�e�P��).�����@�����O�&bUz�Ie�T��_0�3���C�ÿ}R������>�H�Oo�q��t۵�X����_�9�����9�R| @J�]
���╸:o�|f��v�~��`��p� d@��6��#6���t��a�v���Ҿ\�����WpM��%W4-��F=}e���y�_��<#�/�~{S8Yu�@E	bS�~�@�zS��k�P:M���*���?p'�w��ɪ�8�7��6ڴ�E>����������I�6�3���){Tp4������ݏ@�"I˙T���,Y�Tr�K?4�?�A6ʰ^Ԅ��R��|_���;D�.*<o�h:�%^\9��[���_�J�,��P�'<���~�\���Nd��ێ؎��M-���~�5@W�E-=��{����:��[Z#�� P�疍�o��Cѡ�GpS,�#�k2.���)���+��Bc(��`f��اZ?"wV7����p�XV�����i�q17�6Q孳6T1&kaΝ9g���D�M�F��|�bd�Ht�4�%E�o�E�,lz��L��R�.F����NcQ�rὢ�3N��X��
I!�eQgM�p�nV�#/��}i=����(q;����2�v�f�i!r���Me�BN��M:���'~�Y?vK�8��֏�L���U����,P�E��"2�ʉ^`�꡹��X@��2uаɅ�S1�2µ�ª2Cr�He�R���"տ� >{�x7��a���KA���'��w�k��zJ��Ee���Q͞���T�T�)���t\z�W3���A�L�_�F��L�',��L���[�z�U��'��&�M�h�Dk��Ke�Tx?6��|�U�b�Љk���O�_�����)���D��9Gݍ*�T�Y���t?^<z�N�f_���Ċg���`\�&���X��B�l3qb����9��]bz6�]�Ij,���M6|����.���U�z¤��$_�����LLR�ìw�՗H���"����/�>�.H�������6sǦ(�'o;�O�+���Nz�Y(�>[�un��'U�BY"�q��p�w�v��ja��͠�����
6�H]"�����昜s�;r2�L+|��#���8��%�f/rP�=#�����i-�_1���b��(�2��9Dݦ!��|{<)6���Z���(�gn�n5@TBH�~�Ʀ�����l�H�Y�t*Lb�^%¶��x�6��ՓH.��Q9'��P�W�����[�)�xy�f[��G�\�F��Ĕ���k���ʨ�@���C׍A����X��Ĵ�x�ß�v+�I���i�Ϩ�����(G9Bh�Z���K�)M�2Ņخ�n�\���R���]?e`
�-�$���>k5���\�Ո��:��M܍&���9@hH8��.�_���%L
 j0�[k��9Tޏ�.>�혪m��+(5:j@i��R\��9i��^W�$�=�<t �~7��W�Z�E������Ȗ�:+���F	��ߨ���5�3E���'�|��%[&�%D�Q��b�S�ώ���Q�@^K�q^[$f���oSLN�ڴ���������`�%m���$Y����ھ��-H�f`�#h��Yr�����T���;�+	:�75P"���+3��Ϗ_�x��x�k�3�2�=�pY�z�,��m*�����B��O�U���G�_�t��溜Խ�B���|�X[�w���v���U9p<%t���m���(.�(�ƕ.Up9@([�L�B�ӈ{���dݯ`3-�=�hj�`��m�����%t3Vhfp0��&�N�IR�� �в�Kym!eϹ��
���w��~���ʧm���V�9:��}*�4|�q���-M��+�f �/�:?S�@�3b!����q��;�tWgsC􆳖n����cZ}�i�8<ީ��}2��q.��#�231n�(={7�;>"[ɢL�����~�Q?ro��e��y(ϛjQ�rM�S2�y��,�O�L^�܎\�����O��:?Y���5� ���.��%=�u�Dm�����*����#��K��k�����t'0N[��������X5X����ֽ��]
��[�J��w9UZ6AAC+k����̓��[uVJ�)�����\��p3��߆�v?��S�{-ߓ��X�|�≩e4�	?SĆ5�,n�ɭ4�"����P]��C��|��n>�,���v��2�gX^��8�$��7�oA��2�D �����+������������܍\
���l��.]��ۏ6DnV���[��4S�0]|�&�r)���	eLut�N ��S{�ػ����h�p�IG]��q��YWL�ݔ�MM|(��H���MSMl�oj_D}���om��J��|H������IW/�l�6�E�U��*��$��{WNZە��j���T,�2x��A.�S&�ɬ����qځ��g'v�cmG�U!go�\
��5�n?��P��;���,�.ۆ���5��]F�/P�]1Z��Vi>?��Z S��O}B��� i-`�*��=��D��<A;}���Ծ�7􂍛�z$�a�[2A�W)qR��o���o�ژ�>�w��Z�_ uf9aϗ�;���i�l��y�ok�����*I*�j��e&am�ė&+����dɨ���h�)o�E���ǌ��,r$`n�\*I��>��6��2~_=�DJ+Q&�-s"��Y�p��sװ���nP���l�_��Y�X|W��o`�%��1��+]EU��!��Z#.�2B
�R�"5���栽D�M*���]��g���r<ف:��ohO�DeȠN�D̞��p�d�u�4�|H�i�n��&��"Z�������=yfB�v�d�F�n����֞�>�gS��C��7|�C1�����Є}���"7v����4��Gk���v��.��.�b>[Yw$Qh�G��d�<����Ud���2f�(�@_���L�"�A��~�r�e���#w���^v��-99�t�ݚ)t5�{���C����b�$��������T�n)rI��Z��J<;���;��C��Z�]!eD�1��;�Mn'�Ƃ}��E�qEz�ż� Y��� |l���G��gVu�k_�. 
�="�u���������-g���6�T�E(�0�G���q�T��S"J�$G��4;-_�^��c�w�j/*���_�<9�3:4[ߡ�n>�3�
��h�Vx���:ɸ�H?�YDw� qs��Z��������gm��'\Z�>��a�[o ��3�Aa��Ȱ*�[^�c
���֛�M�"7��3����f�7��p�)�������߬���s鋅`1����'�~
�J\��b��p�����������Rd������>�)v���'���<��P�\���H��<�i�������ݩ��K�3��>d��t^�J�������g��S��ǘ�g�Y���:;��i�V-�S)4p*c�}bG�8j|hj*�f�8�a^Hk�� �k5�$��,�VKo?٣��d��[��,������w���_ۖ�6�$�y��E���o�^�������2t�1�Pf$ �y!���oL�Gs��WV����Gt�7ޘ��[�/��8k�s�����t�\���\D��Yi+H~ƚ���������l�������A�nL�W�X�KF\��2b�2���|��2W�t
�&=����-V��k�p��$!K�g=]��ŝ��:
�j�#D���쾏�T�SZ.i�Dmʶ���r��8C��j�Y���peWe��>��t�<�zXt"��[�����)Y|�?k7~ɸ�	�V���/���T*��v���e���~�$�ճgO�j�{��PMXlj"�fe���rZ
�����P��G@GI�+'c�#��#�:��N�u?�X��@�tW��H�i8?!m��%�5Z�S����Ӿ�ܹ5 @�zo\�6��E�t�=*�#@��{F��d����!�sg[�9X@�?�z��֍C����Ɉ3�h�6�t�-��ٍ��09(����H)7���&Y[�ǭ�r�6ֺ���T,��T��,ҸӾ,�"����:�G����s���__�x�Pj^��('��҂n����(/�>��Mm����ۺe]�>�S��=�8�ߚ�]Z��Ԥi�{n�06�8��c�>�:��x�!��9�3
#J�68�\��"��,�@_�i�1�"���J�o#°l��$�����8���l M��rp��+�9ĵ����N�~�'���=?�t��Ҵ�\ƈ�s7|���� �r�^�KFx7}:�P�`��wߵVBu���F�����(��	�J�}�#=���)�
��g����ĳ����ak��3a�}=�8m���:�q�Y��C�23A�����S�m} ��)N~��:��� ��P���lgM���5�͵�ퟹw6i��_^���|��-q�/N8���Uɣ��5CM�q�~�,x��G�/��~��p��܎�i�D#h#i#�i"��]�X��EP�q�@K�kl��`.6����o�[K֛9����Ǩ����9-�o�*\��כ��t��IE��B����$���� �i�ѭ�)7r�=�\?��ڂ>� w��Jø�W*����n_q��b[����DU96�c�8?Z�R������Hw�=.'l�d����W�Ù��秈����Meƈ�����[V�j_w^Mv$��6&��W���c���,���J�.�*�w�q��2�o�]�b�&tyG ��_��ѴtF������$֝���J�-�4�J�b�/k��^˵s���j�;�]��5�9{�y捩�Q׈�t��f�U��Fy#��8^�#��-3a��0#)L
���?v>�8��65:OD�_b����.�Q�����z��Tz �د�3������ 
�ODM�8��'1}Wn�_"+ѯ��l�m�.���q,�:�v�1gqu&M����௼ oݲ�(�J	jз��V���K;���Ew��c�3{Hʳ�K ������.cdwm͙r�x��ԥӭ4�﬐ϫ��l�G^��;x���s������AA�!�v�DS��i�'5��2���fX��+	��#*Ss�D(۪�4����+r"�s\i�8sT�cpp�U�=P	����l�ʉ��9��C�ޫ�����޳:%K6�23���#E�2R
j_�Ŗ�3���`E��q�%���^�!.�)�>Ǖ�O4t5��a�c�_�(�g���#��3�X��T�/d��N�JG&;p�����?���v�
�<,���F/�Ķ��	�=(�����Q$�:I�BQ
��\����ϘN���7�aM,c����@3�}�MQ��+�^�*��(����Ҽ��I���Cu��T�A���� ~>5�8�嶩l�9����=Q9����q�K�"l!4�qV�k��?��O� $�A }h��(���@t��-�-
 �\ ��y�����Lh�7�1���ˁX��oN(���)�f��<�A� ��N˘�ݚQ�,�н�:���Z:���Ceq�˾�k`�@6�K[f`�{r̸Mp��#o���g������q�j�O���lϝX�%4g�}o�p���o����7J?�_��u�Vl��m�l�����x�q��|~6�rjz�n����Ɲ^6N�)嚢w�ݯO��#&z����ͥ���"�w"���P�� ��WO��z9�+�[5�م�y�1��/,�f��a�iA��� C���h�,`1+Ĵ�ݙf�ۢSp�������x2�@�ɼ�Q�!�[��!!��\�[�������|<ňP�-w;�P3�D �q�����`��d�+p��ߦ��"��u��aI3�²�7H�D��9�Kp�i�J2Ȧ�{�)�h=���%�����A��#%Њ�;���Z|�\��U����bU�Ҩ��SD�ʶV� h�B 	(S���K|V9�T �V���qgv�����넓n9�@w�m���-�K�� �������á_�=f����L����9����#�r�=RB,��2?ms�2u�axf`��}���Oi��^'�ʢ��o�yZ����|R=��*��k>!}�ѻ���	��+�'v&}dE
��\R�((qR��e�DsKcA5d�����3ڃ'�ps�f�f��t �l4���r0E�}�)��^R�8~Ї���.��5'����� i�H��4�y����2�1�yM���b�O5t�_�� ���#�I�9Pݼ�OH�vV���^Ǔd�����pÀ��@0��~�:�H�@}�Qp�,*���,u+�|V_0�R9�-����Cckgu>7<�8{ZQ�ɫ�{Ӓt�v��H~
#�^��B&�fj�{&I�wr��wI����jv�O�����j[��kx�`�����r�u�-{L�af�*qV%�7h}�~�59�M���K�����͕� �F��F�_� GҐ]Pc��$hr���L$����Q*l��vO���9ť�4�S%��3�:��۫k��[T�G�s����&I�ݨ����]�4���� ���I�}n[��wK���(HG���f�P.���������G�k��iII����葁c��Pys6cj���?������ο��qk�NԥE��8�_��Y����V�ܝ�%��J��f�sz��"�8=��F���6�t�hפ:�T����%qEQ���s���0~y=�"-�w���Kt��޿ܡ���Q�Q?-%`ߣ!~ZMvN藖��d�{U�����_7*|�/�J<-5���PȆ�(�#]�����G�y'胛�#�`�Q�@b�;���;C��=ɫ�k��Ӛrce49��3E1���E��R��S��bb�|D�o�|Cz75���k�@ۈ���|�\�0���<�z��g�H��r�8z�J�))J<�&���9�j%H�$�\x�&�UA?FCS̬e�g�"�t�n��_�j��$M$a�8j6hsZ�օcr�i������@7�w���� B�����^�7���ih:H��'gaX���#J�2$>G�u���}o���~�tb��f����8m��4]5�Ĝ�nGP�,M�������s;=���޸�+u�$��5�P��E�c�%�e��9:�*�(������x�&O���b5v����6�����W�����;�ޮ��O�Z��S�L���������<Z@�[�P�|[����`����nf��~$�!��qV�Ty����p-����W	"zL�e=��b��ɑ��4�:����Bȸ��߻�5����-'�U�4w9�Ҟ��ڊ����ґ�j3�G�Vv|��a���v�Os��9ǿ�h�g��R����>\�!ZV�H&�wz���E!��r�Oy�_������R ��uU���}L3�]�	���]�6t��/#��]�_��������e�mw��{���xwI��ˆ�x�C8h�J��%��RG�Y�jP��Ψ�Ȳ6t����s�5�dS=QU"�ڒ���)�˳�fmf�j��~&b��
�ܯ0�L>-�v���z0v�&kB��X"��t ŚI1'����9�dq����dtn*�P���mDS$���de���B1	��D���$t� *���<,���梋xLa�B&w�$9��[~��k/�9��{�A�lm���F\�-�Gz�1���[P�V536��TU��Q�Q�	��xH-��\\�xv挻��9�~����ϴ������T���3��;��jg��	*�!��̎ƅ�>� ����p�����Ҩ8ύ�{*	��G����:�Z�4.�/�$�c���n����s^.s�C�o�I�8dI������,O~�:X#��gA�w:f�F,��B+�eQOxH%@jB��p�8z{D�7+%��FO��7���g�!*4��m��K��@_zY�4r�~I.��A��&K�0+)��&(�kJv�@���S�ȩ�ܪ={������V��V�|�]�u,k����f0�k;قc��ҷQ�"�P	5�c�q��B��J����˛���n̢�:���Y�)p���w�~��%�Ή�y��^��(^����Q?�{� ��ڹ�;�'�� ��
��
h���+ܿ	����N���J OAw��E
�=�C�5�7Cy�>n��'n,
�[�@�{�ج�@u�A�nfjS�B#�?CA��k���=�ga����Q�AN�x���8u6��RñD��Ӄ���j��)���$NշEt-�}���ܢt�D\K�#v�U7��<�]��V'�v[%�g(��J$S+�"�&4����7z��6�1��%t���&M�,,zNZ%����i]Sb�sT��e=ḱ�/:���m ��/4#�0U=�[�!�m"6I[�D6UIX�/����^+#�ve���z�6Z��y�4�$Ӎ�A�W��v��kX���s)��<-����@�����T����9E��J�r-�&z+�5�Q!��w�8иS��\�$�����ǿ�����P�K�X�F��ܨ pK�ǐ ÌI�'kn0�a1Ċ[G,k�^cP1�_�*�o�E	l�D�EL�>9�M�Y:��g���dW~��/����f��e)۰�J�<��*��7�+Z�N��Z�@�D�b��R�}t��2j�\��>�j��T�Î�kgV����V�[����dAp�I�a�p����~��B*p�-��M DJ��u �	t��|  �r+%��^=2�N]��[+���Hz��2��s9�f��ݢ��οA�4�����q>�va��LjC{��'�8��x\M���v�ĝ ����=Hl�V5��l8�6�
��JDs���b�����N#Sk��I#�&:,��d���ޕup�?����Q�Ll�����}����������*��Pz�v��<q��f�Ǔ���Y��F�0(4��3y��6;�k����]�`�Z��d�"�_g?\kAB���ԡ&��,qFG4���H)�+�$�o��-��%�ZM�xڑ�R���g�g�7Vn���{إ�J�.KQ���{��X�IW76���M%n���g�ꄔ����LS�N�N�cS�Qc���7F:�\��P>�uFR`ǄO+�N�6�����/�=xk��z���!��Y�
"�� ����gaA驫/>F�����r�gԟ[����$����&N�ɞLŹ5D6[)�YB�2�%7��<�vj]51�u�e+G������P��;��M�����a�$�.�0Rڴ�>e���9ʧ��9"q(��Y:������V��8�\�#>*=�x���"�Za�O7��ؘ㊁i�#�Szs�o�V�E�YH<�ͿR&���$��� To�����Z�o	�������j]6��ȉz3������n�(���#<k�d���J|��!��qFh��J��XsÍ6��tL�B�U}�x9�����~�v���� ��H-bsv����kq�E�M�YE��U��B
]֠�ڂEz~Aa���@�D�������B<}��\�^4�ɠ��Y�l*���)p|�TS��R���7����hߘ�ޒ�;�ՏҨ7�i�S��t����o�pA��^rlI.������%��p�|L?�$yq���S��Wy���JY���/!$�G&\��`��?����x�6��S*�K�	�%/��!�,����BȰ�~�#�c,�l��0��y��0���y�����g,K�"�eȔ�d��h״F��?�굡q�S�a�~f�On�]�������M	�V��b!��^b�3��U��&��3��8�a����5f�~kG��tS��-���A�Q<c�D�����ѸW��P�m��E9�����`���n;�u�-T�^\㡈ɏ�V~�uC�<�]��$̧0�m3G�#	�FO���ұwi�P��IAۚ���t*L��h�o�r3�-T�<�|���#�Љ��`�O}��z��|9�=��=T�-������h��q0b�7ᩆ ����ص��W���[��IB�ͦ&�.^�5B����k��S�=���Q�~�u��J��>?��	��a٬�s�¯�3�����P>$��8��|$�<}kܻ�[�4�?��<�oI\�I5�����D��=� %�v�s}��j��*�1����Bf"5�m���N���BPo��s����*��4�:;�*��\#�ˢ�<�y�ը�#��F�y/]���FP(��ĮP
��7]���דe��U	G�w�8'�4��G3kW�s��Xe2�c�d�:��)[�p�r���㊫��<�pY��a���ΰ&�8_�o�TƔh�����wo�����ު2�ґ �0FP[t�W&���Đ������i�\�;�o0B]��/7|�F_F�ϓ볭.�����ᖎc_¦<3��)� [v�'��l���eg�����?x��u�ߤ&��d;�B�2 6ӯ�\� ��Fb�L��G�n���	�IGk���^4X�p�\��Z��vx�j��tA3�RNQ:`�F�Ψ��dg���Ty���	�,�!�U��~�W�Е���#��k��.����9��]w��1~{ŏ�äl��{N�o]Wҕ%TW�<�/����y��@C·MC~�AG�(sp�xg4�����J�� _��|�jֲ�mm�����s�7�@��T�<	"e	���()	��~�n��"Æ�f�\O�Yb���n��,�rS�� '�~��%�A=�J��M��3�Cp�b��R�#?�`u���v��ڌַ�s�n�.
��e�`|I'ƀ�����ڌ����;޿Y�~�Zq���,���۬��p��W-cnh���yYJ�VG��t�F�Ғ���َ �DJ���v����Ӳ�e{u��Ce�X�Vi�']Y�/�Y9_��c�
4=5,qV�@��4'��\������˼��N�פ:�$n��pX�;K�6ו��>�c}�"���΢��\��M����A�3O�����`�D��5�s���S�w/���Χ���Q;�Ç�T�d5u�r�rx���HS�ׅ�ۚ٩|ݦD��[0�2i�WHձ4p�1�{���U�Ѳ�3U�ǁ0���v����a����1=P~2>=���:�6:y���E��ߏ�u$�H̾zJ�r>#l���n39�)ɑ��Yn,·r���V6���e��yc�62���Rz�l�`��Os����-�r�[�)��k%�'��(ȘW	�Q�7����ٔ�a��8nDУ�8������R�v����è���Zb�'5{�P]�q癒a�_����}|���HR�/��o[t��7�ni�ĺ<);,G�>e�Y��5C-�xT���p�� 9����i�o1�S�Yxx	"t����ih��UM:#��/%����ͧߋ<��� �}2�rk��ǣH3�lΆ���)o�J۔�=R��1v`�c�˝�yt�up�d��ʷ�L��ίT�ώI~|��<BP�iذ]]Hl�o�D3}�^��`�w9U��儦��滝E�ØZglc�3��7���&W5��,�r���xC�������矵1~���K^��7�j���"��`�y�7x#!�?Nf5^_Q+�6�n��h���ȯ�zB���_�-���8�}��lf|Z�e9Lt���(#�ş�4H�Ϣ���3���x�EΪ�_S�v��L��0ϯ�t�j�'v%�z�N)�
��OD�����U���.�������Eݟ9 ��	}�8?k����	ap�KC�2LG�⾭͛c��������} �?���<9�	*z��x�I`q,�yu�����W����4��F��5��#,:�h��$f��=��o��gCwWŎ��l�X�4�v�A�F����_N�+��6e�/������D�}0�/���aLR�%|�3ջ`x�~�"S��qP�u%��đG��?darZ�Ń���:�;ˌ6���v�S�ڼ��5jG���n���g�harg���.�?/]?`}�m�3�I'Q���+Ð�e(��ʺ�d����T*|�z��2+��5l�fLr(Rzc�n�5�ݾ�R�/�[1)'qػ�������9�ã�-?�E�cp�y�\J�<g��( o9��*/4N'���y�����;�u�u���x|�k�!�=�3F*I
�w���2�Y�g����<a�B R���v�����wN^��n*^|�γ8Q�>�"m��/����/�8-u��P��4�-Hq�\��|��uA^�d����xy��B끂�}�RԆ�u�+C}�F�sW�����y�f��Gn��d���-q�����S��م,��L��-��&9����v��x�뽖��ĉ�>��Ӑ
N�u�v�IF.����jM�΄�zi��շ�.Lۧ�Q���,6ON{�56��q-��hWi~��%�Ylvpj8���$z�fr���s!P��c����Y=���^N��yU��ò7ŏҚ����L�)��k�+�����C
������*��%Ɩ��OY���KiU�-�x�kY*꣋��h҇��R<a~�>���&��j�{��t�^���!�c�Ɖ�u%��/բMQ�QW���I�[Lsf�-o}n3����o�P��=y .��6��y<�y$�A�����r`�y;|�&V����}IB��ց��e� ��/0S(X�^��g�q�OF�H�WP��c�ß�� ��
Ywg�g\�R�9��}�ו��A3UO�w%�dT ��?r#&�̆�\Ӂ��:�3a����m�����'��s��S�<dq���Wa&��N�
�W��~�ooTu����9������\����5�PÜ�[��W�����i����8`��K��0�MN�h�[4ڼ��b��}�=��lٓ�y�E���*�9J蹰�VՕ������23-����T*JF�;��B�����h�cT�NF]���M�M&gu2�¿����?nI��.�@�'>f�ӧa�u
���W񔜮h����V�����G�8>��5/���ϋ�;K=��D3��E}���2�2����W�_��� <F�y��!�CiF�S�>,��[�Q�(���k�p�Ѭ����>G:&?�����6��
n&
I��a���#�j0�<:��%���(��Rm$\{��|�v^d����o]���QiN.��a9��bi3�r����m��'X#75)"�.����_�N�9/H��:�Ap�P��\�B�d�X��?b�}��9�^z'�ҠJ�.J+�s�c�6��~O��Sg��e�)kp��ꇎ�-Y��=�z�5X�Y��X�rM�n�#T�:��X� �d�<5Yh���C�Ѩ�tX���O�֬qst�UX�)6@� O�-�+'������}��Q����0��EO���&�M&,����8j�U=��^�	D6�������(x��zN��U�r�͝�=�pނ��� ��*�*�8�?�}n쿔ε��,B|B3N�e8�)�TS�� Ƅj���=�{	�h�n8Y��e��`��V� ����u�. �M:F(O����x���<�L?�G��t�������5�핇��,#�*d�@{`�<Sp��T8^�Lm9�6x�\&r#f�@��Zp�k@|�{]�?*�%ο?�^�4�lW�'i�^�����U�\�a�O���6ØI#�s���E�-+��ק�\4�ځTT�r �Գ�PT3����l�cգǸ��n��>��_���,�G�]r=�*�yi����C���i�L[҇��t�J�����];빓�7�7�J�р��W�],NZ�͠��S��6���'R����m�t������V3�$�UP��U7��D6�R.�ק��<�D<&;��<.�d�J��n
'⬣=�%|Nˆ�|W.�!M����W=����V�=���^�'��T�+���5�\��n�����ȫ>Nf�1A�t��J⺲i2{]�:o�/{?ĸkT��(�q���8��+���]���9� �����u?+t%�x6�)����u�`�6�p413�^�n�b'w���'�r��h<3� �����s�8�]��R�Nk�=nn*v�Z��K�Ycc���mg��5'���ߢ���CϬm[��@IJA��:��p�'��Y헉���ޜW������&��8�iX ����q^ih?oiO�n��(��T����Hݻ�O�Ý.�"�7�n��_�|����p�X!�lwj��E>�k�X��L��t�/W�3���m�y�ؔ�t���)S��r�H��~�Q���i�F>=�)c����&ᥜ�#������#��S�	���m��[1VL�������WW�T�񚴨k��U���hb��`|'u�!L�x���J7SB}~-�h1I�������}�g_��=gI
R2�7�]r�C����֦{��M���O�f�_�7����N4��<�p�U�ě�;Τ;�-W+��<H�u�1z酆�7�������2�9�R/zN�f�DsE/-�UJ�b�f�L��f'�F���x��pdI��	]���yci�&�6L����l��C��#�]Ҷ�ń�1�R
#6��Fw���.���j��ޤ}�l��Yp�)]p�5�eSu�����`V�K�%�4��eT�����E���^dB[ߑ�Y�����<`Q��&:�p�@�
����.�����_`2�9,��<ߗ�`�V75�=�PԞV�_���e����JBb����w�� �B���8`3���W�7m�Vq�~���,@� N�Rײ6���ո��zS��e2*!K⶘=��C�.�ZE�R+���U`��ş�3��e �(*Z�����eυ�&?��e�i%�[Z��#��͞ɔ.y��R��j�yhX�6�a�{u����?�����Y�)����o]ux��7��9H�v��&F�^*�s���,��d*�����	��˵�$�w~�F�K{xQ����,��,E7C|�$��@�d���_u��k;�n�*�Q�Y�[���;�1�Niul�V2f��L���8����5�=}���?��*N+
�C�Ŋ�$�r�������'�[�&��y6�T�Ըֳ�25�^U������/�r�kW#���K�>6a��Uk����PDL:4��P-��W���δk�ז����ڊ�&,C��VT@0h�?���y�b�e���v&%���j�A��.܇7�.�r4���6�!8��j��!RԢ�;|�q�5�]a���%�u]�疵9��ZF��"�����T��CZ����3{V���;q>��g��s�0���3K~�kO���U��rt�a*���a��K�mq�ʨβ<��Ң/���=����Ơ`���W�-���o�ԃ5���=�޵���$��"+�4U�5�[o�R�L��~��-�.=��l�XT`�%QW��B�<���E�䤤#�tŵFm�ӑ�Pڟ:bT�a�ކ�Di�K���Žf��[|��T�����L�Մ x_}�i�k���n̝����1W���]�K�_�\�`t�5�*$�m5����S\e�S����匝*X�������d���J�ګﭓ�Cݭ{?$�O��3�SsGW�H����y�`�\$�i^����n�]��]
+PŗYt�����żWirl��i���{\��#���|;��bf�N�eT6���)EV�b�w�_-b�?=)�������\����D�3��,��nuP�# ����z^E�1E0��)���?m��߅�.>K�CͬU��g�,I|�R���1� ${=���0<�Tܟͷ�����(��õS�e�_o|!�;;�5�[0�ܺ�����?�Fb!U���2#����=����L��~�!��mM�[/�>��3T�);�'����\�Sz>����T�'��T�Ֆ]R:uߖ-�,Ȇ���U%q�j���#%�L�Gj{`��vꕜ�3Ŧ����b��|?.$}�U������O�qJ��T�)��=n+sH՚�3�ѱC��Q�������������{?~eN4?�5�fduN��C�:��D;L�ʚm'O���a���� j�{��
)�V�ݽ��V���ݡ��P��ݽh����Kp������d&���s��s��}&�ةHZ� m5˾6��m�$�t� ��R���'QƸ<���߮�z���27�-�k���0��� ��q�b����Y�LV�����_	ɉ2Q1��?����������	����|��7�����j�\����x	�kc��O�	�jMl�<�0��L���n��^�iD�Te�!�\1N�;�����_N�{�H�K�Ja�z\	�oi�.V�p�9��&y�%�Ia�s�� rv��q97;���4mI�/S�[BJ�i������D�(2��(Z�l'iw�E(�w�8=O8��������0b�sF��I���Y�6a!%�����T���
�Q<�ҏ��M%)��c=��">�����]�f{Y�Vg���iWW+����!=Z�Q�VWɏըU�aW�?P<Ib�<��JG��V��UfU���z��8�_ѧɂ%<���g���F�� s
[G��	&���c�PE�p��G ����pE���^r�Bt�J����-ͽ)��ճ���`��r<U}ŧn茴eA�)��K�_(p��/<�|�x �ېQ��b��0��"A�#*5[��շ�"3�X�`9$8}�h
A1�d5�5�_dd]X��q�n�sYo�o�:����.>�J�����o؄���(���)�b8_+ׂ׏n阬5 ǜ)����rS5Z�}B�NtqO���i�k���K��1�?�E:� �a�U�Q5#�O�v�<q�F��C&���B��Eג�JVj�+� f���	/�y�0 MM�rJ:W�)K�̷ߒ����He�~Z��ֶ/��sN�����cK`���:��ҏ��! $��Aĺ���V�ކ�Vru�7R[��N&�1T _RrfE$L0�ͱu��~���� �����Ç[���X��.ų�	\�ҩ0#1�¾��0��'�o=���'��9���[y���~=ykGPB����yؓȿߪ���4�:^WXm&�6�Ç����+�\� #޺�a\H���;��vc����}���>�R٪p��a}Z���v�<������!�8���S�ۨ����*0g�i���;"��3�'�7'����u��A�[<�5:����o����OI����E�+�:��O-��8-s���#���9o�c:���պ٬uM.m�Xj��HF��Z��4=)X:��3��ɵ1bvCw���O�� �b�z���U�����ǁ���q�vn�[n������.m=lC���8�0�m�9����]O�O���L~� a��lQԱTk���!i^$�_)��m������K�;<w����;�B��p�ۯ*o��1��m���(��emx���6!E�ɝ�������|�i���ݶ�atC_
�37�Jx�,d�D�o�ʝ=(j����]���F������Ot"zG��6z�ת�8��P�Dӎ��1����'���U��)��&8~
l���MC�,ju�3Y�������?%�_�����ܣ�����:�����i/0V�9�rsU^��۩ں^w��%����O����|\8��#���,���MA�e���o��[�҂��M`�ۚ^����-�J���L�A~7Iw=@1�ȿ��_*�ϩ��
^����uZ�<o���W*�QGl�}G�Jj��i��@z��QB����׾���',�&�dU�N�`�7�ܑ�k�lYs?��m$sv���1��n/���@១�{gc�MR����]��� �HV8� ���*Nƾ����fUi��B�L��LT��"�+iY��δ���I��PAw��s�=z�CdB1Cp������~�T�٢=oы~|������ku�2 ��s?�<2�kbE�����y��i=0��X�W���$�]�N'6~�#����R�/,v ȸ⿠��a��*�d�n���x@e��m\�lP:ة.3Š�n��/��R�\� �ۚ�'1:�V��K
8���pA��@
G�� BJ��e���^�Y�k4i���1�J�>,HČ���f��1F��J��=�ȱb�s�&D����,��po�GHe<MPH����������p��z`��{��*X]Xl�r��[�~3n�j�M�鳠���*?��ʷ��0'���/��w��wu&T��q��[�lr��1۲Z����;�,�J')���VN�(�(�Kq�z�\�:,�ٔ��`ɵ@�Ϣ�U������r�B(g.M�O�@�Ǝ��%�(P��dz=`�Cժ��B�jZ��Dђ5Ū�9�ll̓8y������a_�m�D	 5<��];�9V����ݹ�i���)0FT��E�,H�����/SNҦ���ڠS�)�]q�#{D�v��3��� *��.�u��6���ɘsH���E�X@~W�Q�r/�P)(����=j���D���Z����B�f=hC4!�z��g�Gs"r5t��:ܽ�m���+�
rD[��R��Y}�Ɓ��Ф�H��͉]��C��j��n	�iy��9��̮DG��2 �	p6��ς��<|�E-��Èe���P�q������+�Wl�|c�iB�WHmŇv���Ź�WxȂ�e����;U�`���h���k|��\ �;���e��^�,O�e�ц�K�����.�W�֛��ڗ��4E�~�L������� ���Yl�g��O�o���_x�!�.˲�:��kL���K�+en4��=>�8$|��n�n�@׼��X�5%��07]b�\i�W����r�}T�n�����N�V���$M���q?f �S��(�r�6� �q�S1uE��\��a�U�L�73}*j���f��ܡ�D��]�YQ}��ۣ�m}y�B5Aw�ZI��u?m}�OH�ܭ�0{k�q��&,���\���Zd�Pat</�m��s�7:/�h*�h:��V��11���r'���ش+��ᷧ�If���ߤ�!�}�.��������]	,�cpOd�h�ۧ��~�b�Xl���H����}&� k�>1r��Q��;�0W�,�����?�I�s)�!�5&q�Y:lk,�ݑ;)e����H;O�Y'�S�n_���~�l
��'��V���־�諺��X%��B��9�FU�$i�L����~�:�z���僘�̳��/#�l8Y����9�b[gۓ��~��B�W��g(�wg+?�v�y�T��4�@��ץJ��f����yaRE��|!=n�T�USh��oM���=�X�� 6�W;S����#^?6���Ȼ,hsW,B�D�XǊ 2g�|��T�� �(ֻk~��t��\�;`�%�/nw^�B�+� �U��ʉ�t�G~��k�r2�p��P��4!�o�j�y`�dHg�݇HG"����҃#�Ka��ސ�����xSl��,y-�>PܟH�bv�����o���{�dQ��#X)u��Z�O��F}�����閵.�Y����?��}�=�S�uyz��~_m�/��v=ҷ����ңT�z����sc���FfM�"h���I\����G��4�޸�?n�^rU?J̚�P������u��	JX�l�>��$�ն�n�����֍�j<9��IT�w��1�D�̃̔~�0>�t�,`L>�f
�#0j�� }Ѵ��D�����_ぺ��e�N�q�w�
!�4�)Q�+B���oWc#Y��hn�xB�@g�<z&��7�J��R#�542C��a�+(��tk�5k��kj�7�x�����-�ʍ�vY�aê���,x�����K���iƹ��6�O*YJT�RxV�8�M��e�MR��\�V���G9�!���ngo��2BG��d�$�?N�٤߇����|J��*�u��L��3%(�j�`�I������b��oK�s^�_��Wf0a��K����IY<�M^Rx���/���U�3~9�U'���߅��W4��L�(Ͼ���_����P�z�p0F��([��I��2�ǫ���d3��a?�܇�5������ɪV6���P��8UN�j	x#�Kؗ�DE��F���g�4��.��D�A��w���D��z��K.k8Z���B�)`�]�]�Q�arϺD���f�5�!�+��uZ���6�-��}���6�t2'x1$8i"-{��>�?}\|)y��ts�;�&<��zV.X��.x�:q��q!^��~=�ə.)�~�]�P�a��\�ÿ���,���0�_��b�<[J��_�ƿ�Q�U��'�tsjlƜb���ne�݆{��3����P��do�L͸:'���&���pPQ+�f�ǿ�<����Q�EP�1}�*����U�~f�x'W�Jeh��ΠvX$��uuZ�����2b(��D��hؽ:��"����������Be^&^<��8��Cr��NN�	�R5 \@�BA���X�M�q�p�"vaF t��Z�a�v@�(qpy�?v{!r����2�K��B! !���z+d(rn-sFd��yx��(-�m{��@
Y�d���!Y]=�ZHn� ?��@�0E��tiq�\e�y��c�jޢYh���Jb��7:�w�"M���H@ݎ�u(�z4מ0���ś	N9%�#����j�Rx%�NʠI�����+�/�DM}
2�4��c��� �"a����.:�8X���<�$��������z�8s#�P���7��\�׵5��OT��h�>���=bV���� m��on@�ceY�P���$1[���,
t����CWˁ;��^�/jS���	��-ؠdHՇɢ�m���P�����3�`Jʥ��`�a"%���b�9���ڟm����TS����f���7�s�BU���oC�����m%�¡{�k6����2�;�Ã�\��0Y�Ih�p}���,S��ѭ�0is�s$d���~�V��I�o#+v��!+N����l�n)�%ۏ����vx͆��IH��W��Z�#�fl ��
j��'��?��G�:/�\�#��]c��QF��[)I{��4�H�q��ڧ���Y��Rfdt�̵�������V����*�֖�0�g GQ�@�K��9�|��=�  qz�Q�*�R�U�L�Wb��N�hg�L*}&����rZ��܈VG�sPZ�^�<)XiF�˿�=���N������d����s�vL���C]#�[�1�I��x�*�����d�-<<�F�>�_��֚յj�z.(�s��а�KlS+̚���W�B�Y�Q��=N�W�^�l�f��P2���3� F�iVׂ.8����E����;��	��-�/鞢��4y?��5zʹ�z�T\�5���}n�̓�����q���~�ϯI\�ͩ�ѓ���lD{	:�.�g�,eL�����M��H�o����(rҖ�x}9�y�ؙ$S,�ϵ�C�����u���Ԇtu����v����N���ҝ�y>�3�d��8/}*7�Dj{���2-h��ɀ�[�{T���S!U�2�>皟�;����6ܠڐ��]��Z�� �{���<Su#�ռ(#:��N�����.YW[���N���V� H�e�נ��[mԺ�ǡ��P~`�2��&��2E]8�V�I��1N�}t,�)�}�*�8�PB�榗����ĭ���U�-�(v����;�Nze�li����r���g՞��Q:d�aY���o�km�W8�,D�yn��W�<�~�F�u�l���*���+%�	]�7��w����/F{������n^����8u�����/��I<&߭ۗ0~�|x��9������bָ�������z�J>=���{�{e�ƴ�=�-D[�+��"���N	E��_�w].q��2g�ƚ6�jiv�5֦Rl\ /�mI2WA�нi���5��������/���3���
�!�q0�il�K�A��ʈ��,ʀ�/�a^��E��|>�Խ�&�g$��ϊx�ED4!�-�߲��N�8���!�`+Q�K���\����������-}��(�l=��|�����O����u�@����@Y�����>�閜��wm�e�^��S�F�X6��ҋ8�Dʌ�
�bP�U�Z:��^h�hR��h����fՔ�സ��p�c���`��Dv�}_W?\Hb=O�+r�S��/�؅��+���n������4�8���TL���\����Fe������Ch �Ӊus~2o�q᫆��>x��H/������weI-~��J�T����:2"a�7�ND=E:��8���a����>X����<�T0�h����6���]:H��W��7
������_e�D�����THC�̫qe���aC��ڥr1�S�53�>�$rŝ��	X��(�����"��Qb,a�����Rx7W%�5}x�_���8������׹~�����{���|�ԭ��@�q`�X؈T	O�U����P��P�p�������!�B+���\����������?�GP���R6�ӏ�? ,��������7� c��o���V�.��b�t����T��˝)��C��q͹�=����Sc#E+�G_rX��������ǿ�4�H�W�3����!x��e�I�=�o�M� ���.N7�NγS���
���zM�tA�?���W���;y;Ĳ�Q��ǴGlk��jP j�ƨ񑤰�ib���N{{V�� 7�ߠ~���'�dӚIbׯ�QCĵ��m��/�k��zN<��2�V�mVI���'!�R'U�)�7�!�;���6N��V�������f�������*�j����|�FU�*ױ��M�����fċ���Ym��y]Z�D���S�ŀ�q(��F�h��2)���vI3aP�_���-��'�E3�Ծ$�IOn��n��J~�󦅓S�!>~��i�ߨ�z;t��;����������4b��Q���+�/]
�F��3�̳N���3n�X���{�d��1��"bL/���%A���e81�}��|�Y{F\Kp�6���ULG$?��U����	��v�"+r���i�Ww+=�Bd,��4���<��� �+�> �i��R����Ϯ��s��H��NXx��%��n͜�"�#/V��.=�`7c���3����Uz1L�O�LøO]�g#t���+O�Ʉ��$��g�@KzH��L�����iHl�����Q�T��U�h܃���O�r����m�aFl��M�����R���Y��qU��.
x$�ڞ��4�mT��z\��Qw�k�69���1O��%���vJ�����[�'N|d����'�XE��	�g��~��(�~֗T�V�״8����s���^����΅�,����[7&|�9Im$�i92����i�����a��q6��b(�B���+q2g:d6V�\7Һx����|�޷�#d���K�����4(��U>�,WhZoh��8���r�s�`ƻ��!lة�<E6b.T�coKsFR�J4��.Y�VC�V� A�E%d��ߝ�YKf�ذQ����2v@�{��%.l�U��'F�p���]��x?�f�C�XuuE[ye?��F?^��e��^l�F��p��|�:}���w\�*i�j��㴵��D��gʺ����Z�uL����S�E�_�prh��������ذ�FP��-鲫4ڎKM�~ԃ��j��F[���������R �,̀���{���n�
 r�g��_����LC'�u���ٶQ:�W���_ۏsT��E�!��/���e�������c� )�|��S!0h	$Ў��h>Ȧ�r��F-���\��I_�.�E��b��*��ܱtr���Rk��J7B\� �N�����Z��JՓ2�	���`X�^��M�uU��y��iW�TW��>%���5ƅO��P�)�t�������;_��+� �Q�FSK�|���U{a� ���R���p;�o�l��V�� �������݄�*)ml>l�^\P]�6���/\f��p��Q�e��q���D,�i������z,e��r��x�;�yw�&q�e��x���	Y�	�-�ߋ���A�����sv��7Hy��6�4���!�Z�r�P�E��$�<��b���<������p��oԍ�V������^��v������\-C�,@�w��������t� ���tW��?�e�"lc���\�9��ܢ�O��)�F���m�e�OL���!�LI��D�w�G�?��ܭ��vl�ɺD�ƣ�N���R'�G;�#y%B��Ԅ�r/� ;E�'��zTx�h���m�r��4�g ��o�������\�_~j���_~C�R���������2N�VoD�>�X;�!�nR~Ps��.��VY��͐��|�̜��1@}�M_Ay|ѡ7=K�K�C����|�P���H��9�G}��,!Q&]���P~Z��(;�L�����+�yxo��9��{�N�w&�$�A(�
���F�O�m�zB���lK��F���+��Cܕ�n1ǌHGxwO~ϭD��V�d����[^��%���hd۩\9RLQ��:�>�k?*
�Xa������w}����)2W6W�b�`��R�C�{��������).lb��Y�����p'5a�5���g`�,�F�a5M�Q���>��(��D{��[�'ǩ�_�#ɦ�X<C����Ro�8"���3L 4u?$�v��@�h֛<˸K>��0�:ڛભ	��� �
_�l�9��o�v��������޼�`@��)�?����֎$խ�#o���ZK���R���e�/��o��0�j��i��(I���M�v�P�_�u5V\Oz@�}�򪳚��-�V(u�j�H�KE�^�!q؈,�:� �{^Ծɤ"��y�h�5K�	�Iڭ	���z|3�s�R�]�L�
m�B��NT���k4k�M�0<���cfXQ��FŻ�t�H���'�߅�b�@�jܥ>�񶿿�8[JFk��%Q�?L�v�&����/�ٕiCW]�J7R
��bV�+��(�9*�
R�E�0�ߟTi�kq�Q�9�u�"ס[c�����i��K���HQED+��4
P���0����	�W�i���j+
�	2�R�(����f܎̙�5���+;ʐ{��W&�K��y��gocZ:?��v?�{l��Z���,�� J_����յ��8�06}�O�����W��r6����IZ����&*\��&	����4��I��LkK�{{�����`ή�F�p���:ѩ��}�t���qF,V�> �wx���2��Cd#��,9,�hϺ�_�w{Bs����搶��IkM�'�(s�D��ji��@��O��Pw�5=��*�ap��2��CO���Ϩ�*��#_B$��fI�,v�f�܏��F���� V� '��u�g�-�Ɠ������T�����F��O��+䟔���{6�ŵ�Z5�KCڊ�a�ƨQ���µ` ����*�����=u�n[������M���S5�m1��%�x�9+GΤG�}�\�邼��"i�� Lr��;��D�  $����A�W~�+oh��I^�ǲ���B�+�Yh{� ~��G968V��r�>|$w2���/
RU<t�m�[i8��	�lx,9������O����T�vf��s������t��y��[n��1�c5xd��Ͷ=��{߾,�fĘj2l�˰
�s�f���.���Hb]�7H j����&�ӌ蟀����uN[	�����zW����ML�[Cw=�>���!Ħ���������U��b�c��R���)�������!��S%b�-9�Ȝ{'�����"Z5*���B����T�Eڝc��K������\H�ω�>�T�Uⱔ_%l�;y^��Z��8�Z�N���_�E����aM �-pat����,<*W�����X>���i�b?Uk��P�°:�p�floޙUE�c_N/��u:.QX"l�̂"P�K4M}A�O�bo�P����m�~[ߏ�ڊ�0�_{�M�ᚵՉ[�(�9/֐R6�����F��a���Ň�/S�j"�S������x'���D�EN� bBPi/)�{ϰLK4�"s�ئ�`T�W�+z	#-M��S&R&�ɌQ냷	�
n�j`G�Oa��I��� ���J��cOW!*I��RIʵ��ϠI�Ⓦ�t�TϞ�ȅ@�k��`��iW�'�{��<擰Z�bΙ�Z�!�|�e��j����ȏ�Ƀ�#�Y�Px��r�`���i�$�5X��i��fƠ��/��I�z��:o8>!��Z70eq��T���^ҭ�!B�wP� ���I�������}?}��S��0�3�+DI���ͣ�FD�@�D��?�~"OH�����M5����R7N�,�9�Y8�A�`[�x�R�?!m9�uR�0�ݑ?S~\��#7�q��� ���\�,ذ��w0��:ߣ��l��0�cH!ϣW�LK�L��DV��o��x��e�h%�v�^Y)�j�W�i��������AP��x��7��{��u�"�߃�٬�"��6 Tn3J.���M�>zE�ru��8�ꯁA�KF��G�lf�4Ą�!2"���]=���`3�&֍'-T/o��S��pƚb��B��Q�|:f;��PG�izӷ��@�����ҷ^�I�'�Ŏ��>|�Gg\�v����H�$�۴���b[��(�N8
"S ��A�h%A���,嗒����W���Q"�D���ؓl�!I��T�=k~�JV�q��/75�E���R}�c�1r�̙UT5��Fop@	�K'g2Ŭ��� %��q�P���xh��	a����n��q�y��!�1�G�K�ڥ�\� �5�~��"	������U����E%l�n4}��~�m �#ЃW�m�L���aY��j�n<���:�`H��9���Q�ݼ?pH1H)���t��b���϶M��3���ƯN�t����cݢK��8lTc|��0>�z���uwi�?ވ�>�C���<7��Dd�]��/�,G�æ�0cQs�;���^��	���Y�sƠ��[+e��͸m8l0n�|���9�!	?��W�-Ʈ�~!�;Z���P��׬T:���( ����/�����VV ��x�WX Z*Z0�}9+ۃ{>뽟����e?���A�{$Vq�:"��R�9	b֠Q��K�)� ��;Q���a�ī��@��V�������DڊR�Q�hGd]Y�B1��G�bh;z��b�إa���\ߖ��͝Z��R��J�F���įq�(�:�A���;������������F����&������>!��P�	�3�r�w5����w�nDseO�-����.�@L�U}4�;�7��	y�A��� ��H���XT�2i�56�t�]0�~�o녚ւ3��cL�K�H������!k�`��C���7��L�t5pN�)Г��YK9�:&�^M�=�8B?��<�3%"��m
�x��ʢu{Ӏ$���-9�f�[a�@��[������2ܶ��*����	�7{�S�č��|�C����qԯ�p,���¼�N����(-S#N���� ޽���l��������?H�Pq�}��k/�Um-뤜|���)�^�������B�(��4��q��_؍��/N���l2�h� ]j�_{,��p�]��	(��������HY]���5wL�����~�����Y�zϾ���2�AO�R�Tݠ�ru\�J��
��	m�r��0h�m@�=��]�qZʭ]�_MC�h7ƻ[�W�ky%�.�po��*��g�H��'���iC�П,D�����;�x>i.�I{*���	�"m�Υ�->�*���K�^��j��L�4j/�jt�Y̹�/��)��l����?	_z�[.W�����_�Ux�B���KC �m6gy"�"7�cl8B�՟�������������3м�7���.�|���i�$��w$�ϫ��-Y��c��=5wf��ac�t��fAA)dz�?�������X��z�ӡʧ�"����`ת��6-zolVq�v|��*7G��=���n�ަ��IK����ǽ�_��6)��3|`����Ò���4���tQ���Г�+��~��),��XxO����B����ΘS,��rC%�H`��r�-��8�V�]Z;�c#��}�~���!�[Q/vхXl�y?�xÝ�7Bů�>��CZ@!��E����<���@M�`���>@�]���!_Et�����E��e���5]������jw��o/3-�`O�����0����
�mZ+��^ż?��V}f�7��hʓW1VT�wc�0���j�9���@�MѺrc�U�iǏ<r,��u�8�e	��5�V�Xʯ)Һ^NـQ�8:]�<��o�m���v;�.���Tqѽ�>���S�XM"Fh,�!�����@.<Vu'L��P��'Dw���gE׳j� �'��C,IM�'Y���{������9;�����Ž*��>Lm"��~���,:�2w5UZ�=��{wH��K�)�k�m�d����kge�d�����0�|�@�q�0��A%wVJ�
���jċ�Rv<�~OS�H��a5�ͧMۺ�����ۨ�!0h#���'�_�пoPΥ�[� ��G��EAR+\�5�C�������1)�-�hW�Pp�JV\��N����x�yE��g���	���/9����zL���\�>��������?*�}�r�
b���uv��	�����Q��%����>됮���T)�_��L��O�Aoь�w�|�o� F<�*��QwF�����#��2¿}�or�L�/h���5M�+]�t�Z=,�3�Ib`��qLV:��<����ӛ��S��{櫅� E���zݖ�M���v�+�w~sYR�`��=���}���5��{��6j��F�V"d5����8W2);s���WKJp#��:݋w[�m�̳z���)��^z��<���V�1��(��[��j���K�(�	e� U8�`�7i�^�^��m6{��Oy�{�BW���b��ʹ�2�^7t��%�Ѐ,h�p�Q0�p��7XY���7�e��g��WW�3j���պ�3e4i+���c7x���I�ر��Σy�|=�ms-�`�����K��=�`�|!��ˋ��|R���j�lr�x��Ꮿ@R��n-J�G�q�VKQ�xD/��z��������k�;�l�I���	aX���b����.���!�Ӵ�5�g5�!��χX�U��0�@�㞝�z����YR���n�T|q4Nn�b�p�1�s&U��l�W���������������2����aE;\��k�D>��sn!����2���ads�X8`N����iE�%�8�����Ck�~)|xΖ�N�JZi��qU�Z�����G�^�N��!��>�&���a�S��rt�������	�7�`#U+m�Ε�����ZLh���nZ�9՟uy'�&@;D�{�\���k��X�4w��7C�q��{�v���%���~1Y6j�M�8O���\o����[���[�luI�~��k��9�-a��iLD��5Ά�ԜT�rf� ����o���,��wф/���I�
�S=���H;���߰��S �EnyR�4H1A�UǾ�` �k����b�׎�%��X9 Fcg�e�;e��,oS��
�C�T5쯌N_����k��/�cn`�ڼ�F&RW�eg'���Ǯ���ӎ�*���u)*�6��ʳ;�k�� 0��z�����zg��2�����!mn�,�v���*`ޓu@��i�^�a	w��P- �͖�w`([���MO���ge��iZ5$��V�q@����Ui���j�{"�V''���xk��Ex��c�׍H0Q����	%��u܃����(��<��&�L�a�VwI�A��P�R�i��L�5D����n�"=~��Y�P�7l���X����R���WR
�7�e�������Ϸ����؅\w؆1޽$�n�u�r���ЋU��1|�Ä�Hr��Β�I{U�F��4�ma�Jȿ�$��d�cC:�f8l���Le����"�3���S�h�d�H�X�;��L����w�{�ظ�.7�2�D���|�(_K`3w�8p�r�
�]T�z5#���I	/��!'���?�՜��Ab�-��ŊxG�}�I�'��J6l�'a���o^H�<O���/�7�O����f/fR�aR{9_Ԡ��|$Qc��<�4ʂ�wS*a��55T?�#�4�F���bA����!^��̷lm'��$~�L��H�1?ܤ���D��@����Ùf��"j�5��8`2���^��	XP�s:I�(�+&�|���u�Ε�7��k����[�Х#�W��z<�����X���6FzcWɸ.ڴ�6u���G|�Dx�����5�Đ��R�F�Ǔ>��g�����^fv�Φ���&ѧdo�^�1�\���9k��A�\�ƷC�߻����i�͟��v�#zX��;琂��KW���Ut^���3�k�hv��e4���+)�t���+���~,����4�2<�˰�?}!�p���{x����aFE�~����hI@��R��OXDO8��Aڅ�Iq�󩯖��h�ֽ/-�B��P(%�e{� ŋ��i_�\|�<�gC��Co������gnj:��໥���@t�B����9�7]�!�#�
�,��@`�3P�� ���y��g��՟��C@�4d�1��!#�Rf�9"��En	-�Ԍ0��������Q�k�զ1+M��ƢɳR�B���j�	�r����k�~�17��.묾�.uw������4',kȝ�x�����9��2"�ݝx��ߌ���y�{���4�+#Hْ@I���Z��hP�n�3g1g׬Ԉ��E�ý��f\�	bE����?��� ��tk6��������rM�\�jj�V�{�����V�?d��2d&cU�T �����Q�V"&��v�\Br�&� /|¿{�npYsE�mx]VXU(�==7�}��d}�?�7\&_ㅄЈ2̮G�,s�98~?My���"�2��p�3���(�i�ԉ��	dq�&d
<>�f]���
�
A9$Rk%��W���
y�$E�XB_�W�'H��>��U�A?�@���n��o�ӎ��"�^3�F������xM���:oiG���H(ai�7^�Fq�q�
���>!�P���sb�������}�-�}�����<����'���&��J��������(��y�Kup��IBM��lXC7����\Q��?�u��Ih_QT׋$�|c�x[���������t�΁Q���BD��?�� ��<�#�E����r�͓Iw�o5�sn�-��5�Z��!��βpw-GuE�3�:]��4�0���ȰȰ�X��,����r�E�Jke;3�-�)޺;kn~��0\�g��t�����j&RĄ*���(�LKE�����Cu{����O4�mJ$���"��l�$�����Xn�)��mo��>�&�� #B�ȣ<`u��x�IU�r
��~i��m>~����$+��>�o��vx�¬�nc���b��
��b�5�BM�{4l�Ӹ*J���hc��%W�bw��[]1֗��,x�eMsZ�������8�Da���e�}V\[��+���Xr�CD��-"|*+�5G	��,E=+P�oe�G4���~�אÎC�Ā���r�H��?R7͋���Xx_�P����Q��;�;3���U�ǈ	��q7�9^�f�I���0�4�/�H\C��J���@c��Q�1>.h��
R�,
WY�Ke��g��y��P���R��s���'�9���R����m�Z��6�f����R������۫����]gB>w�+����5�g�+���������|NPx��Ǯ&@5B�����UH6� �<Q�@�O�4��j[�a�Ĉ:��������e�z.G1s]���v�PS�b�V��`��U`k����m��;�87z$/��S������Jb�&�&RnC�!�S�t��/���؅��+7�_D6�L�����}|��xG�E��!��&8�,r'13R-���鵯&�iF��=�b`Ζb}�v��v_L���1��+&#tOԶ�bNT���z���0�.���@����؊F9���c�/ƽ�R@/�炑����Wo�_!GX	f�������i�S�f|��jy/t.p�9d�. S�b���t�e���#�c
7�E�E5�$�q�vk�x����snM�<V�b�hc�ȹ�fF�r�vJ�H�G�F�IS_r���S΁���o�/����H3�范�r���g�Wo^���D�X)�|�]��c?� n�A��������ԧ�L������}貸���͝Wա2�7���z縺߸<[˶�m,�ji��Z沭�Zv-�Ɖ��9ٶ�=�s߿�����S]�O\x7P��>cpx6�8���R@�t��W�t���􅲬z��~�>V�Z����������J�
��L�'ފ9��aᕋ�ݛ��Y~�,&` Xo����&X��d�!u��a�+ځPb]+Dj�o�h߭��"RD�1���Y&h����c\���"+��D��q�R�'��L�C�5���/��j���+&P�����;�����.r�"�b�@Õ�$je<)�!�- ł�A�F2d�q�����'n��3�=~�sw�
Ne��Q�f*���Ѳ�OKÿ���uG�3�jͥ�ɠsR�5N�޴�}2���N_ 1)`��K�"���i��?I1#+ �1�G��H�_0~_M��/<M�V�g:1~L�v!����I�nU�w�ŨO�$'W�������#�~�@���5���LR\F/����7j:]O�`P*̞�:�v�|Ƴ}93}=PZ��L��������JZa�U�hHW�
&��~��2��k@U��P	�z/��h�&��� j�o"P������K���b�w��tE`dw���IS߬jܬjTb@~7F�6Q�
Q��v(H�,�_��;�1��G*�Ń.�-�x!bXA�X�B0l�9-�(6��퍄#6e93����bE ���\["v.���)^�H06�@J�X򣖛S��I�N�i����1����[��8�}:��?=��~�
��>f^ƨK��0v$��@fuP�n��r���u�'���5�~�8Xs[l	l88@�x(N�S�P�� �� ��q{-x�3��]՝��h��ŉ|�������d�҅x�KI��ᅌb�;ҝ?H�A
4�\Rq�!���ig�뵓��1ZU�����D��9�ᮬ�M��x��KA2w/t�tDK�DK�{%�!|s'��53�?\��3�J�▉�j�̙J�c�u��E���#��R$.��ڟ��.���T���x��������ٱ$pY�'��eG| �,oM]뻷
D�G��P��1R���&T��'�o eu�����a=w�g����S�;�j2����V�Z�VJo��W�9�j�7��N��:0�D"�Z�G﮵��/�J����s-��wZP fZNᆱ:�:�G�-*�:��*�U&v5U��#7{�ܩ>����t�}��gF�Q�
m	)J�F�C��@����5�j4sS+8�/�����ϰ!*�K:<��#�}.��O"m\�����8p���vgMr���~^e���EFe�!c��&Ր�j������^�����Y��V�i���)P����L���W��
^�r�(Q�a��d����f�W�k"�������q�#�e�W���/i�ٚs����PP�pQY�sY޽x�$m�:��X��g?	�$�z�0���:�ݹu��ĝ�^�/>e �Vfus"~Z��XR��ߌ<����u�^㸉xR���w�1.������a�n�R�oM3gy�[�w�#���?�8��vHC�~�I�~-]�b�}Q T_?Ve��^��q��f�@j��q����Mu�keD��	3t_�z�]s�N0���',���!�֯��V�`�_z��ebc���U�?����Y�ӑ�����QE�`-ܝ��>�s��;�܃ Dg_'�--f9�e�>/|��^����I��xJ�RT�K�[e��ѩ�e��Щ���Z/�Q�%����p��b����&���[џ�k� ���K�D3e���x�?H��G�HMw���'m97j�AY4a��p�{7jS�VR����S~��`�y���##0ӏ���.�U|>.�[��4�V���ٓ���ͩ�(#xkٞ/�λ��ʚ[�78K3�r��WM�2/���\���v䌩�V �M�z����.)�k���SJj�)�s�P���ޡb�~������J�=�A�U��^���]0u�t���3�7�b��dܒ��� ���:����2���6ˈT�u�n�i���2��x�<Bi�j��[;�EHgǍls�ٙ��l�:���`M%a;�����"�?��v�����:�X��j�#�Ò4w�HUp����։�q�"�|ÿ\��u��$�;4��i��T�a��ެ�Ǎ��p��FB�t��3҃N�H�������??r��$*W_+u�v���}�����P�����'RV�����S��p7\�y[:D������I�fj��a��Fa��1��=zYc��GL�^�7�`꼺[u�� ͅ����؍��:�Xh6y<~b���g/���Z����JT�*���٧�{�	�vn��6�&j�Г�&��o_���ML<A����n�7��$�/�h����/����P�	�!����`����-]�gi�De;�'2Cx�/8�S��2\��Dl�^G��y#�����(���cE�X�|Oϛ=�;�Bٙ�;Φ35��;��AF�%�mT��z�#K:Ԝ*�9�!=�_�הG�j��,f�� �p��ip�z��%���rh�d��։���p M_+4�Ȣ����-��Qߖ>��O-���Q�L��?~Ez��t�z;@g��6��O ��8JI�i-Tfd"�术 �����~�<W����c��}��ږ}��#����m����t�����س�6oc�ח�'C5����z�}E�ߋuu7?��X�|�Z���7���u�9�5�ҟx,�E�18p���ʥ�O��D� �^}���뮄�g�2�H�f�)�q�A(�_�:���p%��C�(!������ߢ��}XYX�	^����ԟ��1ዒ�f���kk6ܮ�QmAl�K��(�`�q�����@0w�l��E$��{�}m,	�PT=��q�������pu��B!�&��k���~ 7Եy�9���s�w[�����&#ɋ����_ۓ:0Ďj���e^<Qfѫ�	k�	2�X�Ge�k�SА�����tfu��^΂*v��QX]@1�U�����)}׍�}�re��w)�s�"�p= �b��?�<�����O�]�x/g0t��^��qҢ�{�) y8G�>>�\�@Z �i����^�@Eٌ(�!}�O=r0B�[&�Ay(���M�qG!�j�xH��B�4h,��aaqQ5i��ܴE��U��1������*L�1�S�>��=ќ8|�u��'eM�8���ך�+,���M�5���e߅a�B�� ·�C�j�I�h�E�����'�F���')#\���ד<�냞�i��)��I���8lP���2�  ��L��t#ò*����~"o�?�(���~�b�\��ox:,��j��tF<�F�;��X�e��VA9b�F���G�����C۳����(����?1!�t�K6�{���tY����PA��vG��I����<�VG���W�q.�eҦ�y/�O�b�+�mⴔ�&a*;��p�_��{v���'�5{6#�{��Q.$҅��&&��eF�3�r"Lu�vMa͉�R�s�ێ�&ΣЧP�1,U�yN����r���p��cn�JAҤް����1� �����\�-�W�y�����vq�E,<����v.79�gm�vt�*
��"M��ەI^�EM��.��{=�I�d���uc���^n��u?�פQ��A��i�
u}٬-�>�أ��2��8�g���x`1�fb����V|��M��b0)�C�^0\�b�@N	�����o�'��7U�O��8\Y�X`VAX@�\Ml����4݋�̧ou|��A]�͙����ۯ�����a�9'V'W	ٯ���X��^?��m� �|@�T�~��I��r+x�bEv��9���O|Y]ϡj(/dI�(��G�h����w�o�d�b2�ҕ��� ���H�a���@iW�$�s�R_��P>�A+0Еr<�|��O��r�a ���¼A�p̿���mlŷ:��U�C�� tz�R^����tⵂ��2�����p���A�B�9����f�ss�/���֔�T�`��6^D�щ���}�_�<#���%����y-�Q7�{����Y�|0v���V����G�?i/�os�
_b
�dr� ��{�M���,D<�1�	�@qg�v��pY���e/M-Ũ����BS\f;�����(�S�Q������ɍ�O.Hx�*�E�'��i�Ӵ�����.	3�֡�{A#aW��Uxh�AjNڠ�]Z��֓Inhum�I%���������~� tc�C�Rg���r���(<;>PP[�!p�Dfa�XM.�� �(�ep ��!:=7>�ŧ�3G�8�e�}������:�`v%x�u?u:��Ny�P�!j��kp�BI��0��)(��3SA��N�@��tO�mw��ʂ�I �
��Fۗ��#��7��_X�+���� �Ķ�e���>Ɠ��r����<תp�c(C��3ᦘ�eCi��K�3��{	c3rͩ4XeX�=&`��G�p18l]��#Bg�&#��/����!إ���*4(�Ȳ�H.GC���a&=;n��P��؋A�s��srF�e���]�z�jz��?����Lū�� ������T+���&{,�K��E��z����Vb�_93�)��$���+�>.����N0F@zs�2 Gύ*�s4i�Z)ړ��U!��2���Ln���wF�ҳ�-�Xx��1�KQ5�W�-��tӝ��~ou�e/�O�����;n��@ϡM[�u�1������W��g�����& <���ͱ*��rHR�e]���v�&���{���K8�:Ȱ%�&�iSg�l����; n�DE����z�ey�j���'PWW@w$�}k�Z�G��̝,Ν�23�B�f O<tC/H�<�LY4F4�
%���O��d�p�ؾ�]Ȍu����V��A����f��I����(�&-^+��x��}��T�24��C���8�FA-v�f���Fڍv���O�;�Kw�+���}���(�0<.��B_�'�0�� 2��ICٜ�4#U����щʿ����i��f�q��,��C���֦��Қ��c?%Wfh��>O[r�ᣰ�*LZ���5蠶��n��YCB��y0-d*�e�o�)����`o�x5��Mļ<�����s��_�cRQ�����M<�y�Nd�����
�~�Xw������Ў�]HC_f i+�z�H���Zj�  ��t�0i{"s̻�vx#q�D�}Y�ϱ����浓�%	Z�4�b�+'�BF���q�W^�|y��U�@I.���1UBb�Mֻ@�B�'&�� ��[�P�� ;m�2�h�pлv(�}�K#H��]c�pm�
d����~��d�Ǧ�f�EiE��7_�E)Qc�G�Ï�޿y�2��@Ƴj�q ޫ3�tM�@BT���{v`H}h�0<�������#���2)~s�y!_8�6D�nֳr�a�;5�M�4r���G0e�S�ɏ��*X�cy�ߗ�_��ǥغ���{����Z鼷q� ��K�g���[˘,Qx���W�J���""��$�*i���d���/���[2 F�1�*�Gw�Yu�V;�F| 8�2�5�"�g�ْ�8K��U=��&�.��.j���b�etA��Ye6�`�����>����P���� ���v��h��JĢ����+���E���vpp042"agǢ@����1u��x$�����3���my������T@l,Z��n�+����	`���"g)���g-4H��MД\x@޷k~��^���}���y��',��]�l�fy����B�Ub*/�Y�����|���hc�/�N�S�~k\��Y�M��f��X��8�H�36sͩ�'J���u�+n>�ly���
+Eq?[���v�L�=3�����֙}>ݸ��(v��N29?�A��mA�nB��WշfБc��A}� �\�w���yM�fគ�B
VVt~~~Y%%2}VbmNbmV.|�|�[K�6>ߊ��<�UU�.�]]��/�=!@�
��aF{���L�g/:��'�
���b����8�్���c%���wO��މ��m;���m�.��m�8X��^u�)d)���7��1�g���e[۽�a�ƫ��)o�������� ��z�0�B�� ���e��{<b/��d�p��'�2��GR&}�QÑc�毠�=���v'���f4�lC��O�C�wԅsܥ�bv��0�V�m��ƞ5���X,8Tp¥���"@ryu�3;;�357�&yxx�gb
�!Y�@�\����=��oڥ^�HHV���KNE�����ۊu������⧤Ux]�3�/�e`�.��B>kL��resw3���/!�B酤��Tt-�H��������O�;�ɶE(��H�V]����
}��j�ٽ#��ҰI#IG>�=�dV;ֈ��c�-y�vG�)�2����%�H�A������������ �W��.zpm)���|�2��������h�Q���W�o�iEm��Rr4g$h[qm�F5닺g�Ӝ7�SmѸ([cC�F��p��WWW�&�S��[��G!vMD ��(���c��D�����u|��S2��CW{d�YZ9ud�Z���R��Zl�޷�Á<�cw���(-;�-qO�qs�gw��}�k2�_���q��~>�%�L�
��s�	�h}�-���[�t����/����ck���.��{�,��[�;C�,1�+vJ����*�����oa����f=t˔]2J�V���y��O�~����˝!\���J��w[^���z�%M~K��Ri�l�����)(�IJJ���Q��~8��6\n�c��.�a̮*�
�Vě��f�LB""CC�B8����5k�����=l��1���U��ߕv޷�]�N�>�tx��NZJId�o�,���֚L��3A�p˱���ej55�� I?4����{�JC���X�&�^i��-zbԡ��e,��놵`Wdpp�dI��LYK��)���2�{����p��Pe�|rg`ݷ!��h�eЬ��E�yf�d�^�V��{~gF��T���?�Y�'b0�)������pZ�c7/�q$��U���3
��
�i��a��H#Z�c���e��ѫ��_!�o���|W4����Ĳ6G$���#���f:iQ��5-���̩3XR��|a�E�yة����i_����.�L��5��W}d��a?$��J���:��.�� 8e����C��ھ/U�i6S}5���\{Օ�J��LOS��b5�+���*"��G2���I�De)�h�`oŚ�w�l���_	999)��E���/��[JJjݲkP��E`4��jw�Hx��sji�_ `nq1\>�%��1��6dS�?�m�|����������bS��3�븗V�M���V���>���Ģ�����3���8M]dP��LΩTx�Ghݷ9���(�@��j f&�1�V1���Z)�r�@����>����b<5��� h�y���J�\��F��پĿ�S���Yr�:�9!<�r����S�ٓ{|d[���f6'����(Nw3\D�����U�2k�q�'�LTT ����Z̐�)��OG!�++GuZ�n8
��Doi&}>���0r���a�`�g�m��_�Ъx*w�K�j��'��bl/�Z��i%�=>���9��d�=1���{V'�HF`�Hʧw\��9`�l�O�?PA���V��T�|2�45|~tB�>z��Y�O!V��Y���
����幷p���U�&t?��S�=��c�Ff+,A�^��7I{=n���Ǿ(m��+��ѳ�[���^����!t��2]T�&��ՉK��d���0�������	��%�����S6Naُ<�d�P��]駡Ȗ���M����B�D%��D��%���o~Z��1*��7���}��b�D��|&���0�[����B%����8]�S���Jf5��]t;�*�^`���Gg1�: K�V�C$��<��,�ֺɍ�<���h#ϡ?0gs�	�fE�@Nd�V^�Z
�@��ڋ%݂���n���Q�=�^u��8y��]yڍ#�����b|}�^{�k��gb9����[m����|λ���F��$'(�y�Wg��}����nѸ�=�6�o�׏+;Rڌ*&.�:���b�wy5��N��&�Ax,y;$Hx�5���4�-���>#�īc�p���c�|Ӕ4�Q�Ss���O=WK����дV�m�/956�A�����Q�Δ�5L�W��"�|dO�,ѯ[�¤nu������'�D��E�*�������,�g���g�wd�dZe�E�I����H�j!*4.C�&�RV�T�;Ɩ�@������/�LR�ѷ�O�N�J��w<�s���rs�v��:�l8�M�uШ$A��m��H���-�Em+�/S꿍;��q������+:���X���#���(�q��f6'����
H��[k@���o�pl[��'�\Tn���yxLeZg1J�'���a̚������c��`ln]�@Gt�ŝ���͓5�U���`�'6����P����| n_���x�'P��mk�"�ru�����$�dC%M�I!�0��A�p}&�[Q5V|=��ͨf��&ŏ�������:�m�k"��/��$BR0����8C�G��}�7?"�4��<T����㕫�l������Y�J
Բ�khS,^B��H���Ң��͏ˬ�p�G��ק�<�c������o�xj�/_���6 a���bZ�%D�i�À7��)H,aB�&�U�K�`�HF# eC�!H��L��_t����,R`��y��'A��)��~��
�oy/,��Q���77����&t*N��S&Bt=9NFݕ(1�#���߆�w�8<.�)��
�
�L�LM�-՚i՚"�Nd�eddh�G�t_	EFE��)i,�BGW��p�#��B���hw�=���c	�����/c��F��2	�z|���={�	ԺAN1s�2�=fu2��&-�n\`H��ь&Mt�T`�{/R�e���V��s���E��(���:!�������`2͠��O�\�K���ޟ�S�[����ivOn�6�<��߾�t��M�9:�">B&��`�H��WVQ���8��o �H���m��퓭-���!y�qy�pu�ћ�/}W��Um��۶q�oc���#8S��5�!�$����]�OKS�o"��k������G�� 3����}Oە�I�xѱ�����j^������v�&��E��T44B��45g<����?��A�W��CX~�.	�@��``+�'I󖚋�t�z{'�wU>�$Ҧ����-tӰ���?�*�ƚ3�*y����q]n�)[.��}it0�7gٺ]��n7?D+���w�k��Y2�����#���x�����f�ok��Ǫ��@�����kX���]��ɊJ&��9T��uyyY�r�
F2p?i�Ÿ&��T�wڮ𠠡m����[]]�r�I`�0�������W��{nS.���pz�`<�[a�'2��4IO���pKRA�?��]ֈ�b\���3�	rЩP>tI~����%#��
q����'ݕG�vE0��W�Mm�O(�F� �� gUtu����r���A&�NC�u�q=Y�}e����
���~ő~E$�C��z�/$��H }(,
��u��6��T�E�G|S��d�j f��n�3�1}�o���_�V�JM��3s3Bwo�U*a��u��J�)k8�l����PV�`،�#�Wcw���{���� ����:��9���{3	�2�B��yC����-��TN�2ͪ��I���Ւ�S�}i�6��c�`=��؈+�~*ics��N�ز7��2���X������*A����/m;��u�'�,�Y���9_��yѠS�-\�)�?�ޗ�z��$c�F���X|>ſ�Z�p t2g�8 �CD�Zޅm���=������H���� 
�?e2e��	�`����7�;5;���N�;��8�-�9�8�$+ugB�`�W��ž:B�j?#̤�6�q��&��CXm�#D���'����x�ic�t�;t�`�Q�oU�`x�,Ŭ[��<M�������!�lڎ� �6҇_��*�F���5�s[�!1�)����b�1[�BB�����mx:q� ���BFOw&� MU���2M���zz�pWwٌ�����ť��>w������d2�k����J�ߧJ�u��5;���l�u�	�S�o��$uX��ɓ�.�?�A+F��\���/�۩; ��=�������&���	�޴�|٦J��Ȩ�Mbf��2e��?�|��oj2�����njq��T*>�1Q&g����a*��[��������@D�c�},�M��Lw�N�f�GLb��j5�H���V�| ̺�X�YϿ��H�)G�
��Ad�a[�aGa���t簅k�dа���c�h��A$3{�n����u�*�k9���P���m�Jqfpis3����e/k��)��7���Q�����0���E�����0���S(z��a.�4� �?f�1\�'!���,�����҇�vQXBD��/.ɥ��3޺��K�Fӝ)M9Z��y�i*R��GQQ�2���PT"�_#>:���ON�]i4ض�w�ׯ_����u1DJp/
�.�F\�4ߋ��(�q�����S����ҽ#�ہn��畍vh�>.�����������L���c��F�u[G6�)u̲��H����&��Bb;x��.��{0�դrZ������=41�?("�6��Á����=���"aa�S�E>4�d������A���c���Y�� �B4l%*h/�)����{�ά�X��TΥ� ��
l�|��1�/=r1���L����G*����N�{��Sވ�(�g`ɰ���{��H0��O�8)�`��!��݃0��֌�B�c2�2;;�m,����9���u����[���N�Cnoo�y���ഇ)��P���-O����[�WfL�c��
{_��
m�ib���2�(plW�:�5�� �v�(��G���~��%��~�l�d�p-i_�#NI1	�Z���$����2�� 8��Qy��Q3W���N.8�Z]�»c��Ե|��~g6�qb�#�w
�<����s�i�KIHq���XM��K��l�Awr%K��.����;�j����LD���Ā#�V���)�X6��Js(���Wx`]�����ƌ��W����&/��^X��30��L@���#:�¾*�,��<'��J\o�n�Y��Gk�����X|Ume��kꇀu���f�ǎD���v❝�� xeC�8���d����Ɲ�p/��󷈬n�w@o��Tm�l��~<?C�TwfmS0lTc��U�����Sj�{�-7<���_���1���@�ݠ�cs��Ŝ�B�o��j�*'w���J<����kDa}�I�s�M��H����-m�5�"de����ow,�� V�Xٍ�đ�"�����&��E�!�:�X����_��Gvѽ�)�Fjo�0��W*��o�* 2�]w��� �tFi^dj��R�y�6�N/�_Ǘr[�5I�F���Q71HVN0A9��w���rؠ������/y��"�p3���)#[!K�S�M���<$	`�v.{vk�Ubڒ�{Zi�����8��dM���D⃃�gE]lv�BQ��$/����D}f�m�2���8�h����8��6ҷ��u�A��	�L5�UA�`�L���@qi��U:T�e6����+g]z|�mߑk�&��@٭��[%�)>�7�� N�ud���cZ���!@��#>&����9�2b�D�A�:�U�p��D�Kd�q����r.�_H��#�?	
�-��RzO \H�˵���Z���jN��m���Nxf��6��Ed�P��O��$<k�FV��ѭ"#Q.x4V��U��\O�������qѽ�J��28�y���"��AA�2Mc�ŶC¡�C�ɹd&�o`	���õ�IV��Ft�U����f	�������>�����=~nFK?B���$���/�Is�j��$��U���#O2�.p��ŏl8ց|�+U{R�O�˽�׾"��g�`	x���X`�I(�O���*�TcP�׏y����cH:�� ��e�Z��/�W���!�⽤K��p��41�W@P�&�&�0���6Ձ��Y���m�,Ƒ�01f���%���Lݰf��{tg#��Ɍ�6�-���w-�{#�;�m�ʤ���ǈ�z�H�A�m[���=�+8��q�G<)�p��������mI��D�&����gĴ�)- k�5�4��e���R����ϗ�j�9z�9���-6�U��u�;�������c��(%���gt|}�ʃ��Y���x����@ \�ѵ��͗��}�DX�gd�ǫ,qx#�/�}ˉ�ͷOQMq[�gYᲺ�Lo����N�:H}���N��=���Qhꤹ��v�k�6z���Xn.��uʫ�Bx�2|�G�?	Wٲ��HÆ�k��������; {��Ңԭ?p5D�Qz��J�,][�N������|Xd���"�B� �(�Zg11 ���ׯ�1�XG��&�O�]����z�#��*�rA�JIⴐ=Y��{���>C����XPc�t�����c��-eja|QY��mj����`< �"�K�|��*Rs"[*W$k��
�g��ظ���;N?$믗S�-�ˍ���<99���|jE��Ź���5qY�&���Y%z�[Da��/K Q����d��� t~qo��Zu�Y^��B/�3Zmn�!+rz��
�7�5>OnBW��`+7��3�MH�%�ep^L�A��CCA䗒lib���oI��AF�mQ�B�VE�۞C�)3;G�y4�p�*�0�N�{�Wh��3�m���VS�ٯ���Hu���I;b�~�(+x7�#M�Z�V?Z��@�Ds�/��9�j�a4�v-��:��}�o�/����WO]�C�b����f
���is[[	E���G_1�yl�#l2�xA.X�`��J�����.��e�0U��Ow�!�ϱ�0Z�(��݄�h�������29�⛩�5�)���_e/g����&��dL�e7)�:�Bgі]/�b�k�%S���\�D���ix�J������8��r��][YF��S-]��#��Dز�9c�1�uZ	4	㞺��Æ��k��5�v!j�(R�y�\n*��8G,0k\�n�e�U��ؔv�b�}��.�o������L����?d��������c(��x#�>
�p��ZlB�M�R�'�t��[�W[/�����C�I���[<,���-{}�൩��Ku�(��7Î-����l�	VMLC4N�<3(�;`�ΘO;f�S$]�mН�W>�i~7Z�D�;���-Fz�������Aa�!mʡm!IG�bd��}B]/'�ۉJ��	}�_�KlV��G�J��Zq>�y����ഀC���dG�_g���c�5p��g
���_�vD������3�o'�L�����Z�G�����%T���	�������@��_V1�k�ti�5F���sHY#��~��)@j�|�f���tKۄ��
�m��c�n�ugT����p�!uO�Ϛ��&7�9��^�.��9���'��?8�Zvp-FW�(�K���{��� O�-x�Ļ��a�|΁�Ԅ
aF�}d&��]JD�?B��4�_&(q�	N���G���(��Z�g�ًtam�����.RW8�e��͖�O����l�|%#\^R�o2������Pwp^6l/�d�Yo Y@��"����T����e��D~�p�� ��<C5p2�0BD��������l��$�K0.瑣�9�q{�/�I�
��"��&Y�Ҳˋ
�i��ɐ����'���rB��Q�A���y���U0��>2�Į9��������Y���>a���]�挖6�]Y����0��L��A����O����m8��l��h�8���= �9k�&�2s�զO�U_`����̔�Y-��<~�n��݊>���O*n�-��!��������um�C�_��a�w��l��9z�P���>,�e�]�e_�= l�$�})_ƥ�x��`rE-�YQ'�o�ȳ�k|�Z�~�T�X��|0��{�^�%�HU9L]���������'��h��	�UYFFF@E�jdZZZs�ӗ!SS�u0l�$w^�/�@Wu�
������f[4+��4�@�'��u���M�>������x��`�Wc���o4�	��*%u�$��)SEꯉ}q�=�q�q�~�� 9�{�k3�y�����Id�_����zQ��l]
eؼ�)Cp��qZ�f�G|�� ӎ���q�;㱱5���?�����3Y��T�T�{ZHs���{��O��~ë*�8���T����t������\�fYmhj)�e"�fZ!��I�t�_0�N>2l��u�Y�꙽%ղ�%b1�kAh |�s� ^0���8x���4~_
�����d#�kƑZm���mn'��U���J���n;�M��R}�A#�=�r��>4�.F�7.o-ʹ�L*����kr��:!�|q������v�O.��z@I+*�E��(��f��ɒ���N�_�iy���O� �rm�)%!����侮��Z�:�P�{Uc��Y��\6�VLL�v�0ܺ������QY��OaZ��y��Yg��&�N�*�/��Pg��I��්ˤ�_����0f_m@jJ��3eYm6��
���8��@(A��mMػ�!G�U��?��^:�9��K�1Vjt����#1�e۝Z;���!Tv���]��:G[^?�B����o(n�����8�S� {����{��(o7Is��c����7�������I��B���'A����DAA��oUrR�;O,����
�����C[���	*�e k��7����EN̏���b�k���j�����
�W)m�x��o��K�n��tx��A� �9Uj���J"������s��Z���+ Q���d��a)����m�2��%��f<�:�4#��"VM��d��p7��[��~���΁*qo>>�P�#�x.sԷ�x(CiY �Sn��@�K)�U�R���@Q|�U�xfo9Ԗ��	����aDvf����|��W�ķTO�l��[�w�0�� <����S�FKm�ik}��B'��R+0�pF��AÔ?c����\��Bc�n��h�\�Y_���D���Y 5z�D*'�����m]����z9f��X����E��Z��,(��ʉ�{')����sH'L��ua�.���u*E0u����h�d$�����]�f63J��7.}��A�]]�J��8�.���������8['�������]��گ 鎀Z�s�����;Z����p��և=M"��ք�-�g�9�,�7�����lw��Iɮ_�2=��3����/�^�2b.��y(d���}�TR�h��&���T�d�
d`��1���=Q��W1���K��V������$�xv��y�6!S��~���aOE�$�7��0U!Ԧ����#���i^���/3����]CB�w����sG�I�+���Rs��yVE�r���t(��C����P������D�mC�ޥ��{�� P)�L}�$n���W��X{xY�p�UG��O�-�4�!�9�{騦�Ę=�O�Uϊ/�"d��|�s��m�7�qde�|X�>[��Кo�^lBa�J����7 (	y��Kdab#;���j"p�6��b����p��*!2~1���h>��8A���3�7���W�S�!D���z�#Ƕ���R�H��f����^��]�S����1�Y��1��67�]"����V�<�ж����*>������ �2�;[5꯵&-��bFy�z��p��f��9�Z����ܿ����ռ�O2,��?��b�U���u3l�mFt>]6���t,2�)aK����� ��x#e
�/A;u�c�P�s̦/?��g�o���.��#�ܩ�̓����:��쵧����l�U!�-Jo�V�'��܊�H�:h��	#��%Z��dӍ吐�/wk��7/�Kw����aҧ!��~����m���h��r�b��C���ャ;����F������<�4@5�`���Z0�b��Ҟ���u|?Rc܏t�T��}���1�� ��Z���-��l�kG,�K�&R�+G�·Hx�|�ý��*&?7��~h�d�����R���B��{�N��oT� �0l�auƸ%1�z���}�۠�89��!<~����0�U
�H�Is)�/�'�DBV?/��[f��kk�̃�6��TP0uȻ��lT7�q����jǴ{�%���&�l��k��(_�Y����׽���.��q�r�lS9�t�PW�w;����՘N�������=�F�|�;�Z�1�o�_�]]]��H���Y\�`a�Z2+�(���!A8qN_T��ɉ
=|]X$r�1�ɑ�����G�3��|�U\U��?*��tHw��� !ݍt�tw7Jw7l�;%���;�k�<���;?�x��s�9�7Ɯku����%��t7�2�J���=|��#�����>�g���.�ڼ�.�JW���os\=qc�x��Ht��r(�u`����EΥpRTs;j�� ����%.�<�Y7�L�}��R�.wH�{����2<I_�p�`���ŧ���]�c'?���FHI����?����Z����kw������<3,�9�(��<+�]����TV����߂���M��j �e�^
(�Q]�;�733����ٴ�o+k)x=�ܟ�鮴:Aт�d���p��=���]F�@�y�*|`�OD�ίIkT_�>S}K$���������#���pZj�d���NO~{%V�6��,/N�ލ�(S��Q7Rz�&�w���K%t8ꗟ.ZL�nhm;Z��#�҈1n8n�^�r%��=jC��lB�}�4���YD���{�Z��	Y��J>f���,�}�^3����=���`��lə�@��H(ʆ��^��V�?/ɹ�h�w�s�j��nN�ښGQ�=���{����%����f�����1����_��r��|��| sB�w�����_��Z����$�l��'�����nJ	4»�ǭK����,.ϩ����L�t����yrR��n��h���P�ʩ֣�Oz�=��gyޓ7��}��<���)8a�5��(�rgV�)2�PR����9�V��>�����vh]u�vG�ҏ�}4�4�o1->����-�I7c�Pb��������9H5��l�i��Tv���s���X}R�as�"�����ط���SW�~����%N���2���U;3��kY6�=��i�|����A��������8!��J2p1
��@�����ۋ@��u�qf=<�5D��$~��k�Z�k�I��dٻ��$�s��BL�,�3z��i&�;ެ�$��
�i{��n�W����޷��#x
�i		'7M�g=X��/:t�|0�z�jn�V'��"dY��J,�a�G3��r;������07�k�D�h��~r#��*���0���k� FФ>	9��kZu�=��?���J7��>�1r;�Zy"J��gc�*�Z���M���I�4u�0�����V�f�#���	��:���{ͭ�"a ��B�\��[��E&3�[)x�H��e� ����u�Rq�/2P���?��X�:�*P�����š�Ĕ�eigL���s���~�r�_�l3��i����Ѹtc���Eҹh��d�~훌���;-R��	��o�
&�ݗ�d�q[8��s��;'���'K=5O!nB���e-�{�b���#�+�_~S�.��ԭ��u��f|����Vѐ�Y���pj��ۮ��懽��N���9 �Ru����QM�{bԬq���r7(ƖK��rmd�-Yr9�.J�'��-�󳓛���6$���G{��h�br�'$��Ɖq}�/��`C��>��v��rR�^�Ae���و�Yϭ���P]�t����X�+��1ss��z߿���-ǖ�v\?���:S<�ϟΞ\��?��K��e9��U���l맪
3��'�E�Aq��3�MR]`���BZ�Ex�{>8�UH���续�J@Ta�uI��>R7��/"T���4Y�X̽��]���&�Y�T�U��a��P��
��?���PO���^��ЗI�t׃I+�8q���؟Cvo��Po)��W	��ݾp���[�K�nM��Z7?�t�9�V��x�7o��=�چ9-� ��~�\D	��G�xk�Hf�Zx�����-I٨T��;`�@�78�|��G���Χ0r��(e(1qUUU�S��}vc|�7�d���f��W��%��.%|Z=�6=^&O��/V�h&q�[b�9�-pg�.��^�	I��sQ��jzZ�zݒ�:ˑЬ��m�m Ok��K���~�F&VO#��8��S�z(�����ۣ���y+p%�ێ������܍X��^�9U����I�P��έ�ʱ��į��l��N��n�<�W@��(��\e@p �F����B�}����a��F�ԫ����JQ��H����[=��0���Wvqa�B7OO?�6�QZ��E�徭T���8�[U��6�����$����_�E��wH�u���+Aځ�����LJ���OI떊�qd���	�=�Ǖl�3cϏ{>VKU��F�]N�=p�R3V6��5"%���)�@�2>2{>2k��;BWIȂ}� !�W�l#30j���J�L����j��U�~O�;�uPj����k�X�g}D�m�����5�>��Sc�X.c�_M�mx�>�g��yv�U	T�%$��,1��Ι�����4{���7m̛Ǜ@ʳɶGR��iI���Q@�w�J��B��z�,V"o��C��2l0�E��O���F\.ݯF�NYdk�O��]�r���I�%��?�O��B��B���-��r!Q�2r��zJ�_1�}$Ff�K[�̛��vG���$�?Cy<_���E��?�qsg�� 5�pO����k~}e/t����%�4����;T�"9�`�۱ĐD�rD$�H��W���$�X1U0�-u)�v�g����I�.�:��D��8ܬ�����A��L�i��a�Ů@���c+=���sHAF�����{�J��E�=5���[�WfwF��R�`��ز{�����<�X��e<z{!IA�b� *���2O9�w((��~�j^��h�B�"�bd�$�>��Ds��@��EB	m���6����F?5q��,�Tɵ��u�/�q��6�Ƣ���~#��7�!fhkw2X̀p<N��F���btF/�����~g����+~�_�N�����AA��I߱|���E��t�����c$�( E�$	�29���nӗPw)�c�[�"��d���M��ǰ���bZ�k�`�t�NM���,x��{2��hn��~������y��$�,,�7Ӯ#�J����(b��	IƎ���5��$�!"�H�^���gA�KM�m6s�r@4]JEkٕK��q���>K)�`����z�*C,d����u�6ܥ�V�WXW�q]֣��\�SW�D���_8�?��i����El �i.}x��Ԕa�٪���YL5tt3�e��t��Z���]�(CF��ꊈǁ��v��Ov|�-q|A�'�C�d�1+,,�٨���l�Q>�Y<�#��-��s�		�Ԝ%��5L�ֆ����+q*�a��������Z�Չ[�$������I �TG@^u�)���͑P�j�H.\P��������?���j���R���������)T�re�xd����7恲>Z�e�Y��jI*4��ǂ�H�N�#{z��H�Lm�e�"��<BM��hm�pɹ�;�I:�cҊ��
+�#s�/M�>Hġ��-�X�2�-��;>\�Q*�m�ll��������!aX�v�(3b�7�X9�A��щ��k ��|}���lK����g��d��E`>��X��� =E'��Q���Ӹ�[���PN�W���f�#q^��u��PO�(���V�'��<rm=����N=T4�K��}Gj����<Q�U0�����Lv��|b����=�,cFZe���v{�yv���54$�=@׀�\�2����a˥�͈e����<��O�Srɓ�ϼ|�_��a�.�{���3�{�5����X�e�B��~��L&��0���A4�H��|>�:BJ[����c���ݗ��Y1���ga ��4�5��y����N��=��?�>RB[�tU�}�GJBrﾌ+z+h_���vP�-�/��k�m�c>F���������NQ ��O�Ks,�k��3��v"���:$,��3	����[MJ"��P�S�uq�����b�Y��S���ca�`�=v�f[�r=�zk�u���W����������2�����u������j�>��z;���KF�mػ�~~w.�LZ�j�|y����TV��xzAaa�|�Y�͆6"tt���l��?��u`��׌	:��jd�$�;�:^��=�
�����->��@�/8�eT��{{.k�Zc�n�5Λ#C�����-*��1._i9��t��"4:�WH<�C�����=��K�J��
En9f�e�����on���UT\��{�o OP��'�P�7k[�-��8�éʋ>k��W�(}��:��5 !����7%���)B�LQ���uj�����x(Q~A��bRX�Ԗ�Hu���9F�ztT�'L��힑$�e�*�wꛓ�K��4EQ�n/�IZ5�ޫ��N\�w��XQwlࣣC<i{�W�3�v� )
��aN��Y.�}#�<�6YϨ۝\��g�����>>�Ib���1z!'����$�\,�	Ѐ`�	J5C}����$��(�w��jy$.F�گOuJ�b���2����.���5�JH���懎h���v!06C�w�9ʓe��O���v�I���}�OD���sOn�Ɔ� 1���+�U{F���z�⠼)W�O.�`͞���j9l�X9��L�/\�?�:p�[BW�SҞ��5�����':Kᬐ"��c�x���1��4�FA�x>么I��6��
Fx�J�f
�����)�ML]�g�h0�7����M\ %%=�V�����IBWe���G%y��OHLL܉̶�~J����L�;�=K��>QAAA��q`p�u�a1�3]��ͬ�f�HS�����7Y�jM�;�Iint�w�X��j�#��{�<�M�	_>0,�t�7�v���緙��K}C$lDy���p���N0q�B�8����B�����R�O`�|xa�:G�E�����ڛ��K�Z��h@,�?!�{%�eJ���&�ܞ�vN��c��P�Ŋ�J+l�$��i;Wj:cxP�;T?�1���҄�ឝ��"!%�y�Ąj}c�lFݪ�Wdw�cFٰ���]2�� �T�+5��JQ]����28��'�iZ�x���+�?F3,�}GNmz�6�S�gו��W����L��ѽ�ه�L� d:?�@/t��.�W�4���n�)���P2%,�g���,jOn�|i���u�M�S��IsEb�����&���P"���JR���-%e��,ţYl�����OD7���z�`9��fh8��,���' #m���i��9�qU��Z�=ݖR� 0\��?�����b���_T1k�̔ՙ����lkk��	�)U��yG�+��.L妌�f^���kkor���e�6�3�R�
��^|P&.nH�d���jǫ�a`�� �M�#������k�XJ�ExR��������LTsJk�W�8�Lv� ��#_�Q�|T�-��pW:�U;�Dְ�c�]wY�4s'NiFo��mҿ��v�xc���bG@�
C���$�7�zv$g�B�������
eF��	��a���q�Igo���a24uu����^���8nJⲣX\Z�J��1kǁ�����Ggsjʏ&S'8� 2��͞C�kv-���}��g�]f
]T��,[z�4��,�ݹ����x�W���zg3~�K�|/�%'�YyJ��T$պ�[�`����'�E�Gh{��XJ�j�u�~��b�ܑ����/V��-��tO�L�ͭ�N#ߐ���ԃ%ǥ��ts	lq�d��_����$��b��ꅙ2�Rտ^�d�.�����q������B m�4�7M��-�;���{�K���$��,2)���etwsK��2o6�+�\�$b0�gD'W��6��?��Y����,0���MN(�u�md���dY?�����7��U;@�d�t��ٶV��%f��Ih{��W%�_ܨ�������.oUKM5�(��!Й����(�� ��y����i�P�V�]�����1�>F�jE���B���V��:`h��Q�Q��3����N//1�`���00*�\\�G/Q����~��d� ���:{���E/v��]@�L�9�:��QU��]s�>���cN���ŗ���Ϧj*��D��CT�, �~��*�J*s�\�`���1�9��Kc�1�Ќ(�K_I��c� ��~��|��������dӥFv�F� ��g��?I�l��z0e��8ɛ7o�����ؘ@����ǖ�F~3��f0�Z 	H�5��8U_6~��X�`�0�JǕ9Fnv+�ޒ\��z�^������}�>7��+¶��⬷d%��S}|j�oP͖�&��w��JJ-��B��)�l4M<�HYw��}�Y���5`�G��7������"	ko{y����f8������V?�K>#�S��q&?�i�^u2��RXZc3�_����k�ɒz�#�ƫko�F�9�)�f%�+ZEZ\!y1��OU���w�AG�1��-�%�M�������41V��k�j	�K�4��#�-G:�F����X T�`��ǒ�_���_������ް4=�,�/fLa�X�_��X���p�!Ёb&�/��S4_<]#����Uk�6��>/Yg�m�R���.�6^*페}N6��T�������c3�Vʑ�&���9/ͼ,Kr�I���AӜ\.F�%n���!v��i����:���>�)����G��$>���a�����@����?��Q\-�ߝo��U�BWoʐ��FUi<)2I�������tf�eCC=��H�yV�/P�=2��Uwo�⫲!ջ��s)8�}���fg��v�&�i��
ᷙ��qd�x��d�Q#R��4�� 2�ۇLvL�?��mO��t���EAR�������m<�����w5���/� b{}���XZ�ܧ6X�����x�����kZ،�܅����5��"�B�ZE���zS���Sj)���o5Omj���Y�L!e4�hg>�V���@t�����D�<�h���>��Dh/zd��h��Yz�O���I�D�$TP��������T:?��^��m,���>|�����%ÀG_	���,�����%1��ǃɕ�v�'1%377g�\��v9.*[(�dT��е�' GM.^-e���Шߒ�ϩ��+��8a�{a@�$��օn��s��q�E��i	���T��3��8}C��������?+p?��@l��xmA�K'����B���2XII��T���	��p$@���'�n ���c�zk���J����_��6��t���tӂS��u�A��՗��`�!oTյSr��+��̱S�ަ{��Wh~��˅>��dQ�7yLu@�Y��5i�hw���������t���w�1x����(����c4�c�&m�����p�p��I���_����t�;�+�^˫b!!!�Y�CW����0�^��dvkiR�[�p>�c�Z� rk���r	W2��S��>�&�gnHhe�!����ՒR<c xT�'�ʕC��S������qW%qSZ��b�w}�:L�Se�9��AQ�Ţ���h-�	�<Mzc��;8�ll1�,?�#]8�sň��Q��	�,P��	�\�30 ᆋ������F.���TB���"+j�����_�OM�����U(&����X�	�j5�G�g��Z�뎧L�,Dß��|��w���l�+�κYQX6G�ܧ�^�n��s��d��5�I׸��|�u;�m�5���i�֩��ii�z<p�
|�f�S�EE+������*�Ђ{���A�k;�B�NR�]Z" �PX�Q���#�ZU��E��#�����%:��ֶ3���W��z�0�׳�ŕ&7��;΅���(�=e�,�杫,t�F�4�W����C����WG�"��\�'����n��_����?a����Y/��w:�̷Ai�n�B���
�Kc���T��p>i��OA+�6���Ws�_�;������U�b`!��������/�����F�������>j���gV�l�D*�#]q\WBaL���Ҏt�7jNn3;'1�n&�V����>�}$&��X�[ݢq?f��Xk�W��LY�hc::I�z����)
��]˂��8�I���	g3�����`���f�R1c$=QùX�wz]�cɕF����"')j��\t;퀡h] ������S|��1�7�����v���Z��8n��Ku��c(-�))��e�S�������r��OVS���T���%'Ge��q�/#���l�������႗w.����!�k�5�]���-t�<�HҀ����;|��"" �/G�e�%�|d�J�N({������<��/��c^]��/�&E�n;�R���=�,[<M��Ƭ8�{:�� �����j�սo"�[�-`jZ�X� ����qp��WQK�^���rZ�:|�l6�d��l���X Y�;[.Ѕ{�d���PJ�'i�s�?�����4$:���z%k)ц=_�ǚ��ۦ�rF���������,��U���5������2����9�6n��-��h��ԟ�����BC}CCC���*T�Ui})"�6d�p�=�=&>O����!��)����>5Wd��\�Z�[�	�d�8Ek��I�)��3�%��2ͤ�A"�u~p-�n�l7N��4]�D�u�P/:��J�u��E��\̑%0���
n(����_zJ�^	 ����Y�Cj�GZZZ`����?���0ۻ�����A�i��/o���+J�W�M���������ؼ��S�oҍi%��t��9mFF���"�g)Q�U��ٱ�ö~Q����B@-�3٣ugnp� @�Rs���g��������ߞᮁ��Z��C~Kl�!�;�D������!����o
�ˏ WR����팲�"
$.j;{���yo�]�����8����*�2�BE��o�b�b�p��������JO����a���Xw�&�j����@��
�o��*�r�5��V?uY�e�N'vn��$e�S�����}q�$��[�oy�� ��lԷ7	�\g�^��w��Ο�s�Z !d���L]QL�� |"�
HXTk�ⱱ��v�:`#���9�?���$s뚓���d��ӧO���BA�qp@�>�%��2x�TB�rI�*D���������D:1R�6����0��i�-�4��j���R��>�pM��qPN��*ޅ
���"H��D���#��;���>�9��%�\!j��k(�E�a9��_T��v9���|��&KT�~���h^�x������IQ���n���Q��g,�Ʀ�O|��]w���u�����5���s3��!Y)��4nz3��x�1�h�	���z�u��3�?�r���*c�=u�CƇ��$�@>�䞤�w"�N���[���8�mv*�?���"��Ũ-H.0]w��C5�wQl[�X#���,` Z:���4�Ûm�����E��-�oB��~��a��j��,ˋ_v��Lǳ��GS����c���^������SY�g�	]|kr���̏���v󒵏�����h�_'7̪d�m�� �t0�f�j��B��ՅS1y������U�{z���B��ʢx�W`_</�h�j��,
/��߭���RGz��s�FZ�TD?�L��Yw���.9����lf�{���n"����� _.�����阛S#E&��f3t5�&{�����K��[r��Imjx�׶6Q�,���q�fѡ:����9/$o}���a=����r}�A�B}X��W�ح��x�X��22��>���&�:~F�.�y�4�� �$��cJ�4�g@�:��$pCG�J6�(�k%�s��d���@I�-}�I+�D"p�`Ee�0��|��B��t=�zsiq����a�oy��~��NnP+��ϥ}�����9����L���6Qc+'�{��BlU�u�w�{z�b����ED��a���w=i.>�4o�HBI֥�:V���n9��p���hd�v�c�d�]����`d��D<��e���/<��� �e�=��=LÿȨ` 0�b�R&�^ĴK)����T��CV����֊@�u��#��$Q�]8�޻&fp��jQ�^�˛����r�"�>�+$"�|�r�۠wH{�}0��<i�s@�s�F� [�o�"�?����سPOS4a�����w(p��)�]·��f����,����b�8���
���=���-T+Ȳz�+*P�{�>YZ��a�S�.]���!|�zp��ߙZ�П�$��c�&�^����bfF)��֣d)��!Kh�����Y�	]4;x-c)��<��
����(P�uhhi�U4�<���3,'��0=�]�Y�_R@DP����S��W��>����A�.�ЪW��,(��E~f����+������k�B�e���vJ�,;f����%��M�i�_߬���ֱ���$�BV4u�)��!��E�dP �:�3�k�[�P���0&��#'c�+� ;7 ���%�]]��J?	��8�'1S�а,e���O>P �g��u���� �Ɔq�3X}ѥ݅�ʎINN��i�o��hة�:��t�4Jk��!N�k�4�B�D�b�z��R�d�>�^���}�{��+^�R�s~hCR-�;�O�TYU�><�/pk�k������&�v%��K��C���R�[�-?�w�M[�շmxXn7�?��y�#�H��oX3����c��������vX0�����i9u��u�Ӵ�B��4�:k�:����>6�U��m5>��P��Qmu�l^�8����4���k'�c^w<'����A ���g��m��g�� tU���s"�� �jc����W�α�+�ndL⭜���m����Z:[K7M��FU9�R4��� ̊� Ê
�ៜ�<�(ъM6н�!!����?q����\��ձs��J�z>��-���p���$:`�N�΢>�6x�u��q��'���� ���w	��ʃ���.y�sOB�KIFe�7���K��i>-SH�����c� D�^���0� 뵻�h���+y-M�fU�hm�<>M��%����&OV�ؽ��%牑!���P�ִ2�H�3��
����B>��rۡ���q;w��Nd��!r��7E�2��g+K��	�Ǉ'ڰ��"ـ�@@�Ʀ�+ɀ���F��2����4�<!¾�c�6L���J�m'bm'*�ӖO��O���W�U�r�%��7�h����m��0wK����w�t��]q&�7%Gfx����<:L��DU�s" R׋��nLm�����Ʀ�qF1��(��Ș=�p��K�(r�@{6��u�6��
4t7J��]���x�'f��"b|JJ�x,Ef݌���?�?�r`�Ku�z�d3jPS}����,ܟݝ�'I8^���-z�$�*ܜW�}�u���q�y�xQ�j

��m9��Y�3&����2a8��+��v�x6u������e���+���ӽ���PV�!i˚�a�;��/=���b��z�Qyؙ�R��(s�Ġ���Z����²iũ��w.]|�"�2�fL���l��2eg�M���l�Ƈw�-+�����6p����?���K3�-,ҡ�o��t ��40 �Ÿ�gmH��!򤼵�9��_�� p�T�)Y��=�¯�����;2h5�m�e�����=����DE���s��gp$�kj��ܥJ[���۔�Y�~��<���n�P!N����/EI<6/�+$�*Q�"����X�`�da��47���Y���0Q����b�Y�q����Mg�(��f����Xv� -���`)_�]�Z���J���Z�.���ΚЪԔR��pٍ�y���������c�FD�B~���1��$,��D�a8�:l{0����Y���D5y'��if��r>���ĵ�q�p�oܷ�����0X|P!��ěz�k�f����;6����ܙ�&��N���.���E�؁ӵ@"

p�KبT�'-mW<��T}j�ܷY��/7�oDy~���MC��?U�J�H�7��i�yi}o&ט.
�X
!��,&EBhG[�r��_��OB�EΚz:0^����9�F�VE����`�k�ۑj���p8��3ty�4Ӧh�x�����m{$�jA	���p��RB��!�p��O��Q=�B�Wr3r|��E@�=����Z����S��O�x�W��nN���--�`�e��t�k<�Q�>���ӊ��K�78W�H��D�5n���b �(R]����i����E~�vDB^�}laa̵ie��1^�u���%_�l������H�+��}�/�C��A�D-^�0gs	��e�w['�PSS�'�/}>D�x����/��"\�Zi^��N@����р���W�s#>	0c�CQ|IK�W�����`��s�a��D��7�?+���Ǒ�����Gh�n��K��lawet�Τ
���1_�sr�;�rLH���#�F�M��wR"[W����	z�+�u�o�ҟ�Es�u�/�N��Y�o_Q|������.pR��O���I����b*���� �{77R�U �Ζ��p��2֡>�nM��<�s��&�`b����Ȝ;27uʦ�0d�6��
�n�����?�B�H�ʃ�s`i���h�05߰��R�b,3_-oNO�)��^��fM�J&**:����F��Sf �T���'���Cp	��HVg̒�?�� �@f��,4b���0��v�͉�w���92|�p����(�;ulP��@��䵩�}�2��РY/(R�c#b�RO��
��I�W�:�jt�͸f
���U�]^�~,b�G��S~jj����l+!�"
:�q����&��no�Ŭ�9E��Lx"���L����$	��
� ��#�\��_��"���b*�]F+3�j���%�A�9��] b��<\���Şb��¯LL��"Ѐ��l�~r��X���M.{��8����ej��7�F_Du��.e��Rv��X�-39B<���11��k�9C5v�k͵N�a�L��|�����"C�,~k�7s��gc^�C����� ����7���c :�Ń��Pz�,}���s#tkÚ{.���$��������{<5+��6����*�p{/)k�cPp����Lϗg��
�f��>�(:U11�5zy�V�D�1w,��DA������)���s����蚋VÔ]L����;��W��ױ�(K���TJ��v'��,�9_HO��(Yz���=?�Ht�j��@U�����=��p�������̌���$'?���M�eM�޼��S���xf���@�?XFq=��b����-E#P���}��r�?�p�s��O����-(p�F�Q)��ى��I��I]���ӌ���1K4��ا��yMʂ�"�"�$�K��&+x�.D��[�K|�Ncp�~f��܁Y%�#�[rz�|GW���eU�/����@ez���C�"_m_LiC�'�-d�(�����#�W	��I��8e27?�7_����$��d4�����G�H�p�=��؜���?�r"��աnN��K]�Dbuoc-�H�\S�*u����IW�d�ϼ����)� i�l@;�As:<9"�J�j���_�����o�hg�H��;��.�������å~��o{^*�Ǫ����N���]�+�a�&����?WvQ1�u�gBgma��^�����$�����ܮр�U�D����ť�͜�[�9�<�p�ʉ�21�N�8 ���B�D=]���<����k������׽���6�»W.��>�;����R��Eg^�4����y
�?�u]�L�`-��pQ���o�ُ�?�r�((C����M7��f��C�ڮ�"�Ӂ%����+Mwoo������}=z�W��M�����~܉�a�D��$����W��� ��6��qf�����,��\А��a[S#��v{�>	��e[-�'Ի��3�eG4�	K�`կa�`��N�℅��g+I�ܯu1_r7���i�YVW���G���B�@ �	�U<X�(���P�D�S��G�8f��VQ�%�[l�h��ϖ��lS"[��މVT�vH!ϯ��寿�G��N6OX��r��}}(���*0�B�1q$_H�Z3U"/��LH�bNIk`F$~��N�t�$U����bMք�`S����� �%?տO�D�·�w�=	����U�*U
�c�Ϙ<�h�w�b����[�x U�:5P���>f�v��U�^�]k�w�N��L]���8�ᗆ�|<4>�̬��bb�.Ą]��A�ǐRl���x� �p��s]y�
Ma��/>���҂���u�����ޓ 8��`�U��f��Ghf�L�����M�N��0�=�B����NI��D���D�O����Ӏ{����>W������v����z�PIs�j�,Q*��p��������ө�s/t9i��~�V����7��Bw��¡�w6�u/\V��o�E�zx)�12�h�vqÒ���-�>�"���L���uJ��%pG(�th�����X����I dꫵ�B��>�E@G�U��z2���S+�@�$�P1}����Id$�}�Mp?-���j��S��ۻL;{D�Ǝ��}���q���/}�o�ϫkҰ����.�{�cO �5�97F�Ĵ~����P �{C4��NHxG���п}�0;�O*���U�͛�v�>r5�h���I��)e*��.1Ck��'�f�҃�W+(Z]����u+-�*����z�?w��^�/<5P�����2G�c�K��6UD@�	O�^�m]WI�xԿ�7�q��\oG�w�8j���֦�N��l�!��P�0���ޱ��S��2**��n�t�U�I�"|�2e]��f?8!.��}�{ϗ��W�AS=���Kk��؀�a�xt�ohnf̺�b�͉�'DV��ǯ B�i��#�斖�"����W��ڶ����bJ�D)?���ׯU~�SY��X�NY��.�-U��a� �r�{W�>5N��P,
ԉ�'�2��v�b2�Ġeay�	�L��q�a���WI�b�&3h������s2z�y����C=--��D
��z ���������������K����jL4	g�`�[(ʋ���B�휫6�NJ���&��k��[����α)?�>@Ѐ>��fI�"$1;�2&����}��T��~���8�ri�\)���wս=@�)�/]�.������3-�N������M|Po;W�Ẽ�5NR��4+��7e�DH�b����Hf�6w�6=��)��z��˦q��wd*%�
ʦ���9�!c'*J+��R�{AKD8	����c�ᩣ/cZUh���1@~���r ��S��D!'���e
��bS(	��'��T�WB�d���#O^:�����e{����y�{��wtd�=��f�Z�(��N�Og,�(�{�)b���lǳj���A�xl�}=��|!��Lg���)H��\�%���5RG�8����*�m]���D°��	������~�=׫l� ���56��q��������+.�����f�_&(����X�ώ��#���ܛ[�Ɔ3�9P��!�^窞ܲK}nKU���p$� :�a�w�d��o� miS�})
urOA��ȶ_[���C)e9��f�+��Q�����Q�>��U)K��$��}BUs�F�e���P�:b��Lkqc)�}�o��U{w��N���Fˋ�/88*��65���H|v+�|�O<nQ�<c�7Ёb�,����R�9�:����T'�ppp�o�~��TA�RV(�����ME���%���r�vp¨Gb:���oMAi���[ ��O%�pA1��r�����x{��.�-�7B�|���>��'�6�S;����&�!3��N+3�SN̢]��`UKD�eê:}gm���X6|�DR\��S�_vmB�b�:j����dEY�=/�r�,�8�hk�����ʒc�Q�A�@GR̴^]N_��Hgo�2.}�L�zV=���!T���\�`<��R��dR/__R��[�:;�Q��� �Z-o��Qy�͢�f��xr��~Ѻ��y���L�X)�~����u- ��_R%0c�톯�k����߫�%N�6�p�U&�Ouu���*@i��Mk�_K���j|�<�����Q���&B��o*��p`F�)j��B�puu���΁9(\N���F��	' ��GTQ�gX"���O_����tA��C1o�����f`?��L-9߹�k0�~��r�/�Dh�^�*�9�j��̬��cJ�ʷ+k�L�
�'��R�$���N<=�5i9�o�b�b��\��
2�z���	�M@G�#4�=r����2�?.�fW��5k��"c��Sm���+�ĖUS�zl�yx�.�o��S��&�<T�T�<��G&�|�)�Ga�wi!���dMˊ�2$�E���NEK�ݡôG�+ǉ��|ט ��3,<����K���8��G]�v��i�*+wƙ+�A)M�x��/�X��fX"����\��Б�v�NUj=[���MS��UV���.�t~�0����;K�A�ꞈ�"F���z���%N9k$T1�e�C��S <��J`���>6�W�QW��|߭d������'pc<"e�>',�8}�'�-�c�}�?4�s��� |IX��Dh�t�C�`�_���e��SX��t�W>�����2VcC��?+�(��#��ᾦ4� �x>C���Y}���|ˌ+�PE�+:�7!s,�Y���E7m��ˌt�M5k?��my���C���v8_3���������~�e�q�0������%͢���Q�s�EUZbq���p�Q��jd�O��<s�=У�֎���ϡ�0���[N��A�j|y2����qJ3�Z�C�����Vl>����Ԏ�[_�U�u�"��H�R�Hw��"�����ݝR""��%%���]�9���{��;�y�^{���\{�}RL���<^�V�_2��k��Y0��.<�ϳ�[M������Ғ_��p��%���KeX!��6-f<K�[�,�v߿�n?T�lZ(�t�>���gu��\O�x����A);/��c`����9�h�'� �+�?�?VQ��i�(H���ڬ\��}���TVFM?�U�H���&��wx?� a��R������r�FV��NϨS��v�Gq@D������N�I!W���R���r�L
��P	�����9�J�EX�:t����bh_���Z-@틃���Y����ƈ�:j'�M+*��W=��3�>�%s�Zt]=ll��!w8/�𩘳�S�Y
��c���O�f�'�>ңK}f�g����Y[		�C�����F�1�S,�L*+�u^���A��*+�u�i�ވr���nȞ����hW^55��o%�����V}��U�WZ��-7��x{:^l�*�g~�X�fcYYY ���?e���{PFXѩo�7f�[��{�8$Wl�����9�o5|wO���DzH��I����J��4
[}VJ��]���r���C��Z��!j��=:9��\��!rw3�<_:K/�e�a|Y����M��C/��F�þR�Ӣ��WgpT��&�V�D�i2��Z�����gf3ծ���f"�]�'��$O<=a���0��i;�K�-w����#�nk(�MUb��N#��;�?NQ�p9!''_XjjA�������Jz���~�M�[��و:mWgCʼ�}A�!6�KL�H)֢��G.�lq�o��ϻ�b_+M���@�D����s���C���A�3���4�2���j|�����(<k�c7>0��=w��www����n�c�.��]f3��\����f��8?.8~�7G�����L�<<�9�Wx�+����E���� ��2(���)�����H�g��J��sp!�~���&X��L�h 4���;ȈauU��n�<ء�NU��O7�T�6�3��G��K�~�4��Д��¦�q��	xl���X�tm�L �a*D`-ͪ�DM;���=d�nLeR�������f�^�m���.+]b0Iᕺ�y��J�T�����wy���~J����E���S��;�60��H��D[P!��y#�/�F�اK	�r���nH@��쫋I����;Qh���h��K�7o��o�~*����!?�l��5��~���l����t����w�cRH
�3����v������/@L{؞_�)U;�XQPCr0dH�Ū�����tA9Yn�ؒ�"d{N��N�u}�~��fnn�����M��L��>�-����=� ���ܜTA?B�/�JJK�����J����ci��|�*�lbQ��A���O�m˝@HP���|��3���� �@��60P0���D��:$J ������t�Q�67W90�*l^��1�t���]DO��/�H�Ϩ��X��������D��ku�06�zxl��R�[��ޯ���c�T]�6������V@Ja���k6$Z�b�h���������D������n��L����LJ��#�B'(��7��}e&aؿ�y_��Y����%l4!͎y?���[  �ڢ�(��~��"ĆOS8���s�\y���C0Y�� �m'#LT!41���&�{�H������ X��l�E��UV(���U��fp
;n��\��}}�W�0Bm��c@�M��	�x�5F(�X�!E���M��</�V�Wx8Q~��	�@����Ѩ̕b��G�E&'�3��|�.`r8G�%�(2z�1?ET�Q�%�$��н�ʾq�mk�J>:�����@(��&өV�5}�)��V��+Y�QhH
�b$g�Td|ȴ�G�w�PN9f��0�)}"#�Z	r���8�b�~��)�;�%�h��K�@X�������fg˾S��:5y�1�/&��3�G ���	x� a��^�*���%���'�>��%�Dj����d��}�z���OF٣@����c<y�#�=*<D�k[[5y{[?L��=a�E�#�ɣ19?y�*u�{)���s�2��T�>��jw��k#��}�0p^�����/l������pgCD݆o�Y�9�ȗ��WW�@썡�+.������D��U� #;^�Yͷ�50�zܷ����A^]�3���ȑ���>M��5�Žŀ�^��^︰0�S���yb�u^�
�DX�%�5����'}}(=��-�����Ia�7\��fϜ���CUMu���s�=Kk�/I�\�x���x���_�i���3�r��Dqǧ��|y������������LD�cJEupj�3v����%!�q����%jc+O�������=[-�����=e+��踌�D�P&����[����g!����DC���.��}l���d�TOS뜷-�^ʇk�ܵ�%D�I�9U�e�Q�n��g�^\���,0����{��X��5�����5���[\{�}T����e8�K�G[	�xdpQ;I�[Q�����ǲ�߮o�ݶ��E���oX�ڹ C�*�� �wW����!!t��/�,=Q|Ёle�^����t��;�*��w��N�����������[X��������]�VY���I���:xu{�(\^Y�(��
��}H^�9�i}MZ�sj��8+� "V�L�ƒb�ցL��������x�/�̨�(��/&J>!������o�ް�q=�� �����`|=�PѦV"[T\	'Cg���㫕���͎9ۑ����(J��5*��y?2?�P����V���m��r�|�c�������`�6���s]������k˄#3ςEaB�8�3�P�f��|�s�wuu����/���ݼ/A�>�p���30CUCЍ�≖<�I�/�&�NG%����P8�y��ɧ���(`�~�������5�q�w}�+�����3ֺ���`T�\y�=�`nMh����߅^�v�$Ȍ��e�]0�(��£�Ϗ����ٸ��������F-�f��o�󏙆�
;t�B��9)��
^��E{��$4�(���=���)���r���	*g������4����0Z�����R�A=�78[�aFb��nS�Y����԰S�94�+;O(���d��D���]Ӝi��6��H�M7�!�&(��D�9�0dND��se���}W���|�}a��{���<SG���>F(ǆ��	������#�}����\���W�YH��_y�.O����k��v�]R��z��'ZC�4Dhb�į�PP�����7����;�2���6���;�_����F�IF�i��:<>N,���21Rfݣ+^I��M��{�;�/��w5���x�yg{��gf��� 󢊑 �/"u3B��I3�Q�X��iB�c����s�B�\Ը��i�ϲ�w���_��")�۽�s����+(�a���~�B)(��h���~�]Zc����~�yQrl�%�utr�L6u1fA�����4��#��U{8'-�x�!�R~c��X�U��-� ��?� Xԛ	�o�+5�xV���=]_83�Ѻ�?��t��e���Q�x_��L����E|ݘ�U'!��ע��V�����#�q%������E="�X�d4��$}_��;џ��~Q�CRU�P�������<� 0����t����QHG��s���p}#��(�\a[5���-���X��I1⯙�f���c���H�_�D�-�5�Oh��,��L){6���g�o��s}Xi���94�5������d�g3�ƭ��	�x�܁[��o��L�p6m����Ux�[N->q���|r��V��w��m�R����}5|fpK�
3�;�8�����bIX�T}�1
G�Ll�	՗[[����������Q��@��\�C�y��魬�ҽB��F�RPPP��hr0�x�q�����J��^��aMZ�C��~�ʫf�^��柹�T<S�A2K�7Q����Ef����B�,У�f��M�xT����jvjBmE3\\Z����8<����A�l��3�wl8������?T����,.����pt�_�����O�7qӾ~���K�R�X/�m�d~20�+7i{d5#�?S.� ���Dg֥�e�NF��J��ۮ�<������ܵV+{�橴��*Ǜ��BK���ƛ� #��x�u�����l�՗/�^Q�-
��	��ea��	�=wd������2���_|�f�C����[#ԟK�Ѽ�����(-��]��C��`ñ�B�,���N�:-
t/ 6���"���鏗Fǥ7��uf��/֔W>��g��W������u\�Y�=�u}�w?�?y�ş-�����s��N{��\��9����΄�w�.%w�ޢ�$Ll� 6Uƹ_��L�vS�}-)�[�e�G�^� n�<6��6k.i�!��1vZ�E�"m��1%S��vk����,K�#řb�J��YZٵ�|$�����CᧆWQ�[c\$���m�N�Ƌn���4M��=�]�"�
�c�1�s�.�+G|ՙ��|�+�9�?a��l�%�a"h��ak�q��t�a��ܥE
��$
�pP>�T��<ܖ8G.ײ����qW7��E���� 3�Ɖ�̛lԖ�~��rf���B�ܬ���������c����ƥ��1(-#�O�J��dͦ�{>�xwRk�NA����e:&�����w4"7���g�d�n�r�O��]3�=�꘿sFI����ǁD�/��@ 	#?>�-���|��7�����JI8Q`ѫ�~�~&��^\}ux7m�|]���v����Qu������x�D<��*u0"�R�)�&��N��K���K[�Ye�z��dTz��&�9;;�YYY_��:R�{��tr�f5:���������-J�a����7r#1��&	�G#��ɜ8y�k\��4�{<�_ ������2�0Q��W,u�{��R0C���ʰ|V�.ҠV�S�$��j�sxx<8�M�p6�#�~Q��1{�;�wwn�;4b b�qfe@�(K֮�DDEu�~*O�EeٹE�W�k]�69���F�{�hk۞�b��������y a�.++K�٠�z�r��qBB�ݾʮhQ�8z%�%����_��6د;�n��xnUi�q�\]^�N�i��j����^�L�i�Fg�}v���S�	mL[i�I�;���{AM�E�E�q��kgA�[����W~��O�w�B�V��M�,�7$�΀A|���F���e���##��{��?e_���a�xޥ�ŝ��*b��q������.�=o�S*�wU&���pb�������PF�>U�[1�sɐ�K8�ȳsZ��-�7�0���ך;���>����8n��(U�Q���6a�����r�R�Ԧ��D7����T�5�Z�XXgWd:QO!*?7ȇ{��#Y�{���23<����2r�?�-!@����J�ܿa���ۍ���9��&u�~z�.�2[a_���pwl6kgo�s����O#�js�q o���υ��#�5~����P@�F�$� Z4���| k�$7JH�C�|Wo_C�TWgqu�i��������;^�'��b�֖���~Z���=��BA�J<�GŘBTÚ{�a��
�����í�jZ'৬`8Sj-�� ���]�Z�d��J��2&>�@�)���a�c!I!pjD{�e$u �/�p(�é�LO�h�qk1��-6ǭI>����w�����ՓY��i
?��i�y��824O�u}�-�r��X&�M]9����H�y �
���s������%-L����;���	��'�y��aQ���UG�3.�)m.�D��lm۶F�[���	�&3*w���wW����lǹِlZ�v�˓����"D���od�(P�P��֒%t�\$���s���{����!\�����泽ޭ�_�ˈ�	�K&��yz����F
t]'��"J�4W�������{����i ���}��/�X-�v@]���A�����b5^���\4t��ы.��ӿ��@����c�:��
��64*���W۴j�"$@?�{� ��NOO�I�4�֨361Xݛ�^00��v�lY�A�˭�|���)Uh��O�,=��B��t�HJxH)�},$��q�=�e��B����Q�;dn��1��z���$ddD��j@LϬ'�uu�@��&�S	.�����n�m��� 7S4��q�'`�N������툧��Um��B�M$�W'�S@t�L��|@^����VTVv�h�^�h��Lvq��b�@3��c���>ԠC
	����)��<˕��<.�xf׆{�����.$
�ԇ+�vr�f8����]E�^}�J><ay�xRO�l�2{Ѓ�e_|s4�/]:'g'(γ&ޮ�&C�9v�`R�`�Jm�SS`2��(C���^�O����f��}�mC�D�5�;���T)$v�2��6��>�����2���(�U����.;�K�\�
ep?|Qe�>�x!QUSz
S��'hh�}��n���t��Bjk%*����z}��'H�=}}(+��!��+�^�QF��}��N֤��&#,�+�_)���(��T�m(������	�����"�4�9��%Tp�E�1������q�j�-/
��F'ޅ������h��s�[$�41UgS&�m������*�qgpdzÂS��®��>�����F������7��-�����&�(��0?~��ŧ��� C�֦io���P(b;�x�--����8�����٢���SƗ�<U�����8���;M��wgC���� 49:>�`a�f���;P{�է��%�����S9�+h�P�?|�s��`>!�����Gר�� 2ٖ{�-��v%^�/rϜ�L�k���r�7���n99�w

�@:!a�VMLLX:q��T��;L$�I�����V��r��gs��v�%�A�dd3� �%׏�M��ogX)#� 6��B��g��:Zߺ��>��Y"}\�!t7���@��6��|q+�Z�h�H`g��3��b��mM������l�uu�n���P=��,�-..���9�����<nj�$��D\�;v���	��~@$������5'�pZIQpq�300L4�7nP�㸤��q+�Q0[��>��SuZ7�=V���������^K W��$�w����m��<�9r{,��x�m�=�]��3�[XD���FDD�!�|�ƛ��B�P�F������J>���k!����BT<|����<�=��k��������rީ�ye~�QR!���%`��v�&~���W����!�
^�X"B����:ű����չ쉌@6`8���9f���
@/�H�����4�_UUӝ,����y�}���5��^"�A�M�+(�cI��{�Ei�Y��Ht����,H@󃣗���m�Fw�B�Y�ld� ME��$��w�f��qTS_���|�Z��ο~��;�EBE2o���7���h�� ��17���Ͽ��&��&	�^ ̔��3G����������9s�y`��0s����g����\^\�N.�3�;ڵ�V#������eG�����|dlf$����?��wxԍ�����Q@wWW��Z��wy�ncdJffL�����+ r�n��f�˥5�T�,�0j�.4�e<�r�b\x��뵱�[23�Yt%ӳ�qk���g��?a�����D���ͻ��0kWu>��  pPο��!���Û�#)q�a���Y�r�~�,A����%zAi�j�l9��)�o�ԩkZD@��ny�.�rY��	���f=n����4:�.o�Q��N�=��L��3RD*(*R���d�<�q�׼��U���T������[Z0�w�+mA�N�l[�x;-�wT�\��ܦl�_`#��R'�]ph~Bp�J��"�/�@?W)A�)����ɀ��U��d C��+RE��w@��I���9����KRVV,���O�4Tk�e;��%,L����Җ�LKv���a�_�]F��D��}��!6����x�����0�\#i�Zt�Zԅn[TK���a��iv�2�IN�H�Y'p[ 0��ǝ��&��S�o@#">�Қ�1�DHP0<&��C��X�`-��ظ�NB襧Ì�{|���#lk{�v�[�<͋��C���Nd��o벼J����9�l�6����i��� F>��\(��j�S�T"������,==(%* �c�>�zb;��y�9U� D����w���e�6�4�8�gl�Q���+�	�����x�l��fF&���������G޸ ��D0�MPb��)�]kWM�>����r��=���R��{Xs�bR}���O���V�M�+p.]'S9�ʂ��-�:��O=q�؇��y�p5 �8� N`{�,7`���3Ua1��E����e� q2���x�2/�`�
PR����m,�6����>m�5w��Q��ѓ`�r�'rnL�{W�P�$_`n..%-����)�M\�g���za?���'����J�R=K��-R��Ef�4��ao'<HW�###ш�^s�ugeW??�?�dp)$�Ѵ}�����GW�]M�׽�{q�T��:8��\�y���KLOxi��C]�;6����O���;���\r����ի�{C��u�7	S�'�y��*��cr�&�������~=θ>z��f�Gp���W=�M4?���PBC��R��4\J�4/�sҚ��/.zְ����j�T��r>����9k8R.<!�o���
S���[�l9��ȗ�{E��?����J�3A�=���j�X�]�3�������`��������Ka!���-��9�`1}�r@Ꮽ�L.Q�HB���2���p\"��c{�K�����v�`���[���y8u�&
� ʭ~��\?���i��y����^A-�g5�Uf�6D���-5��;#F˼F3# `��ܚ�	� ���(����������RKS�x�"ҕf�k��2��u.��l�S��F��i��,RZ�ܒ��W7�'���a2#�r��	o#qI1k'8SSӗ��q���˧�b�ε��H�T�g�����N5����#3�;y���(wեr���'o�����r���v�u�O��b#�1�r�M:�677�l��&~��To �x+����]��U��X�&��}gg�򂡢�i�=������c��W���N�� ���ئ����*�����'@f���M���:]����p<(27FP�g�_�7,G�Y��tx�l\R�Q�	,��,�ZX�yN6����'�Y�����6�N��R�*䵏������H�̢�=[���,��9�:v��SDj�nƵ���I�"�R~�ܿ"H\.�޸7e�'ܣ����/�"�����}rN���Q�~7{9��VB����%cI��l1rkIP��f��~N'��t��� ����]��e������q?z�K쑞����j1
(bɌ�%%�	n��+@�ު�?�6�${�E����i���Y�����5.= �zkk�Ll���_G�G%Id�eK+ �	���A���˗" 9���#��9��-�|�hS��
X�銦�~�ň���E����,,�̗���$����D��Wv�����N�'�3�Ljj������r1X�8�ӎ�W�$/�0p9�N�b�R�d�1�D� �8c���s�:'��Y�Dq�i��z�U	���@yynFt�9����_���p����H��Y�ٵ�&0\��3UcN�qT���l�	I��S�O�8�^���
�+����,�-Rk/m��p@�]�j�aw��RQ�<U	���p�
���@���?��BĤgC&/��j֧Od\����"�1����;n1A �A6���D����vOa vj�O����
��^0�8 �< 3yI�))�[k(9��f��01vځ^�
�>���1�ݹ=�h�C|�{v9�٣�����9�>ٌ����H@U��Jb��`s]�"��i������<.3�yЌ�� ˣO���D$5��jj�z�������{L���N��]�ٜ�2��k�Y��b��|�r���(��#.�a!�z;q$���!6bDZ�GpԾ�X�l��W��H�w�ߚ~{��&A!�'���ŕ%$EE6�ꪦ����g�b�*+��9���`�m�j���ت�Y���4�>����̾��,������gO�kz�θ Z/r�p8G�FBB����Fv���dLl��V�Q?([���Eגd�@z]Ã�,b�"�0����yǫb1��wC ����eiQ�ScѫSd�]��X2S�xG���ٙ�����a�����,Q�xU��C!��f�o���'&=�Ƕ�5�Bw�?���)����P�_�J��[�µNO�'���!����XX`L�Cu�V�9��o�E���	`WS*�?�Y87�%%:��, r�7��#�ϸ�5&Ό�&%�/*���\����X���:���s"YW
h���|$��4��_�0�����=�9b��8�_��}>h��d���Sɵ����R��x�|����ߛ��+,t�ޡ�}�Pl�.3����
uq�5!�ȎG��V52��9�ˋ�����sA+#�۝��M�A��&M0 ʵ�����oA@���r&rzJ�X	P+j�PӡR�[�J���B���b@���+3C4#��KL6~�hs�� ����R;���^��'N�p�ևA�e(p���FL��{�
���,�>����О��0������ͫ4';��ѣ��Q~e?i�99z䆇hU�������L�Ѥ$Vu6���(Y���j�)����v�T'���qwR�����N��|�(���5,:r�'�YZ&~i3׈uw�|��"��*��1yoL�\�}�˙Y�7e�c0��H�ep��{���3�d�� �����Я�~����r��z,����t���v�3��B��J��|o�h�e������W��L�qJ����D��RH,_��������YKl7w�$�%cSSQ�YX��12-���͍�xS��9�\��z��v�ybj
J�Jrl�i����L�.��^ =C%(4�vii	�	�<cаJ�ɂX3��hfs���������=�m�
�g&��0��󇧆��"ѕ���gg��Cw�<=2X������J���R1g�"b���?�}
���K�ّ������)i������l�Oʦ��9�*��#���SZ~�x��]sF@�&�asq��{���iY�}��:Sm�/�?�@7�y��p$�?�}zq�������NL���M�@K�,a��#���Ӥ�ќ�Oyo��v��Wspr�4�N��l_�t����W�z�#,��F�ҀV����I_0W^B!�2~��̈���h�&[�����>��@iTbN���=a��ׅA��E�ާ���KH�A0ttv�n�p�fJЁ���h:�j�Ub�5z~��M>'{�2ɹ�����6=��5����\\y"�;�۵YЍEҟ���{�S�2(3g穨���.G�[Ŧ������ ����� %Y//	{����g�&*6(�@��u��� �ݳO�\�GO�-�{��P'?���F�ihj���S!�_
lЧ?��x�J�����!�j��/����B�7}|���f�־�L�\��~����b��a-'c e �����o�b$��;H�(���n��6H�544���N����zK�-ј��%�j_�嗌�}�Fq�ڎm�{ޣ`�RT7������NX�$���l��:Eɾ���^�I"��=wJ�' ����t�N��0��M�� �~
/&6�� �GGGEF� �v��}ۯ��r�� �rj�GT�3��Vl
�%3��L����QL&�{����`��okk'c%}�p�!]N��S�/o|EO,��:cY)��G?䱖�Ic;{ۅ|����9��ע���#?|������*K��\a�2(ܗ��Qh�f�]������	,v~٢!��3��p<8;��lr�����mb��`)�����U[�<y%�.�Qj��l� ��6;;���GHx��Zh70^�W?��������/&��3[B��Ag�$�r<d���О>�%#g�������7T�ף2�p�]�����������7�I.�{꼡�w>�o�5�^��	��<N���M��葩��u��8ecD9��K�}�Pa��������U� �+/gW�y�#�RSd015�$s��h
�{�D���;8��jk[Z�1}�{У����?d-(T���LJ�V2����&"{�D��JE����^�������eD5@�����9�*�6j9�Ƿoo� ��7xp�"�ЭG� ��t@�����{5�ý����׎�<ǀ�{ q���� ���Q��=.�)�o��03gZQ�1�t@Qe��͉`ff��Y닷�\-I�[i�.���i��;��gH��ĻP�\,-����J�0�\���>Ļ��(죍�M_�ߖ��O�l��#��`��8�576�`+��H���KH��-�c�9�7����$���}Ȅ|�]2ee�@Pz2�P_��٧{��4&�� ��OM��~�P3�	�Xd>����?ڟ��&��l��Ui$���)e�A/��,M��yY�[�'�e`���d �5a���,;�*g��P���*Q��AS���F})\؅W4W������5 �_ �S���3�?<&6���y0�������{ee�Q��ӆ^�0 �T+��zF�RE>��������+%d�yyE�(*!,�ɦہ�a{tcNE'u��b�>
���rɠ�3��(kk��q͇z��'a���	���N�ſk�|`]HGUU5��B|:g;�;�����}cJɔ��/7��"�c1+܎Ch��h���g�̊�ÂD�  Q&#�����'#���J�U.�/~����Cu4<<����4���Y� j��~z~-K�vfϺ:n����S�tT}򗜉�U1�]�\�%L�D�J����I`��Q���g5K]�"�ƒ�Z塭��'J	�����?$�H7<==�B��)�::�`K�Ŝ�Qɠ�宅�2�[��w�l���x��j�_TO
Q��y�5lwo��-�\�x��Jh�j�F����SXx�����&F@��?���3��>UWGJ	e��z�xw���9����m44R7�	c,-��}d��.�b�T���s�k��s��%#�`�+�5�op-9��X��3cG�MQ�iE���2���Լ��I�Xb�ާ�A�#nn�]4� ylRby���?ןN�bZ=�3�m���Vykô��_�Yaoo�?(,�R���sr�� ��r����G���22X����v�V�,�l���� ���UH3o���ݐC�V#�,�o��.M`x�he}=�t۲ş�%C��̹�ZI�����*d	``ji/�P���!�(��#a1�ց��
]YYi��}�7����4�H�Q֡Ϸ�MWp�p������0JNA��g/	�έms V[N�Ȩ��[$P(�j��Y}}}�HD�Zȕ=H�CD��a"�<lJ�־���Ou�$�yG� X�>�(�l�r�M��X� �u��ث�s�.LLL����遟}���������=�È�����(��P��Y6*IBggg�-�>����P�yl���ظ�a���k J���
swvN΃�O`���	y����;�g�[��f��$''�嶂@?())�%����Ɠ	��y���{���7��͝	�1�oͮ�'�$�����G����#��r�&�L��� �b{�}p��ǣsk{�y�O��k,�����<�=DE��H98���ʐ<��@3���QJ#������A&����q���L	���e`A/IG-���K.'=_,���׬�X���`�@�[�������o"H@<LlsL�(ᕏ���h��>LQ~|�N�0[���ژ�XXD�Gn��a�^�>��	��x0�[jL��J�(/{���U�Y0�����[��d˸��m���.�d> ���� �5''�F�m�&+I��	���!����}�c���_�Ie�S�����777����U%;:����U)1Q^��gl'�������Z��F���Y耞+*�������'�1��M����[]��7<
��*'��%��5���!@X��Q* ����՜[2���/م�H]f�'>ufd&��Γ�R:���6�\X����a	�Oֿ��d�U�E�����>G�����޷Ύ ;�z��N���r'�d	^�y��\���S�� [c���|--��������Q�~֬�;ZT^�hb�D��v��<�<	��������'*-��-��r~�	�zDٽ���	�`y��e/��3B���	L��Y^Wɫ�C�u��N�7$�?�/�d�eT���Ȉ���Ԍ��ŉ��$�!-DEB �5�b|J1��S�r�p�ݽ�9����J�G���y>
�M�-���4 <�LW�ed�㾧~!v$��Ŷ�5������yr�>>���B�k��l������gW�K�m��	2�;�
´X�N�;�Rj̦� ��(Lo41Cy	۳��bG�m�����������R�
�ך�_"�N3t�t�9(���iF��KP�Eٔ�7M�E[���������,k���$ijՖx~`�/���-�v���BE-��/��]銘���3a.�2���s�{+i��j~aص�i~��G۾��%�[< �Gtu�����//!�Q�ܜ��hjX���C4�Ĕx'';{�333�ŕ?G����F��y��NQ=
ݛ|�]t��х�[�9CI�l���-Q)����b�1�5���]+��oK���[-�ڬBYa=: ��6��Pk5�6Ke-'oiUj��k�)noo7����[3{ۛ�*mi�p���{gu�(�_�7	�!�y��V0$99��ݦ�s���.l��?2,W�h�艊��sxr��{�qR[�����F���k��mB��Zuy�D�;����c�>�iV��y2qj)��(��D�	��p���`���i6�Z��+&!���g|ؘ�|
ͅ.#:�BT`Ŝ�������)p�W��k�~~
�;lT<�������
��c��9��������n:.�B�K�".�����Z5wM��c��W퉪�aii�z�s��&w�k���U8`;&�`�������omgC{$�ƫY�ȵ�?�to��i0//��P��ga��q����k� �+�?K��[|7��W7��FI�s^�^2�L���}s{���rJc2M^( ��	��Ȩ�rtҽ$��={Q�ݗ_	*I[�4|�;4��{��m#�ɪ���_�r)���U�x����a���8�H�n�o}�%K�s�3�ƀ�|�/,/E�l���C_�'��Skx1��3�d�ӘR�IU�d�+%~��k�,�~��.��F����� ��uߍ��J�1s,�4=PZ�~�y�Z�jd���z��3$��u�쑡�5J`�	� ތ����~�����,;}J�Ћ��\���c6�߸FaA�}'&��d)>ج�q;](>��)yM+�8�([��J���H� �n��9�qU��<:@E�V�f��a�*%#Ӷ��3O��V�׶MMP���vM)%�-p?:��ܹY%�3����;m�m������ i�:�JJ�A�.�d^;tY��79�Q�&&fFV�_����o���R,����f���ZX��|��4�5-�HMM=8<l�,5 R� ����u9��`Ⱦ�_�#_�Y��Ŧf��\#G􅖃#{H�~8ߨ���u�w�E��3ka�8�������x����\1B��(�cp����[�K�Ʈz/O��I�PN���G Ѣ�Hh��E�'(����W��i	#���6����&I�!�z���0�q1�=|�^G�O9 ۾w(�"nlD�:���$���(���y���S���m��X����b��Qrx�	6k��|>.{NX�JNK�@��'�T����2�2@��nˏ�g��h:U-:��,#�E��?�du=����,Q�õ%��v�U��D�"�����Zr�xwW��$�G'x��\s.�U�5��x%x���^V]V�����f�f���.?�!$�9Z����tR�����y˪{���³���e=+Q���b���o|kܪ}�Ŕ�z��m�Ƞ��v[�.�Q^oM�D���TD����R�ŊiZ�?j�������,�@�b����@b0`��
�vbW_��g��}`F?�~T�2z;�m��F���`Y��n�Y�i��c����l[����P��Y�����P ����UYx����֮�EMx��C��l����/xK�{^p���ʩ���kc!�h&��������/���}���(�W{�C�{�Z��e��J�F�9gxEZU�)�
s�Z�ۏ��F�)2!jν�CK��:�#�B~i�Yu�'�p�L"��5�k>i�2;���n#)�=��v�-����|L��A�K�f�����Q��^� ?]�\@���z���1���]u;���w� z�֌ْ�
R��ǹV�����o�$�p4�ѻ�����d\&��J���}��ק���!�i�+ �0�;�5@#��5��ɉ����|�O��Ds�C�#�r��741�6�{��D�����l~�(�5-�f��V�;��SBK� *N��"��ר���o�c��\N�ש覾����I��7ewƺ�y���kq��)�����4��йt��N\��o�AE184���xm���(h\e}
���gM����S��+�F���Zn�{8dptwoAw�8v���l䳛���e��텝�vaoP���5��'��oR	-���A�d~�y��_N�o0``�R4tB��;����|���E}�B���s������{k��b�l}jD�	槟�ة�o yF�_\G/F�����تI �B�b�������(�GIf_����Y�W�U���F9�F��ʒsך�Z�Ob��� �7Y��BxhX3D7��4{���r�gc���m\olj�SQ�%�v���v�G;i�O���ugq؇M�|��bb~�H��3�K�~�e�@%���!��H����uù�X ��7k0���B4�Y�SoWׄ�b�݃����I�5�� �$�CAwww�����p6��s�TQ5�W��ϻv���oa3��e�,�Ry�����+R���mj��Ӂ��a���|�i^������?R��,$�6=����W�����&z��$��a�جR4���������[x2��¾�������u�`�WĻ�2+�:@#d~��s��m����9U1�ѵt����%S���dHS�LlL�bª�d�@4.j�l-*)���PG��oz݋ɢ�@�=KG�����Yq�O�ӵ5�z%�LVk�
u��GO/���_�׳gO�ޙ�_����5�o���2�0��_�n��J�0�C�_� K}}�ͣ���qXz���z�4��`����D[���Q�6W:�8N%���-%{=��� I��/ԡ�.���w'���*�U2�G�a�kk@��C�)
#�Mnw�};�Z�P2�d1���l-{��F�	��� �I�� ���W:�����h�-Ŭ!�������C�#L��u�n�q�6�^
�*fh)+hu�i�����^�@�^]7ǉ����ᐗ�^Gy���!��c=��p/��F�D�y:���/���IB'�U�:M�+�j����)���qZ����-#�"A����U�c�Gx)�}��:SF�%�ɨ$~�
1�٦����"#soF|P�:�����CM�
J�3��v���䤥3�qA��W�k�������9%%-�7Xx�0�a�4����RZ-�!�����rZ�K�J��|���5t���O��d�գ�e��d���?�N'j�����l;�~�B��x����}t��Z���vrj�xz��+�yӊA��>�R[V�/�ʝ��K�M3-�'�����[.�@���e�8=���:TL�Aދ�l�z���AƔ��)��	Ke-��-��i�����%XE�&���BMw�^�-�?�8"E pa�7�Z�WJ#츫���>}^�֬wa(1h칻ӓl�����K���k����V*
gL
��	/�A D7�fc����R��{bt]Ի�D���Wr}̏�d�J0� �[�\�A��pd�ŹXV~��;Q���&���kp�F8��k��;܎-ы@�|�$�Hi����{����1�o�,��( �a��[_(��p���q�f� ��Y�}�%�����9����D� =�%����$�Oڶ(��t�7Obř��,�p�$���i�#��&�s�:�_W6�K���g�Xչ��4W��]���/ϴ�Ӧ��2V��G!�W������)~َ�eG,�000���;Ӄw�V��e?)�,U�W�����8�	��If�.E���,�k9{	Q� ���)����A����ò{%P�Ӝ�q���CP�k;�'�<%&����>x�1/ֹ�͠��@�"���E*�<�""�H��<�2��~��o�����Ư��/l���t������6��d��$~���M�i�= L
��Y������]qDGh���� �ͱ��,��q�2SeŘm8X~dWg~��A#���:�4�lC*\�^�}��I^��1�&����xc���G��(�v�R1yr�x)�M�v/e�O˘(���2�.��Jj����9�|�Z��������~�<��n��S�کz�z"M�R9����u7����I���ټ����|����d�0���{%�o�-��Ds�cq�Gn�K����x�Cթ�r�V�F������q͙e�7r �z�p΢��Y�F��[�o|X��(��u�?5�v+�����6���<��(�wə,�,�%V�Za1��o��<z��-s_�A�}��$g��Yk,���Z�4	�Z_������z�׮��q�K´�Aݾ�{wMJ�)�����(�N����Ki�A83\��(Fvv6򿲦Ht)l@f�74|��a��tv�c���tc�a���Nt���h";�8�D�ы�?܍Δ+��A�K<�2,<<��X��K[�h���4s^�	�K."�Q�?�)�ᥑR��h��1Ѥ:<n�a�NE���B�lB�]J�pE'����V|%�u�'��D(A D\���-y7�R�N'?>l	�=�ߏ����7w8bP�PӺli�0σ#���u�kuuu1��#"P��4$l�y2N�nխ+|9�/&��e!�&������w�b
n	��ѥY��2J�� �;�՛��AՅM�(A�MR�l0���9����P`@�.�k��r�؈�!#��U�6+MX����"�����v�F����NùyWw�}��O���hk�PI�׷�����7���\B߯ά��{W$���&z�~H�[4�\{ܶ6���[��z��8�
R���E��dثs����	\����ӊ+��ݵ8�Ā��F�2���'��	�t�Qegr�,��]�}	]c��Q����(yܢm:��#=���v�1���,<C����[{`��hf�T+��v�[��U�xy�{IΗ8����
���Υ�N��_��xeJgLr��F�t`�	j��v`�n�[���<|A9����|��l�լ�ZC�r�U��R�|�5�p����b·��X�F��A���+z
u�$�A�W�K�'Ӿ����P��u!�-<¦�a��F���͹=x��A�p�.Rjx߳����	�@et-������O4�jV��Ci�Э~�rB;22Ѝ_x��9F+k�<ezC6�献��`ee�����?M.ά?�"H��f�2f�='������e�c�'�����7�]
8����Б�?76.>�Ϣwٍ��[&�l��_1v%�[�4��=�=7MS %P	��<\"��Q������}N�80���J@16S)��{|���#-g�w�������MшI@ �;$���m��-�@�m�5�������u�5~����q��L��D��1aqq�"nPY'냭<�n-���'�h<���\��\�	/ا�|G���Xس�/���=bf��Zo��r<�f�3��l���t�3��TY�p=�@}��/_��7�GJ"��X�}�A��l~`�V��rM|ǽq���J�b=��>I��T_+��xq���P#t���v�NXm���T�p�_w_�BO?K�_0��iq\������)_#���گ?��%�]k�>�g=�}�6^��}Ky�*�I^�Q�e�Kڸ�[Z.�W���"��{�E_UM�G�O�طV��B3F�o�2������L��^��S�
�|�߳�d��k��ć����6	�	 *�^`Z��AC߾��C̞�t����ց� �h��:�Z|K��!�ʗZ���p�����R��!�恊�Y�A��"-�D�V���4!�WT����X׵Š�p73�N�U~+�ȶ���fk��^#(!��m�a]h�:��Y
;�`v�%�R�t��N,.T�3�J�l���k����|Xy k�2*�A�q��;K�5�����٤�(U��4^#A���+AYr��r�ʊ�'|��
��}�����דo�m����m���hjjf���"NoS��iq&誶?2��8�
�Zyy�G_YU�a����B���SK𓱌�*��}�lu�a]}�p�A�E����7	��t�x�F�,��A�߱�4�$b0�ӫ9(�y�����a"�<�Ѳ���Rw>_s�>و(NqG:����� �u0'�t8��1������8D���*Xk��^��?����P��)�K{��Ih�~b1N1�/s�q�9C)���wr/���*So���`��Ǚ�E�p�I�[	�o��\��yK�����'�m������>T�t��tt��$�lǭO&�Oc&�-��%�Q$�` 9Xa�b��f���S-�n4~�9�9qh��������I?�a�s9�_���W1�~U~k�{E�,�󑉾@}N��qKz�aU�U��VH��h��|?_ek���.��#�$�n���%$`�'��4uu����p��V�)P4���ckY2��T~�|�n������߽-<1EHO���~zb�[�?=s+���e���e��oV�H��<�<��Ѕ1V
Ԙ���(F+��VS$��hv�Q'�o�G�O矖����A�(����\3c7�n�vM�<��+>��@ˤ8��������Zeki97H�}�t|�d�ړ2�2�8�b�!㯓������H����r��jx7��=9r8�A%]����+ue��&�K�]`@=u���3��E��R�z�����7��lI�T��퉵t��z"���<�_[�3�T��Z���ꪊL�AQM�PίTCߒ����ܟ���EZ|��y6�z��J{�`�n�	魭b��_O��1vӂ�W4���ߟ��� �!�_v0	*�fڧ��{�Lںj����i�xe��U�E�����H�i�v��\���;ܖ�2�g��n�uG@!�׳>���[�¦�E%o��φ�Y%h!y*�$��]����;���O���$,%%�l���l#)|A' 3�7�&j�4"�M����y�����Q��Ҵ��C��+�ϊ�h�Qځ0��G��Ǐs��v GG1C�wv�u� ��0x7d	9_��	��,���� U(���㓢ʂ�'�Z������)�����qD����&�E�jZ���җ����t뒼���'�x��81Z�f�o��On�=���e�މ�φ.�߹��?���
M	"3��n�f|���=^�=>�F;��V������k��t�������DG�I;��'gQ����d��RRe*vSӓ�V�xq&��X˿xp��e%1û�|�0]��akm��6z5I5���QNG�~�DX.m
�9PpO��v"���Rr��:O�gy?v$�` +�
2����6�4��g�zO��=�4�vD�Z�#�.Q�H_Q	���9|��;6v��� ��(򲞆P�h�W`�vˑ,��^��.��Χ�w���ј��K{����6�����W��� ��!	�ό��U����D�['��Ϟ�/���h��S��|C��f�
�s��A��SJο���Z��	Fs��֨���)���ۗBߠ��4{?�~�X8Pc⾽����᧲x�]��Y� �%MI��fQ�&ob?ֹ��f��{�����M/��a�C�C�%vfE:�\��$:�վ{�Ik���UK@��x5��H6�|�c36��a͵G���{u��v6ub������4Ud�19��]�S������BL>hrۣ�Q���K��{�ξ�!HGc����@��Ǫ_7������iP�y6��,s�h�wC�v�Jk\]J8ޒ�
,n&*�m��������I�j�-�1��C�=�c^��YO�ҽjLqY�	@C[���z'=4IbBƦ�7���ܺU��gV��ӳ�ŏ��L��<�Z������іKƜa/�ÿ����"z��抩UV�5N×v��去�d���q�f+���l��\328���/���k雽G��×}�Q�f٧s�pK��XW��V�N�{�O�+�xkg}�h�mD#��I�P��׎\e�-W������m���d&W�$��V�Ņ�ʂ�1.m�n�)��T]׻���\�@?3O�W����k7l��r�%����_�����|����/dP�����B5Fp�)`�+��U��ϯ��>$O!�7��o*�\Q�pUwF���o2��8�#6��j�HxkC��t�ٌ�F���.�C0œ0 �_\�����1o<��N>���d�FI�N۝l�
��'��r�;0K��-iE��j�nS��:�~�֒�/�A�]���=uU�L�4��r݈�ԴJMJ�R���o���C��e��O��#���Ѿ��=)j�Ўy\n;\uYMj��CZ�1��(�(B$)��/��)0�}s�e��1���Ҫ�O� /� ��?!�y�p�3����+y{k	&n%u�Z���ߒ��V[����O|�ۆ�VQm����X�_��Om&�S�.�D���'P�K�FO� }���Nb����O(�h��{�X�pey|A�jNz00՚�wxil��͟�����#�TK"�#jj���/ӾA��e�z�j.�k۶��(�]F܏l�Ǔ݋�*�A�=�(Ą�# Vo*�kg��-e�� ~r��"S�oD�C�{E,�;��.CP,���Z��X�pw瓤�]���ة�P�H��EJ�h�t��q�g��~� O�XM��d���FV:W BO����[���̓{.���4?SW.12|�_9�v4uA�:��q���J&~VZUw���Q�.�zց-���8g��=�Jy��Z�<~��!�H>�����X1�t
�N_I�h�Ѥ|����⾋@+��r5Vh૰oH���aҫ���Gpق��犯ΜaJK!+_�L�ÿ4X����U�!/q�� ty������Ywh�r���BXfY�O�f�l�����i*�H�@Ś���}�P�:���cςH��⊱\H4V;`m�� �%SV�9�"¾�2n�Q�~ikw7�0���4q �)�#̍z�3KPf���%Şr�@D�u�R*<rtI�t�H���ۭ�����~�f29c���3gT����;�1Mi>�o3r�� 7 �b{G]d����T)[���ߚN9v.}o_���Ћ��,��_%	�%��4Iߖ��^�H����7׏�8�Z�R@<�b���J����Ѿ}�S/�>Ӄ��Dh������`#7r�
�W���@�&Hq�G�h[$��mߟS�W0�ɂɬ���6 S.��ݩ8b�xGGR���쀌�˶����5Ԥ�D�~]��IVX��G��~E��-�m�¿��h����CB!���|��..	n9��(�zGI���_7��֩eE��;��Y�"a	����2K�⃽����t �PO,�As=Dd�|G=g��R�՞��$=.Z���H�@�s����m
��q�����(O� ��v��b��AB}��8l9�;�&��������5F�>�=��3�Eŝ7tNZ���|w��H��W�~������[�3Rp񊉉�!��6I��O����Ok�U6�I^��'�_ܒSyO��������i@�Q훠�
�2��c��n�%�
��:����zj�b�Ne�B�>�?t����?)C=├�ʚ=����wnm	љ������2�)a��D��d�x*�M��X��`xtiIAG���]o�<O�l��	��`r��j۪���Z�g�Csp�7�ϋ$��X��J<�ڂ�J��7��,��i�����y�r�|�촁cF��1]�÷D'T��/3��?��r�|��i�۬E�n�����!D�vԄ9��X�))�+���6�>�]���� J���ς��F��'c��z#W+�KO���Z�C��J?�̃	Q���JoˊO��lj�7��.��-�Ϫ�#�{bPR����G6����]G`��/E�>+VL��s���5{:�uvO��l�Y��7L���aa!Q3ir��������3dŏwhg�|��E�z�S&�%�m�Qk��(��nE���F���|1�������B�4=�a���)ڣӳ����%'
js� �s��<}u�H'C]˭�x�$ǠǙ5Z�q[U�	�� ��f&Gr��> ��:�����&��A�2d�&��n�&�3Գ��ڟ��O���.�s̤��ua]3z���S@��L����<���_zvۑO����y)��&WGb��K+� �ܫ������jX�I(�����Wn�b��_ɩ�������&����'�o_��N�����?"�3�Cy�xAuʴ�:7Q�&�`c�b��ќ�d�E��bl�u~)�Ɲ"Q�`uΧV�7yJ�#0o-����dV.�wjD���2�<:�@����M�֝3[�x�_�[�Y�͑�}K�WM����J�1h�]M\<|�9U���$��DY"��;,�N���S�wo��,h�o�*Y[�A�j�|�LGF-c��~���X�qG��h])'5��� �sEsv�n��"n
��\��ȡ�߅������֭�AWa�û�6��"Oۻ9
�? ɴ�����#�����@�(crq��f ���|e��ݽ�.��C���x�����3�_�J�'��٘cU`y���
���sIM�\7w�9���~�	��l{gzj�8�Qʅ��ޕg��`�G��М�/���B��F6=��N��LbX�FP��;P����8ϢlD�뽃�j�Q��5מ���v��i ޱL�ѮF��v�G�<�eT����`�α��?΂��[=4ሀ�Z����������F��+Y/�������n=��V��~�q��?8�]=̏��+9�6���o�ll|�3�+`�J 6[��ߠ-t��IpijG6����h�����v�>H��F&l(C;8#��R7O���4C�����l���/
'Z�7��㉷w��m�,�1�I���1S^f�e5	���훉M)6E/�Sl����^ :㳈�Y�G�21wH��r
���KIyA��(DDԎ͹�Սs7�^V�o�y�EE�>w��T�~m�0M�ڮ��,I��O��d����G8�I��ƫ���������+�5�<��2B�9��+Bו��(�u������)��\�C~߸t�O�#4<+��r���#:)���M9�-��_��qHL�-f�����MZ"C3���KqȠ�Hе�VS�O��O�ŝw��]�}BbJ�F�&
��P3��M@@����Y�0��!9B�Rrxaa���Ǧ�Xa��X��t���gg�|�ѧ���l��s�e���/��~vɫ�T7y���TH�Є\���cF63>�q�I�|��;
�y�R��{B@��*�����F��Q�<�w�Ґ�H97v�d����"�Pb�l�����S��}�O�H�g�o�^d�����s�=ܘ·Ǳd��e{��3�H�48��B���IGҭoF�`���a������ڧC�ˬ����#OB�w8ޱAV4eВ���P�K���
�Cry��l^�r7E��@D/�m }�[��7�sl��9/xI̓$M���V��i{7�LM&r����8�Ο��Xj���&��~q��~��k�a�)�7@�S�;�k��;MfL�UJ��r��͜�E�z��|�)z�Zڸ�$`�h{ႃU#��o+;i��ޢxR�7_��jq+��hN��'����-�T̟��Ӊ~]u�.�L3��G� .=煄�-v�D���V>�[L<,k#B���~��Lה-��K������@�(�������}z~mwzH�zgTt:y�H�/>Fە'��^5�%mR�-���A��#�L���iK3-�	��=6�q���4�=c�M�YɣFW8��!��f�Ա��G]����^�[�� p-��h_Z������"�?���m.#k7C`l��0�O8j` 7�3l�r����}fv?��Bz�}��j�;c��%/��[�cs�\ 3[�W��͔�YP�?U�C>vڤ㨌_Fr����<��1p��5b�̳>*���wh'����r�x�!��t�h�Ĕ���̇��(��4�̹��%��nV�s���?Y&��k%��ʅ��Y��$�џwѶ�ؕ>�u/�R���ʎ�������}d3���)<��`3��X����X^+F�r���¯.�>(�D�ׯZ�D`\I0��>���]_��?x���R�?3�2��~�U��n&���r���~$ඝG�`�*����KbgX�� ^������IU6iy��"���zJ*lD��oc��� �w�`tm��ӫ�*n����k�h�+�o�lhԬ�ӂ���wA���IZ�P�����%�=���?�t�������k��2Q���a���E]�v`^��H�b�14ai�V4n�!��]��"���Z�]�\��d��J��<��pM:|��/l�����i���뤕�&u�&]M�@��N���ܮ��%����#b��N�6L2�'���C�%��%5��0D���z�u<�������O�G�r��� ˦Hɍ7�7u�j���g�>nL���������8_̇��Ԡn{o+0�Ӝ��n��ӳ=ݻ*�����/�J�%��	NJh�*"��b��y�	��#A~E/禖�ѕ��U^7���{�tG�\d���wv�6�y\D�Y��g����8�
O�Z/7��x�CD"��ҙ��/����?&�g�M�)^�E^;ƞ^\�+�Wi��q5�ȇ������~�&��d���^=�9K�6q���o�������ہ@���Y(B��X[L�"���Q|e��R�����i���H�G�1��N,BX�̤��
8���֤���"� |EA¿>�rF%qiAT5��!2�Js+�� 6/����a�����wQ�����\�|���1�u�6
�\:܅7<��vv���g�Ȱ��@>s�=�4�z���na����X,�Xdd���������ۦ�?�E^L]p^�]�h�F�rU� sn��8���Y#�ٓ��T����͚=,�b�X�!_��
���ӈq�_�x���z݁��xV2Q�dg�m�ۍ1��ņ7��	�K)�w�(�1�,��zGNJ���kz5Y�_Ts��m� AKt����)��[�)��d!���yg%Y����J.�ko���޿B�'���ݒ����}e#��K;���y�ӛ�5nN뇥�itM2�`T�#�꡾���,�fBe�a���񸈵v�����H�8
��s|z�C���(2��i����~TAAm�/�v�"M-�b�
�������.�L�zˍ�d.��:���?�pc2?�}�F��G�>?H{�N�H��$A���h��p�E��I�-��4cP$��Ei��Bz��6�Е�N�W}x��"G���\�r����܎���sKZRJ�B�_AGI	G�7��~���=�^�Hx�Vth2�u���<guNg��&@թ�x��|N7���Hx���=�?����
��AQ�	����W��!��!_��!c�us���Z�
�bњΣ���|y!\*�n��E�\��8/>���$��2�)��%�VL�2����fl��]�XHv��{�SWp-� @Q\n$����-צ�cL27�r#1�3Z왮��aٚ��Ә�R�s3v��o7OV���L����I����M�A��᷶3��F$�2E����_p��x�':ήȄ��x/e|�Fȿ_-mkb�?{�Ά
k��-�T$D&�>�O�~J�����Z�uާ7��pʪ��v�#r���u���l��?�Y��÷�w�.Gs�q6��������m�S4�S#6���Ӻ���K��"�7j���pX ����K,�5ۈ~Gh}�7^�(�b�!����~`�YyJ����JKY_�Q]�Z۶�w��]ow��׷��E*V���7�.c���-B�w]����"��HdS5��7x�"X�!��p�B/���fI�sW�F��	����9RMHY�,�l�����K����/���h"����$�L5j]]����� �	=u�����2-�A����ם x�"�P@.�;���J�q̭�/.ky�y]�]��u7��O�4C1�Ξ-�615���y����C�ڍ���D����=�u
璿����v���=�.tP��Ϙ�SGP;����j������w�c�H��/?����G��{��I��"͠�DJ9V��cL %_}��o�|���0V�Ɉgt6(�okW�#��y��;�Q��H�����zY�Q��,�{��b ���X��\�� ��+�ǽ�U�=Z�1��N��!�ۺ�B
>Q�]$u,u�����Y��͕��6E�=���۱J{�E��?�?�z��"M+���eU5u�4M!{��m7��]n���3��K�,G����4�A]!y�@���nT���z�  Om؎�\f{/�W}�O�}���0�"��x����u����QLVQ\\�]\�y��|��rp�_�:>wmr'[��Jc7��d��O�"Q�����FaZwB>��r_��1u\۰�M�s\N��ں���;F�?e�"0�* $�Cw�3={]3���sJ��mgY2|a�a��-��1�Q�[>�9E�g�d��"[������ͬ�K��b�Vy��S�b�p��K$�j��I�w������o���X=���fp9�ܭ��+K���)�(Q���/�4�!1�ų�S��;T��G�!�������fo'��>B[��Zo�DNl�Y�!]w��78��<D������5~4!]�4V�
�CH���$�DM�9:Qq�Ȋ��T���2x��Ĕ��*�:7D����c�e�Ag�f�f����-RNd����]�M��k�&��RPP�EW����"J_��x�X������}�ր�\F��Y��x�`�L��1b��l����sB֋&l�!���qTi�bsn��E-]ُb�転��\�O�->LO�n�� �
���{?[��P��ߞ�?/I��2�J:�K���۞ ��)��$����JT�ݯ�p��߿�V/TVV��V����h_
l�Sa��e����aX�#C���T|޲�@�ė����R�9�.��3r�R%�b�@�������pϓ=��f��7Ѽ�5��H�!�L�so����c��}0-z5�Ø	@��ӭ�+Y9~���ֿ�#��ɑ/�.�Ӥ�;D`�QVьWei�q����°�&@
t��D;��4��S��루[�=c�Nο���6]]=/mb+���V���)�v8�%ϫ4��F�:3�[��ʬؕ�M�9���%���jQ5R��g�F�9�i2۝��9�H�c/���lJ�o�qA�pX��kl��X����5���*�_(VM���}g{�L"fo��h?3U(����.�\ɕ��ęA&��UW�0ZڏO�0o����E�7�O���p�:[������x�y���'9G�2T�K%����N�hǀ�I����\���@A��~���h�P�=06���΂&�]]�ík�1���h�;˧��^���5t�b�[P�l���lt�uy��a+�R!���	����F�Ce��S���~���}�Ac�`�Q��4(U!x~^�yrJ�N�*a!��[x���Rxz.�}-��˵/�D�ё�u�Y�Q���bP�0����-��G8�'rZ��G�o0�%=� �b�*K8.$j�B.be��7�5K�7�t�[��j� ���"PX��&G�xvyޣ�%��q����ȁR��VB�	 }�B�E�M�I�2}�����)�����Yj�&n"@�
��/�OQ��G���v�Ȅ���9�H��Ô���X����� �":ڛNDM�Nܩ�����B�+��Or�>�u5�^���콝����m}�\�)�z�
j�==��p?��ю9�M�ixfϼ���[�~D;��I�r���'�-^i|ړ�������ܹ�J9�'���u����r�e��ގ���S\`Δ��P=��W
u�$-��纹�9*7{�c�����NNҷK���t�q��t"R�m9h��Xo���_�yWbsg;�DGC#��v�L�t�>�H����i$�
݀���!�Ə�c�:�
̅�,�������`�Q3�e�9�.������+)���zVb�i�WPds��a�� kyO/�����W��?lX���a�7]�!cԔ����//%��H���~���r7Zۈ��S�axA;�Y?��o��޸�-]���j��ݙ��4r��SQ�����Ȋ���@�ٗ����C����[��F��{Zܜ�x
�0�rL�}��Dv�jnn�(�� V^p���j���\�W��.�k�팤l7��:����8��V��7��BҼ��:z!���dO�7-_���~���-�9p��AS�'������x&5a�%+/�?��	����86Y�H���,c��y&�c��U������?�Z=�u�)����}3t��;L�^�Mj�xk�L�znZ�R��wF��HP�h��H�,	a)Y�?N��V�xљ�[d�絧��q��B�Cdj���J�4ި2�d_��igU���P�H��� �t~�.m�5uZ\6��e	�"T6�~��r�N�έ_��@޳�R��>cmmu
�u�=(��zbڑ���<}t߅����V��D�7L�`r����b�c��".�ZX�C��~� ��~F������H\��Eʌ��T@˘9�=eA�y����p�xơ]_wV�x���G=+��;�u�nɨ��3��U�2'�E�	 �E;��)�|U�5fU�#��K�0:�jj��%|���L�E;w�A��P&)>��w�l�iX�d�$R���>/݊ K�q�RE)#C�W�\\<�|��yx��>ѓ��V��f�f�X�5�u��5nBBͯ'"�k��1Dl*����;�����ι���ݝ����ް�)�5�@��7����\�|ȷy\�&����i�9�����ʎ�Аp��"�1[��H��J��E���h!۹���pq3?��~�|qz����t��1�Z�D�Sj2�x�꧀�	3���h������TZ�α!��7��矿��1I9\����u��<��x�����>C"grL���N�&Y���-b?��ES�՘"( :�s{h�B�^{�3�b�"����iNőý����C�K�PaW���_Q�?��F�� � R� H3蹹��0��[IUCLK�zb�:���s� H�n�^f���2���+��:�j 1�Ƙ�B,J�'P���_?���O6 8���������k%b�X�~Xv�	�Ri���--lR��E����[91M�l�GƟ1��X����\�����Wg�utB���"Z|)61ָ$��L,�ʐ�ay���f�mV������Re�b,Rbs����$˭���$���&��_w��qq���&��Xj��@O����l��8�s��$���8@^V�L���{������%�#�1A��y�OɦL�7H���7q�o,Y�~fe���>�+�(m8����qZ̕U��Ц1�d:�L�+���� ���~h�^+�$��D�^���h^�t�9��6��;��q'���a���vUc�6���Ѥ���Lz�:"�2�m��љ �}���ut��M�N�����]��Y$]\?���gp�)�S��X��ωg,�%��fŮ��Z��V�<޲�BBBJ��C�[�k��]��������ՅkgIԋ�~�ʆGΆ�*h}���&��M������( ���k7CNóy� ������yu���[�ɟ�JV��8�=u ���@J�'No�b[�o��j�s�#�D�V��j�&�Tq.1��ºw6#N>���mA q�o�^�N��rOw�r�"�;'PJ[9�K�.�{8��>�m&��z�Z|D4���� �O����W#邃 ~(?���>�&g�
	;wj,�~�:U� b�<I�A8�SW�~�gd����;4���Ш�Y`��H���/g�}�e�Z��p�O1��ߒ��ja_sZ9`XQȬ��84��������!*TunѬ�����-�lt�c�~�E���M|�ؿ��t���y�����Z�X��7� /4:��2�[OWu��Rl|)G�Q�8(��A�s"�/:_���K��~U�����=r~]������?q�ZTpJo�`�)}�{a=Ӌ�P���s���0L܎%�F:���C��$e��`aSO��j�è��X��ߍ�i�(O�^<�)��	��y��ڑ����m���G�`NX���1n=2��º�;e�$��N����������c'��Ŀ:fc������:<��d�E[X�/�0�`n���!;��9���$�����"��M�4���N�4�WS�o��
��(�r�)�R�	�f�Y;̏k��^)���^�.�'�#<�)#��}��B
�l1�yp�V�=�C�z�ǅz)j��?p��r�)��a�7�ȹ"����8ä�I��=�z6�hfHX�8�� _�.q����xdn����
I�K�wc{h��׈g�)l~ֵVe���t�9������z��N2̀�9?��/�g����=�
d��QX��z'�R����][�$��X�=��k��U,�~"��
�5�N;ڲm�ӝ.D�PQ�Gݠ���a�+���n��ۃz����!!�t�)�:��^��3
���kϒ�ω"(�zC.-��PU�g��*Wo�n��O�ut:A�'2�(�<�=������swd���'�ST�^�GJ��4������� ��ϬJk1�1Z)�*�g�kOZ^�B�����Ѱ䃘y���"��8�y�<�����؅��d�Z�4�/�كi2u���J;�C�ª�U
������[��W\�u�~���V(�w���AOA�i��������f�
Z����\U�*l��};C�U�sVYyĔ��u�;ӽ� #���+��Qz��^�J ٶU�o,�}C`�����A1c-T>��L Ɵ�������_m�=􁌻���T�5(G�*]�X�?�)�d���a�M9�c�z�x��j��޽�ȔaBݷ�A��o���F���K���0�<��u	O��ĉ���k�fc!j�]8�#k?��y�&g�m�O�%�2^cp��������ŋ4�9����6"��ӭ����Qv5<��n1�4�s:�au}}��]o׶Dtpwwn�]C��]����N	��������[p�`��{�W�U5SC�ݻ{�Zݽ�y@X����D��!ޚ��d#{kK���Td�ol;�d� �����#O�/W�h�k�����(���{MV����m9R����})O��SΑ/�7uV> �������EB���00�?u���ʆ	��p��P�ud,�P�l��~mq<�`��[7���HY`�0I���NQ`h��(({�Ȏ#~�ō�c�ۨ��󻇟&��zh���s�Y�`�}��;q�������#��=a��F�e���o�θ�e34}�4?�\0�����O�9�́��Q�������J��iY���\����_�Y�A��}��6=��op
��2�1���Y"e���Ss���i]lǝ=�l)�f\��7�i�_s�wUNC��dS�蔚ܿ�'#�YE*��YUnͼ;WgJ�JU��~t&¡u�[��!q�2ȫ���9�9~�_�-���z��`j9����PA��|��+V$N�rJD���A|�d�y�>O3L�+Û��Y}��q�g�M�[�k�5�o�r?ܒ5�O�Py;��R�[[/����(����f\�����َ3,��r\��m����� �Qo����?���9I�S����{�
��<� tG����]S
��R`y��7�K`QeM��"��?SDn:�J��}��>Gʌb�=�b�H��sΓ.���W
\�1	�_���Ɇ������=LF�����Vʚ������X3�%$%{��B�1�C�m���*���XO��d<^�w7KR%nvC��(�7F������.���ô@���>�J@�$$�|>�0c���H�&��3��4�$/<�A��"�(�&cը/���]eƅ���=���Σ� ��m�;���W]��������[� e_�{�]l'�u��Mgn�s���wJ.���w��nV}��w�=�Q�<(T׶;��9W�.�7���}
[�TI���U��u�R��s�����噫�t#w4	s~,�7}�� �?P��%o]���3/bWQ�}�Dqu&��U����$y�U��st�����U��/��J�6�=�/��0����\t�ȓ�v����ˉi�Q�շ�ɢ��}�[&>o��DV9�w�O�+���H���zS��\e�ݺ3B9����'�|Y��D�2 t�� ��-��#G��W�.P,�;�1�;`
�?�A�u%�'������+��M�}�c�}��J
H��������-�
n��]3]H�����s;�- "�����S��'��YMU�e5EUx�}�"٘�(�\qG|i�E�čv#Ӣ�" �u=߂	I>ɀ�ԧ�ާQ�Mÿ#��v�����!X�%��+�8�}������&��n��$�����ӓ��2-�mY��㨤(��RbvŬ�(����7O�[�����#H��z� ��9"�����3z��O��Ipol�����Ɠw;�vNf�曆�;	��Q��W�2~"M&@�Ǹh��f�&Q���-���{�b����¢�n��8�@,�s�r$�޾w��^vz�pals�r*�C�Sw�� ���U�Xɓ����z{��zZR����y�K�����|� U�������Cl:�5�32�f_#�w�`�$���}at߈w\�o���0&����̠l[Xn��f�> �B���QrA�P�c���bn ć~L3�~�#��7�鱕�`ii�8��9{�x��]��Q�Oߴk?�L˟ J��1YA5�Ү�+�+l+��)_��cG��0�*���jD���bO	�"�Q��7٭/�rG���JM�ir4=�C���4y�$�:+8ߞI����?˞a�ahq"5/�}-Qfs�^��*�l��؉^V�2�a������9��Nh]y����<=�o�����#H2�Xr}ge���;������&k�w�O�'e%�\P`P 2��ab�Қ��/w[��r�^�;�[�l���;��U��Q�;�Q(\�E�U}ϙ4��p�Ȏ�O����5����&#�.��,���Y;H���C�F|�0������e�0s�B�f��9�Vw(��`�1��'�A�n�S�Q��b�Av�m;�l��oh'�v��yЋ�9f����C��9	��b&j�!b��cq:��A��pr��� �ja�+W��/8^����_l�D`��yD:����M2ұ]E��ЎU��뛼�F��X�U�(ɿ�x��g���*�@�ͽ�����M-ͦi��
=��7�ꔹ^�I*[�K�,��k�X�����?̚��2������Fo>*--�DF���bp��i�LW�LW_Y����ߛ��Iג@��na�l�+V��jo���=:����`�(�)�Y&�=�ȿG]:�H͵�0�f��#����'.�c'V��K��! ZtL�'+䄃�t"Ҋ�N
��l?N�eD��
�c�&Ƣ�M���+>8sv[g�t4�}4Ӈ�j�&�ǵ�K07�WT��>��5�Ǡ��U���D�	��"W�c��y�� ��;^4p��v�ù9�7Fa/G���
�3ѧH�C�0��\������ɋ��{�n�輳�`s��%�������O�M'
�{"ߤN�d�bkr����&S^)�����q}�Aql�[�ȍ��^0Qڄg�?�i�O�����Р��%Ǫ9�k|ߚs\��!8�M,t�?c7!�~ۦ�zr�d�KI�R��We�w���4���^?i��H
9i�2�"�\���W��_�P�G���*<�_:��- ��$I�=�7b��M��*�}D��:l4x�{�K�%6��xh5r|'���2�g��7E�'H	k��b�5m�y�VMj)ws�0�� ��l�~d�âj�8��{"1��H�-�FaHD��_���᎖g�˩x�K_z���Nn9d�d־�lPr]�����3�0�!�Myܜ����`,�,{�f*#A���/%� �}��e�)�D� �H�}BuSR�����Y4Z�uOHo����6b��?�(gÐ^���_�j0���v�"e4ފs�Ys�ͪ�-g�����{CYI]�bc��2i��w�e�ǟ���!��F�������7š��۶�߀E
�#2����ߣ%����O!&'3�#}+ �UA�MMuHH4�ú��풳e��
�X�'.m:���4p�̻IBq	�����'� �$�UZH���VK��o'Vx>]7ڷ�~_�L�s�UY��x�N\x����+qY�
���{���5����xӼ9���]y��ѿ�X����L�m�+�o8J{�	Q �$���YA��|x������z`7��$s0�6�[�=ì̀Aa�Mt�R�x�*�!�;Î����L��"�Id���N��!G�ֆA�`G��Dc�������SGF3�U=(���b�6kMwV�M_���{ ���9,��j4̚a��E"��B� ��0��L_�N�S1���*=8D?�ӑ�}��x��|~._\�-Hٖ�m��+ω.�I_�UOf��ݙ-T��P*ѾD��&�{g������RF��Ѕ���ˉ��?�.��p8&�E9����<�!4�}l�7߬p֧^'R��"�5|B0H��9
�/�Il�6(!XZ�Y*d潱V&N�@���`G̱e)�ʌ��R>hLf-:������l`[c%��ĥ�5���Nk)d��J���#b�?R�q���&x	�fxrJ~k0gq���xw��q�TL�ψ�Z� ]�t��gV/a(@b|Ӆ6�$�dm��m�x�#��h�4)·�ɣ��N>��)��,�=��- ���g!P��x+%n�V<��qPv����e{���^���CkØ�f����0�t�$/IfF��'�ҝ@���g��	�ˌc΢��`�|���7���ǲ`���J��+��m�n0���O�9�@��H9)E!u������_��6ÂȬgIO�n�үΧg��m.X��Zl�bO|�Lfh�(Ͱ(�����JK���V`l>�W����j��G��w��7]��mV�q�N���Y;�4�Ղ�p�=���)�������?N�cbd��1�WZ�O4�N�������k���b������]����n��8_3+�mabp8��\�OY��@���o�T���蟞WR�nj��|!*~�yT,������ζvANv��jC.�yYz�D�,�����:~�6k`R0A��u�-�K
PNB$%.2��>�!nP��Ӵ���wB�h�<+���mZ9�@{�<��Ds����Z�6z����}�X��u��:������PI����|M�?ʹX�J�iI�"��ſO��r�w�9�K����ws'�O��$�ڭ�D9n�n3�%�V|��V\4�mO������kJ@b�J�e_
<����X�����F��P�
0,6~�D�l��� r�L��sYAU%�� �}�h�	!g�ɦi?QD��Μ{W�#��2
e�9�|5x������9��j�V����s�j;Y4�֊f���'!� j���G���b%e�5D8�u�UOPUԊ �����I��F�wz��ЉCv[Y#��
�$���6�k����㶷2�����ovB�-�o 	[*�߶N��/�uEOy�u��禑V�u7�v�˟�9fy�S~����"I�>� �7��P;��>c�w8����K�	p�]�̸S���6�����ȣ����䜃�2V��f��ࡏ"!j��R�V9���t���[א�p��V���^n|~�LZZH� ��Ǭ8-������zU29[$a[ET!,�G8����ec���r�M��DP.�"0��7Q���"�Y$��H/"b���N@X�-�J�w����Xv�Ǐ�(�L�����u:>R���$�k%p�T�}�����s_�]|��q�l����qr4�������s��%�r���D��猾V"��nʘ.Qk߯��ܹCʤ�;����p���Ws���h�ى�YSx��[�l�?��Ln���rڮj���sB�F���3���_�Go#�y�6�%FcH�9���m�
E@�O��1N��k��C������2��X,��ܮ������7��ſM��y,5{!���.%k��a�W��	�7��@��`t�U�z��z�¿U^���k�2�v���6��#�~� �k��b#y�yRr�� �?Y�gOs�m�T~**q��{�i���-����\�	6�Tܵħ�}4@�����z�db�g�����t�����jI� +0���wtu�D}5n��Ql����G�5�y�M<��!�����ڱH7�����i�����?�~�j'�2���V\f����� �T%s^ne�)���U���	�U׷���	�8Ĳ���3���`�"�h���vāΝ%��%�2�7�6D�hc�z3]
�:$����1��:�s&�~�O��~���i�[/A�}��Hs#8�n݊��q��[��D>>�5)#��MR��q�Lשmj2��X�5x5&��F����,��L��҇�R�$�V�V[v�e���N	i�+.�>~�x�ѐ]ѽr����� ��Ұ����l'�Vo��k��Z+��(�]�U� xL���Pf�Ra��W��ͧ|\>��=f�EWJe ��Te�M`�z���+����|�W7����p�F�l�^E�Q~9J��s�V5��}�C#���a��;{o p�{o��a�a,gl|j�#�Ù8��R ˦��)������u�c�7ݕ-	��+�e�)~�ÉOe��
�55�>hU��e��9�;E�VYy�A\ϞX���W8O�nOAZ�ߣ�%�����ľ�iG���p9��B�'ٵ���Hz����O�gi0�1�=�r>�W/�b�q�C��_k�$8�9$��2�; @Տ�A�����x13�u�>�c�&��UG2�����$ݫcs��<!���5<����h�MK �2�~�h͔"%��H���0����ƒ��B)��88�IL�A��$EE�s���2��.�=+D�.�߳������uI4��j[|�>�Qt�}���'ܮ��KG���W[;X����V#� bh=̭S$^l|�c�|Ug|�?]����	DǱ��U�D-�*3F}�?���Q8�aYQ���n]��Л�d%T>��z;t|Vj����\�nф������j�$Xʛ"�ġ����,;݄�o���5:gto���&t����TBu4�l�Dn#[L�EނP�
�Kh�a@���_���"�<�!ZZZ22�~���#"�	�Y%T�^����F��]^�/�t�>��'��0Y׀H������P�T�Xآ8�ȏ����"�/�?��6�����gQ�@�@�3�88�sr��{o\��@L�ZO�d���W��T��I<��1|�Ε��5����a��#(���ܲ�vo�8��3O�)2�r�i=�7v�d�Ɣ����cƮ��ٜ�JC���� �����N���>�mv"�'�lE���j	���#�vn�0��u�Q��x�:�mW,�"�Z��Ыm�ViKoֺ�����.r�1""nC�G�F�0�f78WKX�d�W}%�(*^Y=/��u�.)����\m��@.AM7�Tn%VLJ�_��ɤ̖W�1Z� �c���rja���'e��ffwUו@5$i�T�~�M�>ܬ�u�]����Щq��̌ƞN�J��W�Ŋ�T�RZ�ڐQ)�;^�~��8Ckh�"ĨZ��l
BB����7��3h�|7��8��)��k��7�����R�z|2j80�&����
���J�0bP��.Z��	�-��z�o��0��	���c�p����J,�%Z>���-�b�9�S`6��D��#鉤_?$�����e��R����w��6�a<}���d�b�1{�wk�$CT�����Q�����s�oY�p�N�n�~i��7#{�<�/�ca��L���k�g8�a�!U_��T�ސ���ЉW[Tc ����bP��䄭���
��0U� -u�.�Uk�u����R�S}>�p�&a�FW�>+�cp�GO��qS"i!����L4��M�G#>��N�X�`/�NE�/����*!K`l�Fu� �r-�\����|�ϧst�kD����������}�>]����I���BkЄM}!L���>/-u!���o�fUŠi�����l!����
6�����c�L��ȶ��yUI0�S�5�(�@�	b~}��+%���D>��+��2[�Xvr<��xC�����&�
������_��6~���x5��v��qc�n�p��N[�8H�%��"Qԭ*r�(a�j����z�CX�`N�7�lt��_��2u��ÂΣU�� S��]KB����괆f�߻L�Si��ᄩcV�y-H�3���ɦp��a$$��MGN��{�$0��oFƧ�bz��]?���9� ���@�[NɋV�m�����|O8m�:7&�@���I��(�l�Di){q���_E;)b�H<��O�Ej_�Ʃ&_�Mx��n[����е��s4Z�>z2-N�F�P	��Ǿ�#�[�N�5��t�/*�9q]!Z�<}�~������T��|h��k���T�!�??�pm�R�
�\b�I���!R��`
�d��!R��w�8 !����3�[���ZR�3KnLU_G�B�4�;�l̳��=1F)�c'�_��g��Y� ��Hk���6�H�S���H��r�%� q���aQ������g�v�w-��bN��w�,�7e2ِ˔Q��ľ�.)�B_�����pI�;�����ɡ`C�SR�σu���L�b1L V��4L�2v<�������jv�AWh�F{�wGf�_�Db'�Q`1ZM�O�?�����&�1+��,��X�;Y��e��?�"$�RY��i!�6��Fm� .�l��4E7�xAy�����2��$tt���kL��}��֞����3{�TCOv�3��cS/���k7���'��G<�+�Nꇅ�;,����S_��%,I
���~R�_}��UԻ'�WDϔ��v/��T�H�k��ZTv�D�h��dZ̑���/��t.k�,����Z ��j��#�pn���v����y~��<�-�+�J@Rw��a���N}��a���:HKS�,�#��[x	$Ҿ�	ϸy "���w��wJ�
�c�#�3R|�]��Jj	��|�����º\����TR��ݝB1� A=��-�!�w��W���R=��\3�=x
P_w.q�X�����tvi�ſ1$��wF5LVsdੱ/�~ºt����̜m{N<�K�IXFv���R����lܫ傖W�2f�H,���v$W.���ͨ�%�|�W'2J�x���[��Cyo���mYNf���يP��V1|B�Qn�{�� �ˇ.1o[Xv�La!�Nlp���y���Y·YG��; �X�Ӯ��__>+�Ὅ�N$l�L��(��N���室�񪍚�����kb�B����vlI�4j>�Sp�5�A=DʭD��ƛY�����ϒ�V��Z���Foy�xA2�
�雞Q�0�N}�z�ش4��)h�����+;҅J.$b����Ũ�U���撃����z��s��3~�����{
2��Z�G��>EN�?�ݟ�Y���'m�Wދ<��a U���'AA������[s=9�F�wLQ����MP�M�񻪀�T8������Μ&��`���k٭m|O��:�"I���7JXA��k��&��#�&ex�2��l�/3g$�drU.�f���P��������~�!ɮ`�j�~����ƙ����4�O�e:,�{�,2��_//G�52��F���7r��R6 �z%��}�1�v�;,ڰ�q�sS^WTc��R���-s&��G�&�Lɻ+3�5���r����Φ��7�P力ι%ޠ��	"S�O�A�q�ۑ<��U������ ,%#!�c�|E�.KM[>�m��f�*yvv-�A#�.;�	G�"*j13��GI���ɵ9�
`�R��P,�5=<�z���)s���o}�h�����o�êFB'N�=K�T&r�R��p�Jr��>��[�D��>,���ƣ�/գP&��c^k�	��C�ߑ��\�q��С���Q��-��h��Qo-�yY��
EW�ȱ���T^�alF�}��C1O��rM��u�8�:�z#�a.+H����
�y��(.��V���?��I��H���G/I�xB���caI��0[����t��N�WWϽ��͘FL4���Ť�3c��Q�z Qn}{]Y��˓����8Q��(g�.H�9�rSfXҝ݀���>�۪�\d<|ըn�I�����p���Wt���vM1�@������%������+���	*��I�Q�(8>(Gr)~����W�;	IpR��5�����BRUS�`!���?�|�.�#f��cn{.�y>8u����Z�` �ts���6^@)�U]�V`iI%�ʐ_S������uC���-�v�ߞ'YMW j-ty�~@�׮VIW �o�ټ�� �,gb�鞠�s[��(9W���^�d�$�ǩ#c��_f��uB��0�I�1h ��4~|�j^16��H>�ʋ��J"�<!�t�5�쨧?L� �G�k�z�Uw��ҩ���*D�����I[��$-��(�������֏R`˽���1VV�ފ��7f��\��[�s�[��X #�B}5��`��{9y���EW� _:G�w�%���T�2I[K����b�
{8��yv�ǒ�8|z�9����x[7��yO���(�r%q�u��=B*����g��H����X�5�UE��g2�OI���&0%��^��Z[z�D��+X��U��G�$�����^5��:��KS:J2���̥D�M�+��q<|�I�d�Cl�a�����{�_��k�r�oPd��B�T��3Y��Hn�2ޑT�~��M���,��XV�}�ֶ�!�l4��b��4��R� ��]�;ߐ���>YJh�/����˔4#n����G���x��E��0�얟Qã[�����Rx����<���	w���6��e��Q���G���º�apX\� myy�C��њ��h���������y9��Xh&��:]�!�`�Vͮ;M��C�W�ؔ��s{[>���'z`��U���U^+��n��4"x���X�*���~�.�xP��y��M~�[��2�J��Wm�2�/J�k�OW�	r�"W�P\�^���x�(�&3K�8}
6��:��Y���Q�|~' ��=7��
�\?�������>���ٍ����X��[,��P+�a��O�݉ȡ�C�W#3�8c�w<ͦ�.їV�r���[��1�;�S�������%�ߦ�wbk�~�X�ω6EEh��3{�d�O�	�e+ui�D�G
���� v>]7��[NI�ک}=���^4>*!�����p�rv�L���[G򤢟(�%���d��|ص���mh|+@C6CG�Vש����������_��߶2%T�ld@����tg��*ÿL^��[�o�.�UtG�����Ȗ�,�;�FɈ8=�C�Ay-�����Nz���B`��~� {�Z	������M��T��%�>������g���R�V��Ɔ����P�p���SѨ��hH�@q�ᩃ�E����8�o͔��FٻZe��m\�#��;�b/z%�]ުq��xu��o��o�;��ؒ0M+=�M?b��&+8��ֲ�S����W� �%(˪�������<O��Þ*$㭝���ď͔M#q�,mR�Я�Z!KR�R�gȠC1��r]��ya�&Î*k��1�lӹY�WY���)
��K!'
[s@�6��Yo�+;l�)(��G�1��;h�T�0�j�C���_k��~?+2�@ �$a< ,�������s�����J,�r&[��f���Ñ���J��+��#��zF��~~"B,�O�:��SV	�"7��xv���.�i��?�q-�������\G����,���g� �on�of]� \j��Z0�{���N'�����w����w�.��PPΑ����^Rd��q�P�M��H�)Ms�%L��ڪ��噵k.w����~f�WVWT�7��χ�O���aI��B�4��%ޘ@]�-��|��]v�ں53��DJ
B�燵[�ԡ��!+%�6�'�����XT���5��[�ҙ�Z:׬t"x�5��R���JϳkG���X}ɻ�	���H&���N�n�Ʊ����A����ٍ˩��}Zn?��w�7��`4�i��4G����|��q�B㟧5�滅��&;�j�֘�\[���Z���P�t�L���s#�OI��s�^(+�VA\R�q)fY��vZ��>�y����Z���'��n��I�y�zW�5?]{	Tu�C�����M=��=�k�H�0�R�+~˱����nb�X���JE�CzrJ�s5�7�eaa�m�ǲOl����T"���B��{J�&³<x��O�Ft���ƭ�ϳX�S�U����"q�6(�zhfZ_�lR��z'ab���~��s6������.E#�9a�S�����W�>kj0�1T�Nep�t���B�����C�&B�̖�$�~��gs���!|��$n���ihm� 1�)jg����&�/��#�l�����L���B>f�x^ӛ��� �k
�i��>3��w�:��?[@�^�؇<||�0c
НR�|d:���X�Dڷ���	-�p�t���&~99y	g�jϏ�ZZ�K�b>�/��^�RosO��gB5.�ם�wwkJ�8� g$w��~��j.��Lx�>�͒��hl�����S�W;�vz�C§հ�?J�D�!KI�L�0&�`[-�:/�9��1�������V+�R�vT����u��3bN;���&��iE��WQ[�X�§6[ 3��a�8�nc��,�!	���:���?z7�*d.��}�=Y&�7B����i�d�3"d�AZ��#'��S�/^��]3gL��	����-8I/Ư W�}�h��G�+��]��}��m�>�sr㏀���>D <66�Mg;���é`�FtP	��N��"�{F���bRu�+�3�q��l6�oY�� �L�p�y�,'��MJ|��]u�m�����|����کF+�񋈩p<�]{uMO2�ǁU�0E��l&Wl��&��%i�!k��e��������|�S�]>6M�v�YK)	�n�ڌ�wmmP�X��i���g������pլ���[�'�JZw��.�˸M\jVE��r�΍�^�t���EÂN��pn�ح���9�.h
�Ni2�F!O�������8��f��@id�wHI�V$�Ңg�C���[;�rHUhL`��Z��mÉ��ur^�K Z>=?�	Z�z�<���`&�I�~�E��X*3��O�/U�����r%*�?1��+�7	�O{�_��i��1������}d�U"�5_:ε�vωvQAd*�G�%�<vF7��ؐœ��yA{���c���e���
��k'fe>]3����1!sg�����#lF�
%.��b����N�����?�("�΋�gT?���v�7H=v�#緉J��Z<��[����v�H��hd��RĕKh�՟�u5�J����3����Α�2�@�{w$��fN���8�B�8n"T�e�����zo�⪊�X�C+�����а�EDr%	*��Lލ�t	
**x�I����i���,V�^ɣ����A'm�8�lr �PIjUdJ;�����tt.GM�/P�j�����lH�Ҝ���%�yv�����7�i�5��'��?׎�X�i2��Ll�F=��6�@����Yg�C<��$�p��b���*�yY��'�k�?D�E��s	��y|�rjt2X+��S%�z>R�1Po�sB���k%O(ì���C�P���v(�u��*�w�r��
YcY��2"
2LF� T�1�\�5D�k��0\n���d���I�����u�8��Q��Ɠ�PPv�8�	G끝��h�s��:�vF�S��{UJx��tg������dP_��Io&����o:���������H���r�M��n��-����۵#s�0��M���L&kw���q�Z4L_aX�e����!�e���D�0�<�#g�#u�!��|����Ň����6n[�+r�~�(>Cl�a��a`p�T�|�Fx1fq�	o[�Ĥ��ͱ����Uk��G�{vhr{}k�S�;�ap�?����ڶ:������VG�
���>��"Z��t#@��ز�':Zy�s�U��'��L���ȣ��R}/�G_V�P�F�e��VR$���V%f`wU��z��=�ЅD�������~����~c,̂W�R�����)�D��>2u����O�92�`�{J�#�"��1��\G�>�oP���I�1C��%0���7�)��QE2[����{��~�z�Ƀ	����g�wT�G-��rr�ޖ:���)=�z��5$k�,��GKo«W)�%u|mC{������ 
???`����e�����[�Z�C����;���Mr�3��R�ݸ67�-��ї(��W�j���R&֍��/H�6$��8X��y����"�Rշ����k��gk��6$A�uKk�X���-����Lw�u���Z�2�m�}���$����]T}DЉP�8����_�8o��_�m/�����kŭe�U��̺�D��M&�x:=��Et���_o��� W�fU���*�_��H:lľ����o��`�|�R�\�O��`SCVe�
��[W�O�\ф�cK&8��<},����a��ֆ9�)���t��;,U�n:�Ԓ�C=v*,�1A��+�q��O�nM�~C���:O!�m-�PcH%C[�m�rh5�q�Ow�u�S�N��#l��S�����pYq���.5�$v���6S�����'.�s����O��.�	�����y!��O�?nv"��<�k�H�I��8�+������=B���s��c��:,�~C�^��lo��	bw�$�n���IzA3�o�2	^'7�~��E�F�G]c.��A�rB��ܛ_���/W$���|��^s�k[}���\_zk^9�1,>��jߩZ��S�d�0��8`z��S__?����*�?��E�N8����+���K�Q&��m��nO��`/�eFd�įi���nk�s��!���כ7ĨW�[+����M���K;^X��+A�����]�MV�����/�f#
Mͺ�gR�^��!�fT!�s��q�?-�3�S7i���M���� ���,U�ΩP�"qib����c�J��_���`gGL�(���u�j񸾾�\�}Fm_���� {�0��pd��်�B�VSՈ��I�3�:i�������<~���}b-~��ݴA�@���l GMWnU�=��û���,����pn����Z��O�#>�p0[p�7��1��b����Pf�԰N�q�鴤�#��f�W�\"��y��Ȼ�3�)4r���"�P`y�R�ٜ�3�(�w�w���D���A]�k�X^�-�~��(N���H�����I-+Fg�(��
)���_�;�!/h�%�N��&=�9Y:�k�?�.t_�CQd�C�m�H\�G��`�+�Z�pw�m#�����V�c����y����hȡ'�#�[Wv��`�G��Ko�$u�CJ��KV��S���O���~.��fr���MOi��Y��{��H�	�Q&M�����B�pL�R8lox�Mq�%�L�/�����"���m��?�o<��2d�Gͅ��\@(h�ޓ��1\����$ �m��+Z���ͧ�OX@�;�rmZ�R�&���V��m:=��~!��Dm���L�?X�k~������Bu�]�;��;&��C�2���F���11%	��ȡ{�)��h�/4�W�\bw�����Z�6�:��Bn�đV�� ���N��
�Û�Zy�9sI��	��5�hz~������\�N�g1��k�T�қ�x%x��9���U��kv����W�������q�p�:#�<Ƽ~}��fs��4���P��ͭ_���n��� {��+F�B1\��f��="�˸��x�h�9�\&dJ�/�6� �K�����7�*�L��/rB�$E�&��	��N�[�i�{�m�k�G̗���2٠�72��m���z>�fx�7�n9��W��k4tI/�Yha�z����Ybdff�������E���A�2����cV� ��<�_�K~6���/Y�V�V|��,����n�m���n=�����"{��#]l��qI��)`�ܘ]��Z�7�Qstv�ђ��Vن�+,���(�D����M�2�k����^���
�������A�3���e��WpMG�)�,�U_?�ܨ 8�*o�_�=�B_���Gw����v����s��&���sX�I����є�}~�P��l��m+��'�|�^	��==����ཀྵd/��<׸q�m_%�����zV_O��٪nU�mƸ'�۩n6W�;Ds=f��79q+�ݣ;x���K�f��-�Pس���A,����Z���e�\ O�nb�
�fNr�}W�� s���2���������P,�
��%TX&�ЈvQ�J�gX�'"��ǍRm�:�E���;˶���d�֫t/k���<�������$@��|]S�����E�
�����Ro��Ƥ]�w���%9i�r�~_b-��!�q�5�)�b
�D.��Ñ�ԁ���q���B�ҜCuKfM���2z�ť�!�
���>�z�|\�IV��Y�mB����8�Uq�-?��Qϔ��}Ȧ6�@'��!;��J�C��Mn�;pvwr)�ܾ�uWWc,�3LTY���G	d����%ť/#w�PYSm��h}ca�E����C9$d=ga����[҆�[��2�,g�ce�E^�|]��7Ox�)R��7��/|��M�DS~ڶL�7O�#$"|�>����a��Ų=]���~FcGiim�W��V=���@V��v Q���;�8+�4�Q�ޠ��t�hfR���G�`��X��@���*F�2���|NP�$�f�;f H!���Vh����H����{
���uQ��o��)'�-\��_��X��+�(��E�Iפ)��ɕ �?TO�\�NI[�[Q�ϡ�`�N,0�����r�f2��S�jO���L3M6l�
�6:� ����6���V�X�*I�����[�)�٣Y�e�� �;0n=��}��
�˘6,<�]�;b��H�2��ᦦ�ݫ�o<?�Vg.���q��2��������a蘆�(��8���1��jzU��s��(�ɅI�샎�8[��G�Ml������E[2!%� Oi�4L�������6/�T��*bB@mSV����Z�C�]#.Z��%�Mf�3��f�V�����x�����Y�s!]�8M����IM^$���J,$�7��B���@%%[��屢B�>?[�G�Qh>u��=�ǎr���do�V�]{j�GI��eIQ�Nŷ�y�(�0��Њ(�v��\,oބ��\�͛�j�6��Ua����O�����X�İ��!�|�w�|l��(^�ѷ_�AENv���P^��7��'&����#�^.��g�n���ڿc2~������ssFZ���6}�ٻ�_��I���ZgQA�3�Q������� l���>T/�t��E�[չ-m����[pw'�܃���{�!@�@pw����q�y���;_������^ݏt�Z;m�;a�12*2p$Nc&UsD�U�(�7�U*#1�!�L���4]�����u��Ni����i��|���z<{��i9��BD�;�Y1g$/?d��vՈ<Aa�R�@p��_�}���j0�L�p�o�jHz�w�����1��y�Q�͢���D�2�����յ�+�ʵ,3y=@�K �d��e��gr�ou�	���|��T޹Tl���-����2ڮ�U��-�I�y h��;��P�6z�7�۫�&���D�6��r��q����E~�~ 7qf9�KL
&}�E�R��y���~;����G�>�E?�0�]�����P��O�	�� �$$[��}}	B+���qA/��{E���^�*#ėA���B*:lx��(�_�F�d�s ����c�xl]�P���io�o�4��V�/���\�����Y)�ə�Ѧ����t�|�o�p���8����ww=��Y�pih���&��Q#}����ͻz(;��3�N����m~�����\˧�u�2��a��v��h����4������������*�z·.�������6C4��r~�ٙcF<�����>��Q^���������1���Z��J�_��
hfqq��
���Q��Y-n�x�K@4�0w~�r0�_��`��#_d)�/�$�"���ԩe�<�������wcHnW�2)*
bx�|����$ͳ����n(���Q_z��������Y~M�e_�����(?�ď���e=P���q��:�j4�J��F�k_*dEiZ�Zx}(��16p.�������>�{��ys���V��蔊������S��&�e�7����Y<���kO��zB���V-���>���Zۥ:O��=�̊����"��0㋓C4��h8���fL{G\L�|5	'��wg�yuV�ajV���7<ϥ�-��+�<���k4�6G��^����p��+���S�f����,տ;Y;�,��叿[@�ؤ$�
�n�ё����pws7�~��@��8�K�3�X�ޢNۢ��X�w�)>x�Riy6�=5H�n�g�[o�@����Ϣ���H���hW��Z��yҍ��E�Ҧ-�*�㨭��y2�%voTQr���@�/���������0�.���Ɵ�=�c�]I��<d�(����ot<�ȷ�&��i���i��U�����A�+P�f=æ��<17�&z;��4��NFה�>Ac�vqqY���Y����+���/,����8���f}��R8~�)��+%����A�Ǉ){�C��24?�@�;!�#+G�}"�K���nn�����J�VTE�~!�h�y5t�̊l�R�ܳ?5�c�A�#`�l�N03|���W����x�5�{f�|�R�-/ûr�T��:{`k����nV����0���i���Z����g�r��|�c�&S��Y����}�2?��T���v��*���m�W��l-L� d4�V�x�ɛ,��3`\0k��?;B��оA�%�����
����&Q��X�P2�mW%אc+�������D�^]t����5���`�;�@�55�f#�꽽c�s�J%�ޖ��}�~o�!R��wO���������ʱ�,o$C?W�3�'��;=|�U�-��	��Ax��/&�Ҋ����?8n�iDQ�u�neU/������
+���g��'*#% uAk�ŗ0�D��؇�=����ڷ;�FoMF\o�&���@�ΡuG !��~6Uΰa��)o(���mΝr��C�0�d�����S<_�!�w�ր�g�ׇ�����|$x\��nǻԍ�7?H��ME��G7�'��0C%��w[G,̻���OOz��I�إRf��pN⏱�i9hRh[���DP�~MިQ��$k,,,b
N���g�>�^�飯u����z���9Y�yQ����m��ң�fܻ�Q_\�v��N���f�=�ӕ�l[n`�0�+�c=쿅���H�qֻ��iF��z��`����̂^�$]`Z��!��{Hv��b)�4�HB��>�ZS|�8ĄX���Yt������4�i4�.-����u<�j�1�	t'�$[q��l���e���-�i,�5��~+)���	SXR�a��[<-^�E"��ǹ}����vy����ְ�ŵ0����7��������`oc3&Sި~�B�S�GWR��9�P���R��N����*��
��/�C�orB�^�i���ͪ��/.���jp0ؓ����f����ʝ�������Nly:�+����6�.C,���!��/S�O�O���N�쒩k�Pϭ���&�����7�8cq�����O��	��e�Y�?D�ġ�׽Z}ܪL��زZ���7���+���Q���B3�?�������@當���/�4����͔�U�>VP[Gſ�`�ǣ��~�IOe��/,oܤr�x����	��g���}�h��YKh(B�:��l�Kr����+��1����.�\��� ½���s��#Hߛ �um�O�)&�R#���b��[f!��/[�q�?5H�C#��4u����^t��t�<�ݯr���k�IN9}�W������P�@;|��a�������b�����f�X	KD��t�e5d������),�}���{���^B��xm�~�;X���2�.�Է���}�^���>|@燎N���H`=}Hspb�����I$\�*�����1>}T-���ҵ �`8�mW�n{���7�x67T^�7��o�A��%���zx��� ��CU9Е��s�i�qK�V��}F�F�[��� ^�̏o�D]�����c���k7�	h�_�(�}�p��o+����>�_�>@�q-Np4h(���A��?��?���lc��Þ�ã�AtM�@��w�fq��� �M|FW�@�E-7�A*��������#������$��ߨ��%�6.����&�C�����q��V�7�6s�3ݠ��F��I����[o"E���fu�;�UM�b���ʅ��M�=Z��S(Ivvj���É䛛�F3j��Ń/��
%���{G�IG(����e�l��N�-Q��dC���]���D���H�,\V�앫{/����W�ᨨ�S��/FN�=�s�Lt��s;/��<�NyiaQ�ِ��퐪��AW=�F#�:�S+1EW4,�M�y�qz�$m��0��ϐ��=��RR��iB�o���>_s��X��R��[?�no�|���T��:�F��q�p
ͪ%Ϸͭͅ5/xx�<p447���OS��S�^y.��b��k�H���j_CB�������d�\�o��n�~�Ct�t��Ġ���?O�Q�\�#I��YX�=���/@�ا����p���R}����s��ۦ��	�$i�P����][�/F�=���p\o(��Y��5����jUs�������j�����q�΋����G�����M��%�nT�"ʁ�`�q�.�L^/(ڸ�T+;W��c1""b�I�(-f�*(T�NA��J�y�s{��G�a��J(<b�{�f�k�K[�!jB&*2�ElA�@�^�E��&zZ�i�A B��:�U W�-��l�f6����P�.UU՟mm�((B�)����X�>|�F��^��W
D=S|,_���'�E)�#2�t2��vf\@��øJ{Hc{�.v��L8-%U��Yc7¾L8�hU�A�9@ߟ�ȯ����2��uS��,z�M�oư?�JW�	ڀ�$���q�~I���@���@�+���`���~#��^��`,�����v9(�l4�![k1��%�H[��Y_	4�/8�S.�z8��T����M+·���.v�p���7�gZ�9��v]�RR]�V�Б%�G�~:���Pһ�X��p�~)�hjJ����
o��+�e͍r��Lj�OhU�w�:
a̰�/�������j�o��R9�~��w������I��a��Ì�ԏ/�	����KsO��EiX�&lk���w؏=�j��1�9�Ne�W�gq�3��b����Ǵ�1�䕥cb*(!|�MMwT pf���޽]��SYPF�[�z�G�c�Ϩ}��P\�{�s'�'����a8�����V�f�3Lt�8��ܵ5�}!n�(��9Vg��WK娱+�G�aq@E95���m�e�|ϲ������ŧ���@j^꘰��ŷ+�5���3oF�7��-7��B�@��E$A~�%���oH�tҺ�c
b[�L�-��p������bm�?����n/�XZ�=|���?n��T��_���݋�M�1�[����B��(���%d̋S��3aeu@��
۾��z��1�P�L�tn�Zda����\^Ӥ�h%��l9�v��1��w�����CE��N���f�a���}_��?�/��+�}6�/�[[F��/Rt��:І$��56�UU��.��˫r��}�����'��5��\Њ���LM6!���a-#]��t�í*	"B*��Ri�=;�ߝG�fS'>�*����M��o'Z��HEwTTɴ羾Y��2D���L��ڝ��ly����ޢ���'��Fr�쀰�F.c�!�A�ꮭb� 9�g~����`0&��������G+t��]a6ߕ����p�w��0f�@ɬ�����P%��i�NNm|��G�������Tt����8$�{�n߽6�A�sIe%Z0,*?�DP��������^���}�p��;L��'8�LrC��+Hpl/�?Mœ���lH�ԙ}Vth����s�l0����z�^���λI��5<!тT�����褚�
r�u��H�z8�_�y���Cr�KX�P���l?�����0S/���-�2]^\�B���<�ό%%U�E
٢gUƼY���	�͛�_vs��3�B�Y�	
?��;��lƤ �$�6�X/̟�� ee��U��\��X�����&��$�����]���-m"8X3����� ������ ~�:V�i�#S�6>+xz[Eu����F5a���}��1��|�I�������1�m���B�N�F�Ht��M��Ҭ���3���Z�������ć�{�qW�#�[���i�,U�>�����vߋ3·�/�F�\\jj�N�����۴��M��e:�*��u�K9^.���/?>Ѫ<�ƩW�f��$J��4�p/2�����?��!z����qx�v��u���.��!z;� ��\S�ǐA�vv��2��4���ʭ��Bmrg
za�
^��c�b�׎2�����y9�%w�!I�·�F��G����O����i�p�s�r����ʭcD�Jͭrq�Kڅ2H�HӁUY��wt���]]^���O̻�|��v���9׃N���_�%Β�Ia�g����.�.12^�"�}I�<��ڈ@���dy�l�.4yT���e�0bt#��Vܱv[���N������6m쓸�Lh@��z��_�5�:�(�۸�D%���Q��<��T�B���nFJZNALӃj��q,k�ǳC���<+g�y��y$gG�����gf�e�NÌ��fs��"fw�\w��D�=��|�.�X~ofe&�4�n�½��us0�+{Fd�WX����^ٟ��@��x| ����'Q%�=&��D��4�Ͼj
{�9"���3�˫��:H'G�+}��T���w�q��X�7����'����t�	�B}��&�<�{!srkJ�S�Sal�
=�4<��ٍ�wf`a	_
���&�K�@}K怼�(Z(`��nh�9�f˭J:dȲ46-�F�6X������__:-�m��Ԩ�����z��AȌ���64Q2�ܬ�ح'�}�挟�9=tW-E�/�7��u�QY�ʹ�6Q�v)BOO��y�����i�ԗ�3��t�����k�����H�b�Y�����+��Q_pDs��q�����v)Il��M��mV�K,1�)��7��xɞ�#�Z}��'������F��?��L%ok��W�U蓋K�ba�
9����MpK�������φ8��ܒ���:��%?v���-3����_�iJ8 ���ԍ�[&b��j�)i�X�Q_�q�ZҶ7#{�J�mxo�r�z�,4�B�ȏA���fN�F��� *�1k�����E�޺���m=�2-GǪ�����W����\GNV�/��e!r3;U�gӏy�A�/�e$}և:��@�	�!�/��w$��KAן�&v_� &�FZl����\���/���h'�9g?��f:'B;�h����S�*�}-�T9�4 ����zBqш��\� }�'���q�K��NP8C�<\F��,���Ǝ��w���^:�:�Ƌ��C�!���L�CC��K,�	�R�N�!F�"a�U�h��-�6&�ơ�s��v�l�����Mo��0�s�=,�_%�B�|�ڋ즒X"���MkUM�4H��^�i��8�<lZ�>�-�u�L&"bI�=ƷoU6�^6���
����s�.�Ņ�94У(�s���ike��o�C�⹢o�C�
�>�F��i��;;H ����S��5������A����4�3����yH1W����:�����\�"C{�&D��BB@���b��_ŗ��|���v����G�1���S���|6�\s� Ԉ�����V����0
&��A��5��+�Ze�!��!�L�E��Gmh�.e�,4���Q9
����cyb��幑S_��3���D��+uf��d+..�@Xy���'@�hA��<���_��={@	��-��w�ǋ���"8:v����KWRu˃�����YzxPt������mW�e��~i+�Iȏ����g�����E���\p@��@G��a�Ј�757�ٕM�|YZ^�9;��#¢#��&V06695��β����,R�;��,�6�j\��̿=��5l7����X�`3�8���j�L��-���I���Q�(�q�;��P��~��'���\h�V 6� $E"��NPr��Gpb�V:����Wv��
>Y���񗹾"E��I����7R��!�v~�q,�p,e�5� �~D0�[*t	M��G����6���2����ĺ6�
E�4��bɼ+?9�夰��>�O�
�/ϼ��Ǜ��{
�T9̨?(C���-�n�B!�o��byW`�!��q�������Y���X��|YJ��ߐV���#ַo�F��ٖ��͆��Pbc�bm��50q�E��DѴ֪��[��ۭ��~K�I���1%w�V�bJ��z�rX��sC�K�:�S(M���)eHBv>l�������̇\�J�Ùǈ��������/���d]	������� |Z������	G=HS)��������
C� *�F��=��kB����%DT������ ���y[V�����q
w\I���3��N�E�֌fj:y���$�?�R~~����/Ed�K("ʘsM>Q�L���_��½6�}���P.�"����|� ̔۾d��ZEu�A�����>˔�bTW�}!y�c4LJ��>�v���uw���t��(�����a�����OW ��<s������� �˱�A|�d����V��W�C���f,S���W��˩����z�P���B!�fM��:�ȷXJ�4^�ˏ�?\�D�X�8�ȅ���w�@�H��� 4S�n��8��awa��ȵ��_nS\��6�꼉q��h�ؒ/ޤkr�)�S��P���{��껖$R��PJZ_��#v`r��&D�?H��uې�
rO�{��ז��_f&�`����B��ͤ�X��RG	�#8������MM�q���i;SZ�I��M��W0I���Õ���O���7p��}�����D'/�Ϧ��״X�Ɣ��\�������(�s�|\�Qݥ�����U&1U*?;BCA��L���ೀ(�@0g�`��0��_����=�x�Ilѳ��,-�L��6���H��������Q5����*�_�����|�E]�p��P4�3p��t"o��d
���~��Exk�K�n����O|�쁽�ݰ&�=��xg�P�R���yB�B��B��j�:����&�/%�� ��L/H1upӺ=PV�IF�%���tu�W�trɪu����X�i�,Tvc�x�N�����$��˨c�\\G(!_�^Y[���h�x��Y`����PYY�܅@}tR9P�P$6ǣ�GdF����o�s���"�ؘ_]}����z���H�-ޚ��$z��N��H��̈�X��L�獻wRݐ#��n���p;t�_!�@;1�d�2�k:��@.��YД&fVx!���'�L��M�A�&�2��'F�վ>nTB%�?SƫQ[Ql[����m)�p�y�k������$'�|z�w
F�p��,�x����q�LdJ2O :���V�x�I�c8v��L� ���FGjܾ�1�;AOQ�w�s���-��<X�O��st����v��1������e��#��$�8�wn�w5O�Y��n�qr�m*8	�H�N+l{FhI�+l�;&��Nhi!���3����=d�5Y��A�ǰ�z���Yo�h�8�aII��7uu��w)=���)n����y}$X�-"!�K`�3�vww�n��`�}z��W��𰄃C儥f�u�f�q(O�����ȡ���%�����>	��/��u��:��"�D�{�8Ss�E3�8**jJ>&d�XQF����AA�G{a����K����SߌB�B9�ʶ߉h�ec�E"��!��p��7�!����J)�(,�C&�ݙ���sxK���}Ci���𿢠**�4�x]��IM>�[��w|5���]ѱ	�m�##����rϚ�b�d��}
�&�h��p��Th���A簏�2j�}����#0Ӣ�_*P��UI��=�ț�4�_�dQ#����$3����}�!,8I���?��hK��^�X	�ǹɃrL�n�Px9}�'XQ�*x�٥\D� `q�� ��2a�i!9o}�W�4���R��{�1m`No�mv��.�Z9��A9���_P.Z�ל�c��F	�<R�Z�`$��1���U���`եcn>�yl��!		�{J��d$�	 �M�Z	����-w�~�;//�+���U�����TWwu�p���cuec�Z�G#߀�?����@�0o����ޮָ�(���{v���N�ċ1�! ���}^ij�5�vLH�'=�_�K��i��U!�滝��		�2Uf�B3�x �
�h�fy��`-�>�	0����"6�fw��ۅJ/h��^:�i���G/Ι���_���z+�o�	�������}���1�
�|f��A��!7�,���W����J�켎a�$Z����% ?<��ލ��
���ı/}k"q4!�!���&g�NiE@��cTp�{��}�w���U#w�"Ê��_�\}�4�|�*}v��/��7�fAJ���������\��xuo��M;P��%lO�p��N���W��]�Û��$"^��WWNUF�Dr�>���&	���7t@)e���{tn��)�D��2G��y���R�=N��	K�� ����	٥uq]��������f�����9����T�����q�c���h�� ��}��@EU����HV��B?�v�v6�7
@Å��Ă�E#R0�[+�����u!���J��cQFm	jK]�m�s[��d��Պ.ڥ��G�H!�:�"Q�}��ޱ_6X���I�(�S�ߌ-�x�;�'b��;�h��8��݄| �L[G����}]��5��ҟI�j;��{3���=´\�]r�S�����Vu�Ϧ�2��}j�<�� ��{�7�������l��0Nn<��nWBL�Xj M��c�?�b��̴��Ey�)���hM�j��)��>=�����#�IÈ)��R�@c0�{����q�qȪ7�@| �\��
��9�![���͇N-w$�Yøiw4��E.�F�z�>��Q
�匐�[���6M�LC7�$ֵ��Ǽ��Y���t���>nNa�*�j�j�>ŲC
��Y#j����ww!����q]�=���>�����X-�o#7�}����^0�4D��\#�\]�����  �QZ/cg���ܧ)���MUO:{?�t���K�����`7 /+��F�G=��<$��#y/�4��i��=-�7��.cx���aN]���6g����r��������!���2s��WX{X�O^�_i1([7v��+Q�4�64�O��e�&����t��N��f����\]�;P��ɹ�{�+��,ֶD/W(î4���������}������O�o��H2�A������W��I���՞���,R߀u_1']�l/C��?������zt'ʶ����'?e=����l	!�u���I��x�bxB�b��Oe%ϖ�I2	�u�G߸V���o-��6�8o��?a�,��i��VA�>���7B%z�M7}�i�]wT�X�M��3��������ӮE��²��y�����R�l���_҇zU'Z��&k�o�E�Oc���(-S�QPP W��B����5'|�~���;#o�T����?��v
�����qf��ʹf�$���Dߣ�{�*#!�D����Y��o������fI��b��!�O�,���J��L�#/������U�����$Lz�_������˃'��MË4���;�ԇ�s�Ԑ��JW�8��>v�U�a�Y䅕,%"g;z\:�2Ps��=��9}s?fy�[�`v�H���LQ=6/nnL�I0~58>.���<Q�@�A��nݓ�+!�'�����H� c����"� ��a��/''7�/2�c&c��?B�zS��x�&7c��k�7��=�fs\U�۠�υ��h������Zm&�R���a����iɊ�[�o�M��b�����7}�-0bP?gY �d���h�z��Y��L!��"�e#����:�����~�xZG:�E]�=�z�6�,��e �/0!T:��ΚL!	�����$k9�t`7Da ������a'�y̸.]@ً�s/�
�|�5����q�4�y�&��Z�pw���*H�p!%M�����H��C�,PK�[�ƀ;�������F���?�Ĕ��ŵ�Y*�k��lHU��up`�v��o~�7�A�4��o�H-�$Mg6ҡ�cG|�<�(d3�}�\��0�����4
N�\�IZ(#����n��.�d���ǯx��"HU�ڟ����ڣ�%��8;d >lc5T�Xl�@J���G����ڨ9��e<~�`�:��"feE�K�J)�(��/��F��9}�[�J���*�"2���>�IPTU4��F��ߝ;M��'����[��,�t�y��q�x�/��\\%ݹ��ף�@�Eĝ��0X|�!\��:wrY=��<��Kж�`�O㙪cW~�����(F:h���О�+����fs�1YK���@�WE�U������m���KO�c�]��X ɜ�zD�y�r����F�\��$�u7"//���Vs������Y��ь�M��*��sc���]�k�4a���h0~��n,�[��<�:=��@<.?rFr6z[>�n����������m<Id� �T��<_S�A����~�ɅF$��-�j졒Ä�&8�>�o��������v�}�7�~"�s��i������e�kN�\�tO�j񩂘��M��+bj����}�Xҙ�F���#/��CI����v��7��Rx�8~+Xo���zz��zG�.yV���C��J��Aj�i�QEh��p�0������=i|/���J�S��艚�G�>�۶D�;/Rh�"�0��/��6.'�je�%)Ѝ��]�"��յŦ����?A(�����hm��>?2c�F�ZxH���H����.|A-�)�� P�b���=?���"m�H�  C�"�?�hD��g�V����^)3�?��3\ɠ�<S���㗥��_Q*���.�o���B�����[��;�muAV��\�/��G9A�%蜰��TT�w������؜�Wٜ�(蟉��^}7N�"�O�Z$�7G��XN�;DGt��}_����1+x�3G$���r��h��c�U�%o���X:�$�h�ء;3.�P��qq�L�(�Τf\,���JM>Y�TY��rW)�E���r�~��A�]�Y
��M�����(U����h�.�u/�Asƌ�QD�j��9����&�:�M8�����}�^5@�\�m���%(0 ��	qq/�����S��M��	m<]>ͫ6G�"�@�s�X�T��0�+^d4MDD|1Q[4��c����.}����C�{[����Q0�hQ�o��p�7�FU�.*��5�xkm��S}hQHPMe����6�+�;C��YGʎ)��،�(l�kd
6�5 q6XlASgf.V���A�Z/� �����I���$ޥ��ƍ�$%��v�u�4�y���ōԹճ��
�*�x������w�J�;`��v@V����hG��Y/��Etŭ�R���0��'(�'��b.ϣ^EW�5����p���
6�����ېo���紙��y��)��+�G�
�d�ߣ�fff:��u ������� �y��Gy��iXLg�؏=���E��=i�Hp�N�� �v������%��������f|җ}�wG Ř+.s�#�J�.�AQġ�f8i� omYkG�[���kk復��o+�GdK4�K_M��'�J�:�.:Ma�V���~��=}i� �l}B
3ܵ�׵�B#�PGt?�k7Ӕ�!�ܹt�IY8���R��{�_��YQz�
�R�M��c�V�|���S�ϓ��K��Z =P]�����˓����d2��|��ٯ���k>�$�0���@4@Sew�Mh�7�S���z 
o���2�{����wV�L' �����}��ɭ�g����u��@đ�uZ���z�qB!e�jSY&�IMK��HX^� ���.�#|��e3�A�R>\�4Uk t:��ߎV��+���̅�;��*�����X���rF��&d?G,rˍ��XĂ�J���,2gG��d(�s֮��R��W?��@�AF,�����x�ú�_���`�TY{�d@���Bs�25@��v!yCxy�$�V1}Xi�_�_�����Mi3'v����Ow��Nw���婢�� �E`�k2v�x��g��U�ai��3# xx��:�M��a�t���4LLTi��`�j�QYP�|ca�j�V����2cR���	�B⓺HR1��}�'w��PV����t��	��u��QV&<�(t�mĖg 6w"�jSt��-|��3!ܞ*TE�ITv�@�Ż�#
|3[�u���͉BQwuMMI�j���������,.1�X��8L������^v�&`���0c�Μ.�#u8�N^�Yz��6���y����x9bk'�4G~���u�w�X�%2쑿�>��V-/��$Y���gI.�����Ӷ�yL�+�`kk���Am��)o��c�&����1��YYL�Kɩ'(��Zt����y�n�b��߼=d5c���J��x�U�q�4@�H}���p� y��z���1��-]���d?Z[�l%I?���7�C���v����G�xƀ�܋�'�"�L��N���-ճ2i7;U� ��8I8��|�l�]�ꆝ�	���:�E;����*x������*ǻP�;g�@�.���R�m��w��m�v�'��#����l�y�2؆߷�.o�:��|g�f8�:G�||^�W.�����%����?��BjS,%�+��|eq0C�H�N��6�.S��M����r	���j���d��QECr�'J�fy�+D�r�+<Ê: �g����-���>p����s�~�Ji�|�ϝ&Yh���Q/2��5b��k�Tf�Zx]�S���&l���Y�����q|m.>^�����g�čMڜ����?'-^��@��l�]�6n�,����a�?m��%|hi�2�����X��½/����48D{�J	/���iI'ww�=С��}�x~~q�ĝ~���]},�O����G1���oC��^\�J���׷�����& �S��G2y.��r�k��o�����I았�~�h�w��+.�*�[�,h[�H��i*U��``��]�?�&H ����i�݃N
��r�m-f��������5DX�J��o�l2�^��^�5�Z�y��+Rt�m�[33�2�`ly�z������cy�$]M&>�F�W4X8�h2��C|�򅍕٩iŨ����g����^Mќ|���/�4�4�������M��¿�G��ص���F��@����oX���^�<܁�7��BH~�ϷW��'\oz�!��?⛊U�3yW�� ��W���E��p�
Qk��C<´l���9��\�E��g�pϤ��0�\�C�Pݠ>w���WU-r.p�neyy�,��~�	�ଅFF�6�7�m�`�o�8Lr
z�C���o�P(q3}��~�ɵ��<vy��.�b�oe�#�&{�7�b�����M��Z[}7vO)]���/�>-�eLz�5�qG���N���G���}���ŲH�.��;{��%Ь�O��*��R��%���1�	3(>�#qm�H-ߠ�ҹ�ry��[t�L�'�|ƯcqhZ.,��Xָ����'�������l�ڮr:ԧg�`�_Q�P��G(�L+3w�RV=��o�9�J���֒����<�`�c�`�G~*�������z�J���	��F�t ?��R�~����:���@)�`i�������ۮ���*�Y�u�,���_<<<�2�V��?\^�<���K�#�#�O�y�A������,��T�	��>U]Nc*Y3�8�s�08��\i$C��#�P0�K�2{���t��N���&�#994�!+L��ѵ�:���}�n�a�i�J>����}�:�V�۳q�I�¯~����$gB��~�'��%q�K�+��vkw�ҋ��� Da�����_A��H��W Q�����~d�>Mb�%�ݝ��t�H�b�гl]#>ص��i:���a�it��GC�i{z�?�-���MP�-�t��_���
�D�:9�C�r���,�#��C�ne7iȏ<�^�&`WMvƁ�e���i�����K��ٵ�<G��nK�Q��g.�I��p�cz����ǚ���S��S�`ȳ��7v�NDp>%I:7�,J��}[`��z�
���ڷiJ�A���E��o*�ʜ�`"�wȒq��-��"���l,�����˴��D���|��]��iH�KJ�8�I߯`iN��P�&��r�~�W�k���2>�.�ܪ�i@�aT�ɞ)Tn�vd�W�j	?�i�I���t|�]����d�A�b��O]0���y�}吲��/ʛ׎#�iL�V�4[P������Z�{��@�	��`���7�t
�v�s��}SW3B��p2��Sz�;A[���'��T���W��=fЩc���S[�U�E���F����x�1�J1�k\r/וOഹ3���F�^��ɿs�;\:��	�b� tt�@i�H<T��"i]цF�f!� ���%ݘڌ��Ln���{@�v ~R��qyg��YP����Vn8	?rˏ��8PĚ��V?q���< (�Xc2 ���RH�?R�P"D��D���͹˨̠.3je���b�qy�MKKK�H�JSEܶ�Q�p,e��"<ω%�E�VN;�zSy�Hanp,L�C��	b�X�𩓻�u�r��@4 �sU��s7�sa�����A����}X��i�.Pmt[W]0�uMN2G/W � ����:lY�uywSzs�Dh�>?�p�� f�������6'�OD	�vx�k�ڙ�q,�{7`����!P5� y۪����]�M0S�����Ki���W���K	44���G�P����jTo�e��U�>F� Mf�����9���X�1ø߄��ZG��v�mܟI������6�NP������&���D�)1q�����>K���ۛ��\�?�����Ql?�"���:O�O��ӟ�����z}}}�aϷ�����L�oKY*���6<�>>Җȅ��R�25!+����+����i0���MCL!��{�9�GB1KE�ROa���lz7�'ů�~5���Hw�+C/�G5I:C��<�g�qq���<�@za>���E�:QG32W��vrvN��dt�wS�O������*Ǹ���\K�Q����7'd�P0��� �9����F�ń�������>p�D�׸v��|z���)��FT	�D�s��D=�v!�����P�"�umg�z��1P��1���>^&rWQ�"AU{%�s��d)p��r�}�ad�/d���3���sr�����L�tM�� �~:y���o���#E3	nKh^�'�c�LM��[P�=�����	�}�̈���z�i�-��Qr_�LE7(�>OQm����|������F:v�S�{J:�������Z�X��Lͱ.2^KCGVą��)�lVh�V֎�����z����k��	���	��!��<@pwww��݃�;|C����_E5U3sz���ڽ�ilj�P+l��+{H����f���~)���خs����a�W=�Ԥr%��Ĵ�jňB�sg����W�Z������Y\zm�����~�Z��{�h��.�~��n��U���(�1�K�Ҽ;u�- �o��l~������j�mi/�uJ۵O�v�R�U@i�v�)2x|m���<n��"����ݣ8F���U��tE��t��C����P���=� ySܝ��?�$&�Ua���6�"(k��QI�B�4��ŭcg�C�ϡ��v������G��WYZZ�}vϙf�/����c�M�MGK��a���V����3�\���������Îo���  W��{2�'���$���+���[?�y;,�=�7�	��#G��S;����К�߱��@ݜ.�7�l	2�����c��0b�I!o�S�GYC���ۆfIЃ9^��
D'�����ZY�'<�`�N]_�|�DO�e����!q]Ά�;�+���1�����څI���{h�;��;ԓ���\{�//2օ��l��z��IX�����؉ѫ��2= L	'��w��|��`&;��$1�q��^�lJs<�|�qt�"�.b�����t>�}�ւ�������[[2�I��L��2 @��q������
�8��=
�]=h<�I�w��V���;�pr2��`}a���\.v�\D�����Z����<���Ne�ѯ��:pI�/���6�]�CX'�B�2^��������c8�v�	��\�z}�U��b�v�}�?���V��qo��b�(8�}��B�Z^N���'^�h2���齆�Ζ�X�9�:Ib"���^�t��򃘇0�A��G��b�93����U���Ȟ�󉗍 Y=珙f~zЃ�:���T�fQ���q���as������l�K��n~g`g��~4�mm�*X�J�˙�U�Շ�����~�_��Ha�&W�]z�f�O�9Pt?���];Rd��%8_b���>=>ޖ�`�/#�d��Ru��v?|�7
�N:�lp�ϙ��v���1U=�]d.d��bߙ'l�dlXtu�X�w��m��ϵ@�vȪ%'5����W�{�����
�����zit_ �cߴ�m�9G��5��^����"o���~g��7p����$_��S^�.�� L[ʍ��ax�hȯ
�@�*Q�I7!v���f#W3W��䎰Z����$&�g���N�N�.�M���LF�Bч�h�|I���OL�eڞ���T,,h���Q11)�i��~z�!�-\:��R}.����JS�o|^�	���֏zS������&ѿ����,��/94P�u�I_�O\��`���4YA;���#�FU��0�z>�0$�C~6�S�sGRCP���p���y�}rH*aOk�ls���'�z��V�(+���U���h�����71Up0��D`{#�U����P>=e��/��GAd4e͖N>6f�|��=�Ŝ>�G9>� ]��f��Dv�K�ku3aYz������e��g�]; EƋW����Jd<�)�Ҿ�z�6��1����@�c�4�u"��������ăC 9��GO򇧶�nr�v98%��3;���̯��*i�Ye�����r8Jӳ{ϓ~Oc2�?��F(���y<� <�3��ЙV0c�v��j �~�@�boΞ�Q�i�ޱ�|cp��nx`C6�(��:�o z��Aۿ�s�w�u�V X�{���m|X�F-��u���+П@�n3b�
8Ī�d��jM�5�����/j��.>���`\��&.}�����_[?�+C�x뢭���_��dW3�ٙ'S~�dԗ�b�ɼ5�*k{g�FQ8������o���K���������A=�������@�/�)��������9
8��Ad��F�����-'��;�-�?�������ߙ�<Uc�fָwp͗����ΐ��]2]u�v���up㇜`v�CU.#���u��{����ߘ3ӮWq�4�4��'��
&�����*���G2#.^J�I�J|��Y�I�+�Y`zf+��|���Ǩ���=^,̚v�GrW�����Sr�AR#�J�'�V�J�c$	�S]e�j��f-��3��T�ޜs�o6�&U�H�w1,`_9�2������ڞ$K]�:#��u��1�3/�$Aϫk�����$(

�w2'A�����������a�C$"�0t��yx3�g�,֞�:^�0q�����l��T١M��`�2��u[v�Q�  w�G9�s���
�ݫ�8���Mz����|�i퍤��x�Bqay�1�6�Æ/����y��Eq��|lTt�B��!Sf�n��6��7|Vi��qS��@-
2�bH��$��u�����n�h��>|ė�TV7�������b��`�v#�J؍�*5jV��߁�X�fe}���X�0**8����'-��hMmZ�ݙ����xh�?�R������+�9ɸfqz�ҧ��Jʡr�Ը��2���j��������g@Iu?��MHT�YOm=?J�eQC�Y},�7��u�I�#	�U���	���ĞN��郠��xJ����4t��*�^2�*r���}�{_���եs��%��I�'��(�����(j"�������@�n��@U�V��9Lz�zyQo-�x[;<զF��:�9�l��76:fl6�]���ӡ^XF����G���P��x��0�:����1�[���Y�)?:)�J5h�޷�MH8�s������I�5o����spl���H�6�7�iq�&(�*��9#����XKq���q^�gp�J/��u>9�}��x)8�NkEY��JGp��ۻ��0s7h4e:����tb�L�:��rEz�Hjd�k(m{D��<�ô��#��z},���26�����#���ˀ��s�����6�����I�v��	�!��K��G��V�t�o|�\֭/��*�ăQF&שۼD�{�;^ek�O�<X�Ү{����8����4�!�����zqH;�<�+��^Fd��	fL3H�= �q<�a�╦Y�����J
zj3��4O�si���㳍W2b�y`�-�d���:̶��X���}��S��O�Q~�K�5�(����	@�Q�q���4����"��A�v ����j��x���ec�W:A���G8v!?Eab�ص����@��šc>ޡ�ה���8��N�W���t!��D �{�M����$ւrV`��#�A�E��K��W��C���`ڕ=x�|�EI�T4��!��O: ����Z���K��eSx�4-O��$N�6LK1x�iԪo�W빽��݁�W�
���=��f�lRw^��}�D�y��u*w���Ι~�.'�2��N�ḷٖQ}z��<��Z���Z���7U'���3x^����Φ̝^�T��#O}�Aɏ��	�on�9YA��Z(��E:�ߙ����L��\�&F�0&���a&���r�A�yÊ�{{�'�5`�X;LԖF.lN`��9$❦f�ɺ�A�m�S�m�7��N��^~=ϔ�N�a9.��0g��i�z����D�l)��ۄ?%��+��j�����t�>a�Z/7�Ě���=���u�}�����W�I���1���;=C�O;a������c#<�����m�C��g2�qL������<=�	G������/�����o�eh��&i_g<+n_N^!�j��Z�$0�|��/���KR�ɹ��������b_�S���4!���s�c
v\w0?f~[�ҳ��PV23k���7F�[7��U=�ot�Ͻ���z����n�d���v�_t�ۦ2"bq7�\7oe�b�{�xk2�����V�cg;��#�[_C^UO�U*ԓ�j��e����a�賟�j�1G5��5�f��g�����oAA�L�*����=�'VsN���z7����_ݽ��սY;�e���M�{ ,�.��Z�^��~��3LaF�=�!,)���$h�T.�+��3�o�u��3��(�ԫ��9�ހOO�l��/���c3b�F��.�ݵN]D�V�t�jɾB�v�l�Pz9�i F݂b4E�;�3&��u�f����)qE~�XU2P,���
K"5�c�}�#� �6H��ݳtp�`E�x)5"��l���r0r�ڪ�$A����2��I^��Q�CpT&�:_Rv�Uv?o��O����(c�0s��p�J0"L����F3�*���e��r���LɆj�.��V��OhhZ@�H�E�î�>e6vL�4އ��J���Q"��wrr8sؓQ/Z@�G[��>͉�H<{�ФP�3� �&rc�8s\�2�������4_�����Mo���"�C�T�[iNMy�u�yB��]�u��MP[��.��(�	-ma��?8rx#d}�OE��|yޝ��T��Bm���ɋx��B�?�{�����������C�1^�^��s��n���߸}�<m���S�`���a\'�C<>�V|2[f��*9�l���D�=ͷz�(�͉�,���Oi��y���V�g֤d��{������"�7t�W2����C�qz��ή��W��%�U�E޷D���XX&o�/�!
�~��۰Rr�۲�����<�j�_"�����+D響�Wr�!�g�Z����Yպd1��W'c(ZP�N:��R�9�>4���5g�--�ƥX�4u4��h��P���V�#j��Z&��q�� /w��}vw ?�=��y ?_��s�h�r��M�s�9�FҩK蟟��nv���9��9�`H��1�܅J[�P*�2�n�4RG����p��3cv=H��7kǧ�x�^��IA��|�0)���,nN��V�E+����Ց�(��g�'A�J��M����A��u�}�>p鞾�ʥgg��P��z�
�������o�+9����t�����2$�<n�剻�lhpEH���������0��z%܇*�uTZ�Xb��HP�39ߎ���h�{y�(��ܽ�}��PUY�<׳��<����e�� ���S�:3K�ȵz~\iݍ�����L�_��b'`��b�*z��ozͥ�6�`�%B)�0gŢ~g���U�xڡ)5��J���m� �AG����pL�1��
�ݯ��S�;��Ԕ�CV=V2�ζW�3�f4������cz=�}H[~�Z��w�tfK��Q]��_ע27�������e.)��?�J�b�NS@��̔��x�뵚�:�j=`_� ��Ur⨗�]��õZ4
%�?K���`Q���Q���'_KəK��u�#(Y����?W4��OEDh��Oj���C��7|)4�"$j�����T'J�\h��<�Y��)�=�Q:��W�q|	�����N�1Z�e0��"p%=�Bt� ��?�5��)��?�?����[[`5�߱�CE��@&��bg��V�s˦���q�h�o���Gm�mc >�;�s��E��@_����ᩓ5=u����:�ϰ��ӈ^s�mm=�2�U�(�s�zG��u��p�f��#���M��U�b�}ϗ�ڧH@G��Pңe�L�I's��J�����[sl�H�9�-�r��uU'�V8
�R�
���ْ�0��6���`�R�u��T"�^P��7�y;�힤~6��u����\�%V��%�mK0ES�\N	���PI{ؿ8Y�6X��F�&ɨY�� ����y�~���T\�S�U��F��ķ*o�����!�e�1�b�7�e�^V"����zA��g�q~6̘n���H�KcA��JI7"���M�����k�g���,��A�<����ݘ�Y��Ҡ��O�)hO1����Z�So�Z���C��Eh55��Ġ�������@��%�$�[^�o�������S��B��lƧ��{.�ܳ�}l�1��}��
w0���c����-�~&�XPt�=WP������L�����lq4W�o�URV�Yn����/L���|�m���V:ܰ#�.(�O�*�d�;V�'�@�C��e�8�\򻎑�+z�ZKGTɑ����k{B34�﹎JL���}���_-�� &?	B0wV�g\�m�m�"���ڭH�Ci2�J��.�$Q�uAś7t=���^�N/�o���z�mu�U���M�݉�{�p���F�6�������Z��2*�MT�e��r�J�
*�W#�(n��R�^��g�'��������Ο�����! �[tĎՕN��v>t1�+T"��?�~�IJI�>�j��::���Q�|�I����+��@��dmV�n���E&���q���!���OWDJ�W!6����."�?�n��7���Z��@��00����ϒ%Tst���-�
��j�g��&tc��`>u�#oTЂC���M]��~'��2�9V���&��d�T([����a��`����@�����o�.�ے�"oZ�eŭ�K�ʷtst��4���l.^x�T��l�� �F1^����Fe�w^��?�J|�Gn���k��f�NL��0�1p�Q����a=��'<�,Qs1�\@�6�p��&�D�_�"�0���_�Â�G��Y�
���ثkdw�'�c<Q�c�Nsi�)�/�k�{�J��(A7~�~��-˯�mNgv��
�G��z�����h��t��n5Ӂ�O���D���q�$R}�ۦ����k����t)����W��O<!����v�Yn�ѹ��zV�
��4g�r����X�ҵU��q�5��J\$��rs3�Q��^��K4���aGu_%�eS���Q۞̄����|^<��d'IACו��66&�{K�P�b1�e��6�J_��4�p�/�JL�����1JH)� )��:�B �HKU��w���cA7���zE�i���m^��/2�@?�sg��@YQfw�q�<��F ^��̆[O *��*o�Hw�2U/>4 �o��L1������������DӇL��x�w�fV��R��8�Xw���;�Xp6}�8w�}��D�oTr�
ڢ����v��U(40_��Jɼ�q�S)��P�\Ͼ��Hv�i����ÂO��E��g�.�C��f�0�ɪ�w�V˦C2�I'yXR�T3x�O=�����������3�'��%n�pj�d�h��yz�R$�7��� �Wd�roj^�'�;�Z&����e�����q�|=�pպ�	L.jX��r'K�l���r�,��u�����0�T��y�$�2~U��+�m9���ܪ7�OOa��}�7����"Q�4��`��;>�:�"��QK��:5.��/W�_�5������������$9E8���D��1�VG=|Җu�vӉ<[Ƈ8�rk����4��E�>�&!�M�iD	�C�athB���דC��b�t_f�m� X��#�)��rXl.$�6���}�osh����-���%��{B�+����5G|z��yv������qN �)P���r�=�r##Y"�\��)�j�{�Y��x&¹ݛe*�O͎~��wx#HV6ɳ�kv'K��Ѽ�@b�-@�	 ͽg���^��2�S �V-�ӳ��Zd�ن���X�>Q4,f�)"�)�ז�]��� z7��V3Fm���D�-�b�Ag{F��L�X,�ݛ�sӯ9� �H�<6T�`�n6&�X����Tw�K=��Sl�&� �E9�hc#���r{�_��INkiH_��\�ލ�c�d VY-�����܂ɞOC�TH8u-�S�[�j2tp�|{?p�ą	����t�u�6�G�,�� L��[��h��w#M(H#�𣌕��1��nȆMV����|�6�C�Ł?�H�%X��̟P�F�3~okx����\3:'ec�(%%%)++
��Z��W��¶�xdT�R�����R;c�K'.=�Rz�6L�o�M�A���W�ñ�<��A[�=n�;��Аz����=>n������D��a�T�+���(�xhQ:<�O���=W0����������Շ+��`b�.��گ��2����_b�_�}�:�.1�t�@b9-w�ά8TY-�0�}�*��}�Q�w.������$!�� ��	L�]���-wqFD�DyR%`V�z�un�~�TUMZJ�oW�f�6*l"�&��H��G�&��m��>�G��2"��ډ`%q(ͭ�q�g<�X�6�M_J��ճ���1�{2@�kW�Rw��$�஗���=�W��{�a��2-KΟm�(v�5}�ع���r:�^{�?��f�ś�Wsz���ߜ�x���Q\���	��j>�f�coB�e��ˮ���[p��u�|�b��?#�Z�w��b ��`u�H~�̝���{�e�/�M�W�֧���H���z^T��3H�L�=�_��v&{�*S�u�3�'ϊ__��O9y��h]��{�l|cw�+�P"�L����N���.�����hs���X՘knX���	3z�I�O}���L!�u�7��Z��k�㥆�$�U-5�8�g��%�JS�"�f��;\���N"~�p� 蟒�����s���̕]��Wy�2����]�<T8MR�Qz��z�L�6ͳ+��&U��>���)��l2��n��T�;NL�0�:e�{:�kY38�:!��?y����C� ���<������Ъ�WFh]�SKw"Ub�c��mn?�;$������l��?ͻ�*ˌ���<NR�{�c��I&�u;Ȍ�	~^�[_�1��98#���v�_»�!WX��H� $L��w��Ŀb;W�ՙ�\j�[G�F�Fnu���_[=��N�5�������v�r����^�و/�Kۮ)`@���rr��K;�i�J|dq'�vXʴ���\�{�l����D��K��>M'#X�PrK��g;^�H���mYnm��$����Ӻ��%��|�q���>x�����A�Y�� %��ayk/ݴ6zKk���LY��Џ���/���SA�Ռ��{��o!�S���S�k��|�S6o�zi �eyv�l�ge��$��u�[��ŷ�n��
�#�~�o�栫Ӧ�����CJ�T=\�$��:&�qm�a�F� hf/� UV��#P�)Ÿw��.�p�r�`s¯�����$�V��GCe� rOGS}�̭��#u��W^-T~�^�ϙ�"�Y�ζ@���j�3ÿ1�[����)m��/B���U"O$��q���j���&Z�����K ��5 b��h��J�p��W�ZE�/#���\8'�U�]T޵B1��"��=T�"��U�@)�jyl���<�uT$��?c�,9�;�Zq,�L_�la.ݤ��I]�\�J٥m��piS����,�-�j�gXY��~���Ã+��
�J��i�mj«��@a+-���$�o"J%�j�;�96F,��$���� �IȻ��Ύ��	BaH��v�$�THŻڐ)`�'�%���ۓP �`4�4��X�\�D����֣ܦ}�{��uD	�V	��.b$��!�/nXrX�-R�]���G+�wC�R���ꔵ�Ea4Wn���P��+YҶ'��T>Tj$�eFIA�Og����LhVK����J��G��d�8��A���u=�#��\<Ϳ�j#5��Иc	��|Bj��M{Ý�?��&k>�^���faa2�J�^���z�Եo�M�f���LlųC
�~���/�l%Be�ĥ���A<X�L�=��ʐ�܌�1��TkM��C��nF1>H����T��ƕ���k+��:�Y�=�N��؈`�n�����!�����v����0��D0��� c5#=����tAj㺁����1�|S���TQ�Ș�|���+Į���gf<	�F��B(�$�
��uE36�׵mF���T�fd��܀ͱ���`�I\�$[?��c�~�I��$�m@�k)1/o�_�OJ-�,jTu��ֽ��&�M�����h>��(FW����8����ʃ8n�7�K���i'����)��n��do���ٻԅ�FS��ٙU���`q���JTF&���V���\�!���N��VH��EE��j��m�Ʃ70?�?I� ����7YD=Pq��=>���P5%����h&y����?M�h�n�ï���6���s4	+�����4�����R�7W��(��B=���*��l#|���5&�F?y��#eS::�{W��qj�3!���o�d�=�U��"_���
q�k�7����4�O�����a�і���n�t-��-�6M�+,���"�,^�"ӍGt��k.��������""D��?���j��?cf�(��t�$͢{�F���C�<YyS�!'�͖��3>����⻤^e��$-`����f#}
 �s��P`ܮw�C���f"Z?�x���t��ڤ�s����:/U��/Z���,�2�@kU�vmc�ƭPñ�76�J��7�1��SH�K#)�x��U�x��	�� �yS���,ȁTϕQ�����m��lO��$�K�c��BR:���ٺ�Ջ=�X�����G�3���	���H\�&��4#"�`�,�M�
֝�Ns޾�8/��!.��������Ew�����y ��<@�>��b���#��������8�VW�νѪ�;q�W����Ð�W����=��^��0w��߲�4��λ��%,�����}Eĕ�Ȇ�	%�p����)?��M�F�:�CD����� Ֆg7vA���P���z|m��'���ϵ)R:��SD�{�b?��a�gR��'���>��wZF���%�a{1�؜�����NވoO���I��9�]��]�T��<}�y(��g0
g�^-v�$�b��C����tD$3�����ǈ�H6��Kh��amJ��3-�z5��GqQ�LS�4��/�*]��k��\�>W���Ő��10��̪����G=����*5x��i�O./�S�u��ܑ�kQ9U���7v6B
�v�xTf5�|�{ ���!��C���
d�$��fPC��r��=�VAI���Ǐ���?�E>�J�]���+q΁�7���۞b�#V�AW[dn�'~�z���/����|�]�3����k�s�9���Wx�|�v�uz{r �����>Sc�1qÅ������ή]a_�yxu��H]�H�9SS��w�/�h�.�_!��@NS�:)���;/��=�/Q�aA֐�m��
�7Ʈ�V{�&��潶EpQ��%�<ÈRdB9�<��b#V�Fol�	�;��(�C����n��� �8�?����x���e�ROFO�g�H�������"q	Vi�HzFFd��L�>�b(
�{�@Y�c!6�ĶƷ-l��q)�ҁ|t�vLٳr2���@k�6⇳�*��	�����V�i�x=O70�p��|�N:z�a�{6�r1T붐aƙ<`�6�Y!���kKK�]��(�a�f��dm���x2W�=�±�i%��o
�'H�-�<���A�%�<%���sp?h�����`A>B��vDm����
,SwҒ�����m��bd�s��{�e�A�V���7ٽ�K������%{���0 3�c�O&
ԃ��w{�{�m�@8�;9P����J�ݒ��$b��f�Ǚ�r�@��_�b=(����� TȜ;$�5�tE�n���X�j�m��{��	��Yu@ߑ���Tm�F�"�)X��d��2�G�m�R�+��(G(+�%R��{vR��Sg��ѽ�T�8�C�f���nZ��jB�[�N*G�棠����8�%|O�܍֋�����m:O�_6�̇�]�r@W�ݣX��e�扲��d^���� zǑU��u��e�O'�gf�� �͏�;e�1�x��+��}��q��%�2*H�n2��J��t��y�����g�׷����<�@�D?V\�p׶�+��%6�L�4�#J�Y^,�v<�_RV��oL���8�]\\�G�e2R���HX��N��(4��^�CÒ�w��s�~�q3�ݨ�4��a�0D���zYI�7a����]n�����˰&-X�<�UpV|lz����*��G׵zh
�=(4���� �,I�g\&���RqA����n��=d���&������s������DO+�~��#��ض7�����3��z�y�Jc�~6�LYfbh�G:`]��G��)���3�-��?K�V~��/p�$���:J�<Z���,~����d��}תC�f�d�帤�H�!�Y n������2�n�$!����O�D��?����W�u�Bp%��fXd��F@>`�Z_7� E��LC7XANC9&��tm$�!�R�iz��[��a�i��j�:E����Mhʙ��s��-�qt���č^ ;l$w���E�w����Ë��߾z���fm�̻�{�e������ە0,�X2�f��cI��s��Z7��[WT0���_-&>��I|�ߡ���~9`�,��,R
F��g�Ko߃�%A���<�E��>�#=O���Uy��͵�Ll|h��oxnwͅJv��b���	���8_�[;p�4����.ɸ.�iA�Y��g�VW����._�2��,���`� չח'��o;�_��P�����b���HFʹ�nZn����R`1�>�G���}/���R:yh�TE\4����
{��%�?���q55T��-�!�>}�?�?`�%5w��*�7�K������(��	�w���i�^yV�����G����w��:>�!���������O�eU��ﷲ!L��Ϝ�罭����g���d�k�~��J�7���� a�rK\ώ�0�,߶Mz���/JVc/W��z���`����X�
ă��A�v�2��ǁÚn- �% �?�O�y��$�V^�B����XqqIhL6$�U�TC�y�<�v�����J�a�*(�+�fl��z��s9d���fg��|�ES�F�/ !U���+�J���[V�8����҅��6-���h|N�^�@pJ��Q�u�P����f@��(�罁@9�F^���k�:p/wæٵw/ ��j�4����^?���hأ�p><F�@v0�tZ4}Y�fM�ʮ�E5�?�q��7:$�p~S*j�����������ǙN�����XӳNeL߬p��2=�8Ӫꞗ:5���(��V�U Vnn�_�e6WeS_��i��rC��G������}\��Is��B<�t�Bw-���#O�	"c��ԑ��;��s%?
B��}_1�5[y��z��J�*r��A��9XB�gӦT����D��:�_v�p��f�a=��Y��`�8��Rc�˲z���̈́�d�5�Aq�n~������ldy�YDS�A�f(����M��DI���f?&N�3�W�;��o��f�����Pe��hU*xx���	gg�������ն����k ��YDn2Ti�б��ߟ!����W�E�.5tVrj%�	^J%��xa�p-{�Ҏ���U?E�4�����>�>�ke/��oՃ���4�m��Cak��e����,ؽ�?6�4��M<-������U�kkV�'BJ4�׬��'\7�'�]�q��O�x�|t�>�<�EO���(Ќ�x��VWy!H�b�9��%���#�iQѤ�fk���X"���?��v�?C���o���t
l�ZUe�˖��2������Gվ�s# f	
�`�]���`F�D����2u�������[���Q��Z��l��b�����G �o?�9������]�"��#I_r"@R2ž���Җ��aѫ�_��w��.�������1T����܍��=6�B�>����Pl��v^��u�k���U`�j��p#�G����0�.��{�]t����ݢ�R�q��)C��A3�x]��[���@0�v�[�mΖ��v�;�ЏZ�{����w?����
�w���x���XY#����N^��B�̸~8"߉���3}I��zo�`�����L�� ,r
�5��n�LLo�z��� ���_݋W�?>G,����yVGoƱ��4R0}�1%(P~uf&Q�����:�U^�7Un�������>�[6nc��T	��oL��H���;�tr�/������{�p�i�W������T���o��[��Dp�L,����l��n'��?DkKze��Go�0ﭭ �<Y��ؕ5�5oo�8�kϾ�-�+�\�)��d���	���́f�p��b�II[;\,��z4�N�_�gP��i]�y��Dg<�	���ho?�+��-��*�#�� �l`Q�6��O�]|�.��, ��p'�oŎ|���8�AOC:�4H�i]��@��BL�|/��yV�I Z�O[�pw�_���8M��'�G�h�0�,|��m]-��-��`�����u{1��I�Wa�`��W%{�ɥ<���r���+)GK/�zO���p��b�Z��:z={���'�Ն��p$<Jb�8�L>�j������[�
<T�٣�e_�e�g5�}�����I
�t)�l��neCj�+�Ii�����-G����K����j��UI-M ���=gƍ'�	t���ϲ[�6�+_�v��Z|�����h�k����M/�x��]�	ӨXg�/ۿs��`�İ=|Ue��N�~�i�w� 7!]]�۳��U];׌�X��r�����J��KRTT�����$�c��?\`�Y�J\[�E�`yioL���'cV��CM��;�6�M�4�!֬n�~k�XF�8C�[^B/��'����<�wF�.��t�冘��`����3>l���m#p<
��C�������NȠ��z��"C�~޳m~�7$��GM�sT��f��ħԻ�?������ǹ=�lM�~��ɯ����fP���>�������g�]T�&�%*E��∄�RX���:�@�M������X[0lR�Q%.->��$�+�����cǦ]�ǲs��h>sW�2y&5cC_�P,61QVML�n�]@T)�,���9�Z������ʎ۱��C3Ug����T�a��`D��4."���Ļ/{���#l��ޓ�px�#8�cC�L���A~@��3Q��(g9�::4��'�[���������&Mv�kW��m�=E���G�E�Ek�Qa�i���cG3� ��=՟���u���

**X���@�����5��WZ�A����\�>��\���#7Og�z��Ҟ����A��ͫ�Pw�!Ѓɚ��b! �S�O����c�0��68�y����3��ي��|��b��(�\(����B�+שP��G�x`٠l��������)������7�g}�1S��,���Up��/��i�V�<-�rW`��Õ5�~N�]��7��_!vLL������g���xV�G�hL%)���y�����+'�玻�@r)�"RP�`�ܻX4�j�S����y��%�:��{7w��Tl��c�Z9T��R����h�q2����6�:�j]����-ƶ�Ɠf.Y��r�Ny�O'Ĭ�=�D����*���S�UPݠ�t �8���E�JN�`�2= �S�IO􍒂�j����ܠ�g-���dX���tu�x]@[s�������>���\C���j)�o���H��A ��d0W~�����d$F�+���q��b2��?%^��90��R0	�s���ܷ2��>Vv�����k����M����89���b�"0��c�ҭ�h�k���Z�Pf�&��1�U1g��~��9,~� H�Q�X�&�l�ƭݗ��uL[~�s#���_8QG*��?�s)�ɜ�����lw�6M�V�9ˋ�lZ"N ��R3�m� 1�8/��'�_]'<��t�zϭ_|�)m����4vQ���l�w*���[zȩ�����l��o����O��7�N�*zo���J���]ݏ�������h� m���GD��wv?^�1���o]�osm�>y��M +�:5��}	�������n���?W Ҍ�9@�B��}�Y���E�eC�Z6��-��&�ӂz;���9�Rg`~eB5a5K	���ʝH�=��`�i�9��T�N[��9{�7�)���b��P���#6��?v�_(�e�n+(�V`m7`��]hm��vHݿ�O�fL���gf��� 2��X1_�����{�q���ֿщ��{�7n5\!0	{���".2l�R$/V���wDe|||��{`�e��z@\x����6kԔ���1��m{�m�d>�rr�bq��b���B��9Sz��(bk3A�NM�d-��U��n�	��;�����Qx ��F"J2���}uOY���$�kwE�볉_N[��G �a>�@��
�B���m��6n��i`�����t�t�o��="�᠘	�ֵh��
���p9RX�Fr�����MY�*O=0�L�wBT�v׍����QY�4cF��U��X�� 9xU}ǆ��(�����)�����ɷ�zv02�"̩���v��Ӂ�b����x�	P��[��k�w�ݰ�݅�D(�2���IeRJVLa�{�j5��Y}�}�2`�%� ����U�|r��f�K� ��g(���s���@=§�a�Mg��5~aɛ����e��f��4�F��愊+yBU������+U/��咵L&�9��v�A�ۚ-�cY�g� 2���E�@�=)�Ĩ7��j�466�?D?��'�elȄ���=�&pŒ/F]$"�X��+sa
&ކ@,%���<}sx��um�XW�nW�]mo���Zmc�����նV�z�=���W�&���ƹ�9���8�CU�ף]�~æLۋZ,Ǻ&��"y���.�jPT�5��
�ɂ�K{h��A>�ڴ^���V�=愂FZ������nloדs����h{/Z��9�.�D�M�E-���#�	Gr��4;5��Ӻ�>WXpI�J�ڧ7i�����]� ��V`�D��]^O�I�>YWy#X�.J$�K��j��H<S������r66����g@kK���!%?��4�
���z�K�d��&t�Ĉ9���Іꭟx@?�ى�wU8��;Ĕ�y�y8���������? ˞����幅QǍ�#������~��>�&U?>��uxܰxݟ�<=?�LK�z]t���(O����l�:yDɿY�jR�b�W����z���wxI�,��_��\�t~� �d�B$;�P�Kh��Y��L�׾5��.�K�g�.����v�n{X�/��z��K/K�Sg�^�.�i��|�j�W,��d��aK�\���t��}��<�}[<��'ߝ�jU��o.q�z�����6М�ڪ]�w�@��E�o��t��<���Z���dǗſ�9łꎥw�6�Չ�����}���w�j��ZF���8U���@�ђ۝�+��߱w�I�ga4<�e�c�J�Ik�T��U��a/��
�X��퓉1�J�;�Һ��̰��g��˩�x�)ӕ_���G%��_E�X�bvY|�o	}�!�g�R}�a�E�ě�,D�� �Oo�-��Xvv����=�e��Ѭ����L0X����V) ��a���(������0�ǹ��F���'��Z|��Z�S������:�����s.)i,��n�NB¢���0�����N*���Pd�6�&�^�oߧ�X��t��!�yU��v�n�Fnw� jf0�(���O������5?6�M
s@2���q=V�|~ݺ�,�H�*����gA���Y�p!B%	R�h����e�á����8���G��:��EE����P�'B�Xo��ǺU���%�S�[��GH�U��M������:Y�/�k�ځf8X��<��$�]8E�����!��_R�P+o�5�s�v-����;P)?�Nh������R�[�vc����2� ��j���x$D3�3��b+���.�?>w����;Κ!�绛�ز���O.�mC7y����D&���ޏ��1�֋(��n�����E7�4��l�]���ɩ���8+Mtm�B������=ѽ�>���/�*�<��)�EF����t�c�G�y1���&׫~�Ϋ˟8�M�o�:�H}� 	Ӎ��?��\'<@�Y�����XrR��n6��~J�[M�x���~��`�m���f�It-�]��I����X� �|r�qrfM������ʱr�7���u"���Q�h�L����&27L%��7�<�4��#�NRJ��VY�/Ԥ���O$yI�IF�|0P�	��H8�5@��p�h�� Eߡj�+��ыmh^�jȈ]�bl�=X�js�HE�����ԵX���F~sXh�T3�����	�ƃa���a[�o��D�E
�u �K矃x)�l>���B�֖�����vs�x�Ƀ�*B�^� :�5]����IH� ���q)ڸ8N=�9[ 1���w����J͸�����[Q]�+_�?�	����9�rrb�Nȏ�noo�|����<�S���9A��<��Z���/7�P��(��d�n�����)J��_;�������P��r�+a�y��ne�|��C�+g�d,�t
J��Wb%�?#%��T$)���ם0qf�Mt������Z���\w���ܭ��6Ր��\-ݭ��b�0�l�%�(��w%�;��?��]��H�� Q��+k�AV�r�ӡ��xM���R��~)�{	FCv��2�a{�W�3@��=_�FqC�a�_j�j��y�3q���Ԯ�%�$�����)��i?���n�_"F`��-c=P�J� �N��.�G��>���֚�����9Z`_t/��\�4ŕU���'�g Ua�eXƅ)�a�[�UTT�H��t�lʜ?c}��i�����)�(/��B"P��a`
FyP��7J���oy���/ ��a��u�;8�0_���V��ﺘ�9.�~7j�8�����6�%����bl�R��n>X�$c/p��Lb�](_�w�7�����yVh��Z�g������Fh�l��Mf� J?�����]v�F��K�p���AX/��GP�3��fN���,���7�1�� 	 r-z*@�!��� �rw�k�,�]E%���mۭ~�{���Ϛk{y�u��ʠ� �)��l8��A!G ���󝳇�f��R�c�^F~��I���)ұikX�u�c))�,���,~^�Ƃ#݄�C�+i$�ke�pX�����x�e��(A�`���]���1>���ܮ�("b�b�4�J
��F"X����)�$�����@������X!��Y�Y�[����$ZU=�����EC�����;����6n�����P�;^��6����Pܓ5\�Y�P�'n~b�Y�D�K$�@�����f�S�C��'���m�6���-�H�2z!䱓��;�7]	�����|^T�-f1'�k�B��[���b�j��>ݯ�Sݻ�tK :��� |/�N��H�����'�(ܘ�2�#��V{�v��0��MYϲ�ŢZ�PZ�l����bX�  ��*�MM�8��>m}S8N�g�����ln|� ��g0�4a?��B\s������ؒ��`�������q������e��#Р]�4 �!�G�8�7!���@�x�}�Sҝ2N�8�s��c��6!w_~���X �Ͱ��l/f����Z~A/�<:!�OW.�BO>�(��h��u::����۝&�o�;v����J�oX���]�AVnG��?;X匒�e�`���\ݥ�w�mn�U����+�����$��UD��&���f&]�9F�s�k���I�#�)�����o��H d�&�A�,�Uή}9eÙ�vmS�KI@�rB��R�]�q�7���J��Ks�`�蹂�˽Y�.�V��u/FS���dP���CV�n\�7 ���gK�������������z�,�]�t�I��|�e�5�B^5�M�IX�{ѭ�7�`�|g0�q?�PET�@��~6iI`u���E�I���T.hy$�­��!!3M�c���m�c��-�u� ,���x3βZRt��h�V�)����霹�s��C�&s�����s������P[��>�xޕ��&R+I��%��I�K���J�L���lWo��'Ҟ2{n�d�D��~37�^�}���U��M�X�I*�,?ւ�;�f?����L��Z��tϹE�����6..G�������i78�!�B�L�x���0�=x����HHJ�^2=d1����@��� imR�[�h�0���]�KY5��|�5�9�3�Ps�7�
�x�d��ң�\�������<~��L����M\���HY�#P�ǭ�x��ņ>yx��ha?�/�8�3����Q�^/��)�Gk��1DG�K���L��ƶ�P{���|p���Z6<C�D��1>���^�-���nڍ.~p!�G�2�N0�7�[��NCw`�JK��=ƿ�mK!����������\�<*[ZZ�s�w�>�=�X�Zp<�Z�}�<Z^�\�o�J�#&�L���ᶁ=)�@k����iV�L:��˂�r-�����[���"�/�>>�V�3՜cϊr5�K�D=G`j|��@e��j{z0��6_�0|0���l�0�?�R�UҊ<@�<�o(�<�i��Fed|�l�ۉq���s�A�с�9Sd�z6�����&�+漙)��ݤ-ۻ����/6����1�?4��(W�?���y��?p�G�a��(.
���O//�!�`�;�׾9������ܱw�'�"�x	�' ��~]1�{G�u�Z�s�u��-�5�JE��� Q���N����*�XN�, '�����~�� w��E�ˋ$F��D48�������p	>�8:�,���%~����T�����M����p��_����o Yb�\���Sߵ�T������Љ8�����y4��w�I��6�����f�Q�ڙ!Ҳ���?���Z� ٿ��ŷ�LBIEV�򤸷�{׹B�G�1/�n��R��� b��6.�rF�6�η�'9�P�g�:�y�z��XvS�j��Ag~2ɋ�f�(��+���lݾsl4�\J7V"T���F���z)����'�"���B�A-F�d��]��j�y���z=u�~��N�&�waqx/Q�e�QE'	!�!��NY�'''��RVz F�%M�/���rT��?�M�)8�ڑ!(�v�T2���{�����O��-���5/��|�rخ�Ð'�N,g�_U�(Y3"Ζ���^��\hUTN��W���4*K%��}�\���!�vk\&��b�L����r��O{���;g>��2����ם����?e9�{����c�\������I^��&���/0���A fڐ�����i���y���������-Rm��ؼ��7^����⏰�Es�T��1��+�<Y��iN�)U�&
$��@��b^z셻Y�ӷQ���0��%��Q�Cl�P
�P�r�		߷:�(h9!Q�{:I�Ep���@��� F�Wh�31M��D�0�)���E��5H�c��hbbr���iʅ��4���q���.�
�Z\��ؙ�I��U��J��"�y	���[:y������㾚p� �bnIJª�k�9'vL�`����N�7���<���"h,~��|V����s���.�v�n�R{(��\P��g��k��
c��]�.I�gFHBՀ�[J]6��'��ܡ/m�U �X�y��%G��;&J)�>d-_\'���"0�%����>&��;e��5�A��.	���P'����F�6�
��+e��X}��?����a[�m9��C��Y����j���G��-Nh�T�L��>jIU��K�;^M��p1��k1���vS�����㣅6�s�]^_�~�V��)�Pk��U�]����]�>)H�_�N9�$oAy�W3�9�� -X���N�;��3\pn>�/����Z��I���v��#��fu��w|��1�`ЕSK��@a���
pTC	L���`I?U��i�¶��(sT�����~�j���#=t�S����& ��YT���7�%�m"��M�����ц��	����١?�>i1�sO�t{��2@����������Z&!9�v��BG�������k�(9t<�NHΡ߿jD}rf��E����vxؚ7�^����8��h�*��k`vS?L�/�����_\.tBu�v��־�@�q�W��:�I�P�zzz��X�Ȃ��c�(Ra���{%;�NON�\�*�G���}n��qU�NW��@14��� ����5s��"����A^���y�ؗD��Ӣ���8ȥA�|b��P����_>�?zhzs7QJ�U���������F�eЮ�B%�m_(���Y��G�7x��k�'
��zC*���� z�_Jb"���zߝ���?���K\7 �X��Uϖ��k�d����*���I_R��_�w;�n%D��a���N�Ʋe�+�2���ޑ����U.?��2��F�����-��v���%�����uY�Pc��X��pH���Zgv�c�Z��!�7�_�-S���R�����:a�戥q�v#F��=�`�kZ��\��i����i��f��)O^�9�=��[ߝ,J���6��n@%yV���Kl�����.:�w���ވ�w?@��c�Rg��RI\iM���Ҍ�S�Mĸ�[�H��M�s��,��3bk{"=�w��f��-���y g⊑S�/8����7���@FJJh��ɉ����Tddd_v�AiQkw��=]�=����;��E�-S�ߪ��'���j��/�L�T�k�~���#����Y��ԻDn� x:Q�e�z,B�sE!Q�Z�S��/q�G��Z�	,wOpQ~iE{�XF�l�M��'����5eJ��g��q�������0C��A�4_������p�F9U�jiz�,q�~A���;ބ֝�d���=��^�ф��[��w��&}�e�%�2���+.;Vo�ϲ��0>������p{��n�k�]���Uj���CfN�[�Ǒ�}m���L��ZZx0�� V�&��˵:U�p�ɗ��}�V��A�2�,=����v�4�q�p�aHO��];��l6��\)�D���`�4���H��f�㟔4�G-���@=��O���g�+@� �{�{��ԁU9��J�I%��\+��p���B�?=O�����*�4�dsb�!���/#��V{�E�8v��.�؛&x�V�=���F��RM�w."�Ǉ��E�ZrNת����}��h���{,xb�6�fF�r1J(�Dhtk6�ёܤ#=s� zu'9�- qH��j���M�Lt���Y�C1����/��@��ݏ1㽉d�G��&B./�8�>�'_b<h�T�ǖ���%�N�Ƒ�nv�&�iV���z&�X��o��H�E��m�~Y��-��י@W��C������?Q8�O�������= U8���h��5!�U��s:֢k��"<3��[e[���"z�,��l%��}
��8�Ĵ��}�əM	i�4�k4Z�ߞ,*��\��TJ9H��/�x��Q�^��X�A�k(xq�
*��9,0#}�J�	�㻝9����[H['���J=К�\�68p^݁�a�m�El��im�]uծ��T��kUNr����K�;�Ƽ�{;w�U�t�k�H����4+��9%�=��!!�V���sࢼ�]����p��!��aBk|�Nb(����Q��]��aFE�0Q�Eߖ���w�⣋�}�5on�Z<z�K�V%�1�ZLdp�8��7��IEī�_,؀>�A{�|e�?��qW�i{�x��`e�H8Ƃ�؊@���G���{��� k��<��Z�q�o@";{�L��r�Y�Q"��Q��|؏]-������1��܄�>��]�����~R���f�:��]<�H�]R�!���:���,`d����v�;{�PD�޸�&	�G<�!h	^�dF�ڏ��Jg�0�g���seD�V@ls����Z���n������O���8h"۰#����?s��-}���r���+a�xńb��]����nO���R!���勏��ɏGЁ��!>z��D��ۏ�dz����t�O^D�mx���OVgF��oe[�����#箭�X3�%S���`*�\���.��{SJ���X=�m��T��\_+��%�991d��-x������D��Z/+����d5ٿ�S��n���Մ]�˧���,nx�9z���Y&��E�J'�D�@�F�:=��/���<>Q8ڵ.ۈ�*�U}9YپקrUTrq�j*�D_���u�іԄ�2ҍ#�p��Y��*�4�X����DSOHk��V\�]]$C��9L�vTG�Ѽ)��v����*c�A^@�a֩B�4k���w�����$�O���˟L��H�\o���ܫ��2[�sKZ�e�E����qp�<Շ�H�$%�^�q��������Ɗ��Zr�?���H�|L�/���	��Z������O_?Bd3��78��4Q���d��h��v��e�{�ofV�������ܘCnЬ��)iεEo��Tc,8�!�dHY���SO�'�Y�e�A:@Ve�B�5^멯v� �YL�i(�Q+wq-�b�ߊor�{ɌfX���dldqK�jp~U�;�����Oj�O1���O�������,���D{�a�"Z�#��K�<��X>����E��!!�
T�\�U��ot|�i6�?z�X$�ux�-�Erl�$��Lϰ��!��wžWH��ۈ���o��Z �Y�o���)Ō+H�m�2?+8�A���l���}��b�߷��dtQ�ml"����v�z��~Taq��t��c�8�&Rz�Ԅ����*���sjs[��_6�X�+sy�u8U�vN����/m!a8�.C�T�a�>�F�a�ܼr�Y-����E0�k����&�S��]X�IW�ff������{ݹ�~�/�`�w_?1��&�ڭ��>�:��7�=��_k�?n���(����>\J�T �&8{B��E�.b�1~��'���o���_�?run��%�԰��������������nPi)�e�[3���%��0�_��T��X;c��{���:^�I�|+@��;�tJ�S�؍N�Ρq߈6��"��	�!.S�k(�E��L��I���7��C��?6xZ�/R��5��Q���P�"�9Rm��cS���|�Q G�N�~7H���^ȣI��A:�?��R`F��-�� ���f�V�]$�&|�Z�M�	�`�~�3e�ꠥ�"c��"m��F�a?猡��-:���Ai�c�QL���`;u���7-�W�OHܷL��ߤ���^0m�{��7�@�'lW�|�&l�L����s����u��y�����i��vv�J����P��
�M�?�M��%���D���Eɵ��ح�[�x��7�y�h�'�)Bh��!���ﰕ��X���gY��Ƕ�7���Hx6=/brZ:�n!�B
����K`��;����`���}���/�������lfϬ�)�65�]���'F�Ƕ�Ƒ�l�ԁ�%5�����Q�=t���K�[{����N6��~<�o#���s���{2����Џ�S[''/s�E�ɗ��������Ԥ��C`�n҄|��u�x�[A��?�����v!F?��0�)�Ճ�L��v#�ֆD�D���}�����I}�n��rQ`��؟Qy�xv�h3 �Be_�Z�d���'���;a��[X�eSSb���a��u,n�(Min��x���ؙ�nf�f��u�/�@·��R�S o��'�=�la��s��04������k&vJ4;y	��QqT;jTv	8�����|�]�"8AO����~��f��'3�*���2��	��D_�w�LA6����!���t�P)f�?lx�:���c2���%''w[�1� �8��&��3����'Td	��E�f��ly��V\s�;��,���_).=�{k�D^�O#v�샂�r�OSr��؏G�[v��N���[�a��u�67^��{K̶�)~����=��g�e�S�@��yW	&�T��J����p�~���ԩ̺D�c�����x�K����Sv��x:곦@���G+��������`бt��m��F��G��l��o��H��W���}�Mf���s������o�N��C,'	k�*J��H�>�<�&|&�o_@9c��$>��+�GR؄1,®�O��.�<Q ���A]��]�<��?PL-|i7�����r��A��e,M�`L�1f��$��/b7X;�bq��AWm��S@	� �ԅ6�8�u�W�;߻����v��T�3=�r:�~z[*^E;\�P�ͩ�2�d�(��/���͚���/�μi��e�_T��z/P�EY^C�X1;b,u5�n����*���c�<h��i�7�[[��g���g~~��xi1q�Q�5VRqeYfnG��	(?�-��l��(5@� ��`9.��%�n�)�?P�?�ꔅ ���U֤?^��@��H4ȫF+�wZ�e�����x]*��%��N����۹�6~�I�J�P���>���Q��	V��������F�j� x�M�d�ሸ�׊ܽ�	$G���r��B�_=*��>߱���Og#�����lu6o�\�X�V\�s���@�(��ehv*���0k�ՙ)dHݔ1Md��~���P�޴_�U��$w���B{�^2��d{�(X�~.(�sf�NzbCj�u�=�$R�/�b��� $wa �d|E��%ikF6o(=4^�
K�c^��G,�u����`_<��������A̯M&W��nJ(��1��=��F�)�����Y@��X5�j��ZkuvΚy?ȴ�W$>�� ��X�@	���<�Z��LLM9�#�D�(�>�+!�d�
j_;�Y]��7oX�5t�V�m�6��u��|��۵J� mY~�v�V>��of��	 )?�Zԙ{�5�,�K�ĩm�#g��5lM�A�m�	���ss<��������������FZ����Du;�Hzm��������i)UVBRI��R��h���w��ƫQ� #��V�PԂh*U��(�M�����Ѱ���w`"=��l�������(�R�v#�e4������tQ�)h0��z�̯�&�M��O5�����.�W{n�e�3���?XKŽM���`��UA������TZn����}��P�F���@l����g�Qt L3$�n�CnZ�0S���?��vt�6�ZcE���¼�$[�x��C��Β��)�r_�#���� ��.d4^���{�
�~�>B���Ztӡ�	��G�9�G�^~{��j���B8$�9��A�	�j����vѰ�}��B*T��õ����PX�)�̎��K"1�Z��mA�R��������Q�q���ߙY�Z�&�3��`ہ���V��bޞ�92���#Oi���ڤ{������n�X%8�����53�y��R��JL^<�^��׳�?q�|����tgv��3�/�.@��k�~�fM�x�X�W��$Q�ܐ���;��٬�_ A%@��c���rJ����Y�.;�����^^]�Vj7���V_,�A�6�̓K��:А�Џ�a�����>k@zQ��S�"��kWKI���Ǉ��	-<~%X��_.���F@)�|䣘��x�s�\��ωJYPY���2TL
$�����:4�G��H?���sD��$WדSO�-\�����,���͖<�Τ�q�0�f]��H+��qC�L����q��ܸ��&ά�׾�4T�gS?���)0����jN���iD�!nh?8:���|��+�(�oJ��D�ɹ�|!pG~��g��q�{O��2�J���=(ڴ�a���^7�%�q6����~_�:i��c�f�ަ��~�$"�q��0yr8��[c�rRwU�Hb��4^V ����;�V����������g9F�������M`�<�r�⾷_]7�e�F,�p�� �N\Ĉc�˵�N�qN�Qc a����'@4ɬN4���W�k4�6<������&����2����b9@�ju0�q)�q�2���m����^_������\-�+ �?��K?�zp^����`O�B�N�U����&ڷ��-Rg�w��k�2���w�O8��5z����Cm�ϱ���B 7E[�e��XλX���,�y�H*	�!��	s�q*�LO��k�j���h-*��BT9��{~g]2��ed����v���K�H�����Cߐ�5V�J����D�Oc�P���N��X�Zr��#8�Ā]�������4���@���.pօ�0�R�-��΁=�p������@��_f�xA�f���߰1|�P3�3���)��}U��ZB��>V���_f���Z��>+��z���2� Y�*C���m��}�j5yr���"�?�s�XR^��W�q!������{�mF����KȪ��QArq����4^g*�����&��|���V14l?��� �F�@��y�X!h0ߗ���̆<U[�|����mk�1>�j��3��	�S �y��1F��i7)��o�;!�#�,6�M����ߍ-��B���-���]�X��D&e�9Q	U0m��.�GR�&m\_��,��i�`H���r��`BS
��Lȿ[S1n�e�M�t�D`���b��Ӑ�Nʇ~_��
b�[�1�k��5<�B��hޘ_��^�;����(��v�6J�e�RH��L�R����R����l>��'�g�{��/�8,� ���I�/�Y'"!i8r+�NK|����ٝj?��0�}���ރlP�W�M��xv���\=R�Of��/Z�*\�0��<�>��=I�&2{ϗlM�y�����Ct:�\���5���s�*%��e2(c�w]�H���疣��>b>KA���E����_�ymE���4[�W���/�z�\6xǋ55�@�����|b���
Z��5��H��ƿ̂���&�)�2��}NBw�8�-�L^�2�KxwyG�z�jlA?TlC7��l���qiT;���xZ�7�9�g4�;��S���r���U�^���QkJ;4�:ވKaL����+�� |�^��(t�V3���g�f� D�쒊��!�1T
�u5@bj^lTv���Q��X��KF�@f@I3O$�&挗I����B��m�Fݔ]ϋ���:S)d��X����w�B3�$�y(�^��(@���a=��9J ۧ.^_�^8*,��%$Xg���W�O��l2�����U6|򓓨�~�L��}~#[��F_4ջ�9�T��+-V���yz����@%�t�
6Վ�1D���O����q&�h��A� �]5���QJ�����B���������]�s�e�1�,�3���x1�� ��h�Y���z>�9ly�5��;}�����)K3�n����oi���D�n=�w%���1�G
nX��Xˇv�|���E��3��d@��w�b/����ou �ZPh ��e�6�H����V7�R��s8�qrG\�͖;r,]��B��q�n��,B����c��2�%i�o��:*n���{o޻�rޜ�;Fx����!�{_��c	S�(ccn�(C�ﻲ6R������4{Є_a��{�a��#�������ԶV�{�T�������7����)�4Z�R��~�]mjlrړ^ksEv�L�(���|��طo�bN�X7x��	J}G����<"� QmǙ��f߂�jC!�F�F�wkT	�*������Y:����<��u�"�,����/���ȟ�bĞ�ořɸޚ����-G��6<�%�d�:7���1���^�*~�]|;�0�x��9�8
t��Z݂;�� �N���j�!�8^@�:sw4���� �>ݰ���u:T���S������s~��o]�c�o���=��/M-1�GWߜC��\� ���O&O��"��8Ȩ7���%m��D����{�F���	���H����na�����N��Y\�
O]Τ�p�'�j�u�O��[^����e�Õ|�i���3��.���U�g[�l�P�#@t�m�~��}�e�ub���Dk���Z�������;�6g~��5bp�Y� ܨ���@uR>��DT�Y��@��{�����v°B�#�m�{�P�? �j���ֿB�b-���:���Rl�r	Ņ�T�Ȉ�j��j�`�4�����Uq���<�'5.m<�S���<�B*�h�ls�|y7�T��F-��l�1��S���+/@_?��j9����Y'��-_�2g!併���d��Q��U[�6��l��E�v+�{=�MgP�B G���S[����N��D��m[���3'��j��&܉϶��!��	7�u#�N��-j��
�^�LE�������qG�������]������|�����ͥ4�b��pf���/��%J�q��S������Y�;��&$,���5��&Ix{2^�&q�4��Z�˞���*]# 3�LO�/Z����	�[��.u��(.�Dmb�F{$�v������-In��x/)�yɋv��O�-;��W�����h�����ubb!o��*~��::�V@- G$.q����#5+����Sv�KD��;v$�`N���0�\���.�h	T�|�HE'�U8���)�&*�D/dO�%�MY�	=S́J������(y������u�� �L'�7W&20B�	�rh�sm����ّ��a�@�?�8����|8�~w�Xڳ�&��;
�<��K��C�X	��;��p��c�|mj�&G���mT�7)��g�.W��W�:`:�ErW��ӝ<���g��!D��'am��Mk��Ԟ���t����B�*����7tq�(����Z�~�(�+ܶ�� 9�v�~�ÍA�%���p,*�<
KJV�Q����ٍY�8���e�äZLR-Q!�:��߆F6H�9��9RXx��߿��$��������(<{�����2<S�Vп��pل���$0���9�BѕeP�	v=�	#E-��r�&N��DT�~%��X�K�?*Ƥ�w����wE��rB�a��z.��g�dV���[)썘j�j�Е� J���7�w^� ���2���,ԓ�eEv�L�r(����DJ�&1���ƍ{��ŧC;\h������l��0� M��503Ȱ�윜!iř�Y��X�)��l�nn�;<n�Ϋ�ѩ��v����X �zPPPK�~����yڍ&p����?9��v�^;p�Z���|�7���zߒ��\E6g�7{����K����T��P(߅7섻��3>����/F�x��;W���۫e��@���!2jpʙX�ӥq���\�y9 ��+O����ƚ?�HBK�Z�1>]np^�!"!���I��5��[:PG�ˋ�Z,��??�o�'RXM-�	�g���?��ۢ�xS&,���/?��:o��?lp�`��ܣ��+����� 84SeL�ǵX
9�+��>=����H�e�S��xt��������b�<���.:0����x���>np��K!ӆD�Ժ�;5�W�F�w�'R��OxA�Q���C���R䵸���~��b�	`q�@p�����0�gG��%��xV��,���8є�P��4�-u�@a��FP�vIU�!f�s���������m��h��Q��,26�y%>;�ЩV��v-��A���L����[)===���S���4�0������s��)g�&���j^�T��sK]�J����:)?g�%C���U��p�1Dh�`1���W��~[��:x�q)ew�j}n��ۍŞ�Pc$�W�!��SÙ}^z��1�x���Cr�$ٰR���H�"���0�%>���Ȃè���	$���@$��J �a�Ox8R't�@O/������+�J���#U�=<>p������+���֣H�|D�VS��A��6z�.P��S�*0�it�H�hu67�v5g�����es���_1#����g�[@)����Ô!E����I��
%�@W�ͷ�y�{>��Qjb9��r�?������,n��Q�%��
An����!����}���ik�L�����}9ɵ�9`����zY�=7E]4\�-�|y����E](���I;�Pg8�p����$Z������ Œ��4Z-��J�7�O���`�\��2H�%X?,�øU�)|�t�h6.��R~#�z,�VC	u�w�EYh��E�M�ڼ�R��H&~�� ���iE�m-L=��m_d��T�W�rd�<4���㼮RM!�sE��RIK�_�p��v�7}�/�ʴ���̇�W�?_�Ln����W�[��0�(�C=��:�22�S���߃�����v�c����9�?�y2������|��H%k�8��1
3�%�c��(m�ȂJ�U��J���~�T;��؄ƥ����R��8� ����K���'A���D�S�(9t	�k�uPߒY:�ݘr>e��og���WGI�G�$�fbE�J�q�q�~�=o�7�1�\.ʮS�ճ�¯p�� 'y����E��sZGBIm�*��Ԟ`�X�{���1,���7�W/Ғ��ֽ��&�S������b��O��b&�e���7�65�T��9�ޏ�6�e6"���p�]$Ȳ�	��g{/�(V2�&�͞��6�m��L:�&�;tX���	~=�s%_�<T����Tt�����6oZ�^e�@H+���0ܞJ��Lg~�e=|ټ�.O��0hAK�4����ُ��Wl{���%������Ki�ɰ=�o"��s�����nF�]̃��Շuwgp��|���E&�7�k��Ռ��c��X��f������#嫐�w3e��Ǉ�.���7�~����"4%�P�@\C��h��?��݃i"�~f�
�t��*�l�{��-a��\�3�'��)dT�_���ki����0�R&��tE�s��v�����n�e0�Q�׈1��[ⶁ��?&�&W������u�O�-�������g���_�@��&��l��"D��b9Y	������7`�k-�h̛B6�}�~��B	WKA��D�(�,��j0C����n��l?�os	��x�KT�/L�@|t���]���g*8r�<�8j:X���C�6u�^9ee�����w[뻍���˯�*V�|(C��5{�]|�
�(�Otd�;����?L|�1��^�[��n��Hȼ���9� ݤ�����_"Ƞ��W�r})o���@�i��M4����P 4���o�	R��\���j
�.�(B�Z������V�[U��� <��OZ�eWP_/PR�]gQ�]���wڲv	=�N����N$�P�7c�`Azu�C�fo�����ޔҨv��Ο�^�<��@}9#8���=��;�m�w�*5:uk���q]u��������9�gF-�9��ش�^r��:��yĀ
P��?��1:���:N&Fc�ic4�m�ml۶��Vc�M�ƶm'������f%s�u_��g�C��K�r=ް��O��.!�@��iȪh�M1�����@���}ƌcUb��!���k���D�����,�ʣCEn^Ұ����T��|��[�3��Wt!����|ۍ.�ꋥ�
����dBp��S!E*S�R�.���|M���T4y�����2���U��oxyx��l4���l�tk��S���1ȸCfF�Lq�;���S/*|k�>�O7���l*TD��4�E%�gl׸�暙���q��M�%碇ͯ��CEQY��=��l�gY!'�_kw�3�@��im��z  5�Y��?����z�a�긐TU1aX�Hf���5���b�dA(����@��itA\]�:Ԓ����!�Z��`j��f~�_ae޶�u����=� ^홑�������f������wω��]��L��V��@�Z��z�V^�-�0����h�M��r�Q4� �d82w~X섘�n �nc6���
���ꚩ���V�
�~������(�*��H�	���1s�����P������L��GAӃ�d/Uُ�4�D*���4�/�Nχ�Zj!8E�Tz]F�?��Xb�N�}���H@V���G�\C�'����h��W
x��	��Q�:>b�7�@NY���c���u�C�΋r*c�X�p���0��QI!≵-;�ë8w�(7�;\����|�DǑm{�
��(�-|�t�%%����v�u	:����/���h{xp}�I���"��=R���d��u9���@�����#�
�`�}����:��ȣ���c�+�/�oŻ�NKQ�{�?�8}_c�Yi�Vr�bX}TB�?z�q��WvOA�b�J�)��8q^h���<�w>EW}Zʀ~0�� T{��Sj���/:���ү���en�[�lvfo�����Y�5�ES��X=\�)c��O����g�5L�4�Ը\���?J�t���r��s~�ʼ�Ī��wz��Y+�l`��~c��@��]���n9��g�L��U0l��k"��Z5�l�E�ѓg�f��:�ܢq��A�^�Kc�]�Q�������������Z�*����l�S<�C[��l$f9~@,�L6b�;���g�i<S��I��j���!�H�e�&)�]K�/��
�c��L���d�(�`Gɳ4�ս�s {������������ˋ��#rS�&0�C������J��s��π���J(<�T���^����Q���h���N1��k�	�xi+p�[�֝�_�Ua�:���%���;�C]B���|%/"�e;\����g�����Tm��Op�/�j�c�"��1)�֞I���m�`�3t�;&>�D�-��Mvj�1MF�#��%I;۽B!P�鱎�.l�{��-��?�� �8b9q��`��F]i5	>z��X�3z��~�2pp=}�G\Y:C}�0`5fA|�����q����Y��B��tQ�^�!x�p��pf�E�ݴ����d7Y�K�l1��igT�\>I���[�Lz@0�O��z�*���qaT(���-�} `֪Ui���8r���#�1B�7 ���
��	������f2���*:ђ']-���2O
�Q<���\��]�sF��s�z`~o�o�r5!���9̥�g�����ۢ^�c������[R�Q��?�
{��?<�Ɨ��I�SPP�03���=3�%2�1~L�D��~!� � �/��
���%�oׂ�^A�lд̟K�KsѦ�p�nϳ�	�Q�82�X=.�(��>�K	��J�7p<BZa?�,zq,nG���4<�D��8�8/��2��[g�g���7a�|0ĸ���`�����U��ɪ�SL���}�ne�.��K�v]u��w����s~�SӋ�h���p���x��A<������I���YX_rY$Sk��o-�Hw�{LK��� e+ȅGgp7�����Q�O��(K��6��q�e1৖\���D�����x}�~ха���v�@J�+��d��r�H��R���AE���׭O�x�J�������UL;�%�ӧ��r�=��Ǐu��zi��	�d�m�o�BM��+��)��Qgw'S���m]L�2Ņ���x��6�0�%��	\Q�v �`o����}<��y����A��ú�"��`tevUN��b�7
�9<<�e�=G\E��SN�Rj���m�fo��N���qq� ��t�ܗ�Z��Wy�I�D:��!�����͊&����Mj��v<�ɺ�W6�ykP{� $�s��I��������������55d%������t&��h�uj��׻e�ލ�m��{��y���Ucm�z�-�l����g��}��W��oCȱ��c���jB���ڷ�|��z���_]�6����-X�/Lo�cw�B�'ӣS����p`
Ģ�&��S��%��.SV6��у������[�$���
NlMs�ÑŽ����\2���gg����G�0ҹ�"Li7άo�1�ҋ�l%��k
�8B\�ڙ���38-R��Y:��������ʼ>�h�-���B�J��:8^
�h)S�3C7<��1�z� a7�d�q5Ē�b��/�1i-��a��h|�5�<Q�}2���O �(���g�mTvI���[� �Z�Z�%}$Py��Z�U3c���+"����1EZ��2!1�(52u���s~S�O%e���2s�^�����~Hz�qi��m��;���E�c�����U��f�7�]��k�
�%� �^6%T�s�l5����{�K����nt��ĘYl,�6)Ml���d�_$*�77l����z8�+����v�b�Vף���^��J�8(�����b�w�Q@nZy���>C/FZo�ཤ��������Z�X��*��A�OOu�����j��v����8���j`����;�E�7��Dud|%��H�����Α�yT��-?;{�&�����S�HMCׁ�h ���vG������#�?C���3�7�/x�jx��e%?��p�$D(�_�1�]ä�oy�#�{/�q���s1�DÞO衔������Ǖ��.�.+����q-p@B;��-�-}�Ȳ�\�tkl�W���澹ݵ�	1w��g����޻�]�x�Հ��932�Rs[E�7�<W��&���M3��;j��ugP8�.&���u�K�(!8���{�G5�q
�[8����o�9�c�-5M5U�v��S@��;8_��_������U��3IIIv��L8R��R���3|؉��� ���vMH��9z;��K�a9~��^މ�|�ֻ�Ɓ�!�j��C�����)�(�)�R=�r�mT��d�D-(j����ܗ��n�ӹ�fo��3s�B)����:-~_��I�W�M��eϭW��@�Sw�CF�C�ۓ��ၡ!2f�����=���⧐M�.!�	;�[��L��*�m^��R��N��h�� Ru���o�@]J���:ףj-:
��\֭�E�I;��� #Ӱ����߳�{�:�����t?�y׈�8jE���y}��>i���;��l(7��e�������&:)\kc"�U���@n G+�|/\|b����T�gOm�r4W�9�=l������(l�4=Rw8֡�%l�(�k����{�?v��`r��N�[�">�H�l��F��Q��\yǫ>�`��u!�|�Y�si��&@����Ձ����i5��l���~�㩋���Δ�G�� ��Z����ۿ�[�w}V��`a&���tZ�x��R=T�/!p><�=?t�k���������*���K�N����f�#I�Qj
zl�S�����ᤙi|K�9���I'R~𮽬ŝI};������g8��l.g����4v["��䝡���PXP1�pp����F�S�%�<<ʳZ�m������D\Nb:Ez���0�z+��D�����mQN -�p
��CLM �⻲����J��p~G@E�.��z���ϴR��D[�	��?]��>Q�/^'�s1Ķ�	�J.w�|����[��^�u���4�#ƻ4ȓ�������B����C?Ǧ<~ۊFx��ؾ�R�5�Tk��n�������<^0T:��'N^�a����p.U6c�4#n׬:)��� �l?j�N�<Mܠ��]��޶'H�QW�j���UJ���I5SD�L��?��t/��w+�C�H�OG)GS�^���<H��)|�����X��\�R���m�N�v�W}��C����m���f�$���Bc&��ͬ� ه��ֺ�`�wظ���$]],1+Gc�ܪ l�T�uF �6�w��Ƴ�.���b����"#����&�g��qc�x8��1&�VA��(0��=�h��ּ|��/�?�	�J��Ў/����{9�:���&��Q�X�7���E�s��E��l]��.G�U%�;�1.LQ��O�R���W��$����|/�mK�m��(�4c3�|Թnl)�-�tۦ�����/�*�g,'Êӭm�m/��7 �7����Z��n�L��-��!���w0������/����%!M�H��N��<p���v<X�H��q�yΙ������}&����q(�:RɁw�X�S�}/Y+qE>�ÿ$�'#a�pz��.n>���x<�r�}<�2�xGzU�D�S!��V�!�n�m�� LF��h���řr�@ꡐS���5��P�t��&�/$��������:9�9���?��!�z�yڋ��AGp���2f����؏.�>�o�|��� �aU�x�o����֓�b���u���6�����3���*��Re����r�ړ
��yƇ�Zoǅ#�D��`�+������*�j�Z���]�T��@�1�~2��L��y�.�G�>|O� ��@8������/z�w���Z�w���']�yA�k��3��3�W���4o\��[n���w-�~ s�'<H�q�*�W{��L�	G�w��NQ�(�FeW�Q��.�>��C�ܗ��؇��"�{{{�׻�-v[�L�CQ��]p1��A�mJ�M����FcI_�V��̯�&�0Ep��*!�$�}��v�g;������Ð]�/VόǬ�W�[�����	 $�?�g7����t[�����:�rv8:����ᗋo���H'��x���v[���#�:Г������߫)��'�tlΊf�.�=/^]w�Q��o=xA�r�:���pzn[�*j����E9��
{$1y�������1���~B���`g��[���s�H\-�AHF��v\�I��N��S^[Q-���h�,[��b#A_qO�1T�,�W�^�����Ss�|<64�vA�Jm�ց����Vn����s���9���2cAC���>n���S�G��anj�x�X�>�N����S=f��Jq��3�N�LD�Pcm^q���Tc&m��YȘ!} k67��_��b��z�n$jG�#��8wl-"٘R/�ṻ���:��dy� 睉����Z��%��:P�������a�HT�����O�:�����<s%��c���*���-C�!O�p-�����a�w� ���x��n}^c���N>��ǒP5��/�etK|��ǃre�� �M��Ve�s����<+��G
�F�#]/Q*ct>VYuۉ�V(1
��S�>��J�N:�������8��O��z�ƭ��Ms4��O�\�p�n��؏h���A̚,�u�Zy��Ŷ��Ƹ�xI]�!�:"$!.�рf�>�X���1�'�f��s�i^p4��6dT�Waoj�(<V��bY�)�L)�0���୳�j�V�.o��%ӯ���ѶG��{��0�oܭo�~�لGh�@�
��i�s��-�u;*ن�Y?6y"��hA㺟:���Z���Ӹ_%�B��%掸�~���7`x�,�+��v\�8�����]
���=c���D�֛\i}}�wJ��9{��ok"���9����Ϫɐ���!?��s�U ���[����s|�t(l�K����P��S"��x�����WG�}ڕ�moM;����Ӭ�-1�\bմ�w�ݹ�ͣg:Ϩf��/�.�~�7܋|���g���sz��%C��4D��0ԓg�-ֵ�'���wV���<�O�ŀo�W`��m���^lJ�u�H:T�����F0S��?�͍���0����ѩ����9��r|+wE�u�ޅ}���C�nT;��{	u�2X���༄!}�x5�^d̖{�Jޞ�+jb��6�!��L����<�?���}2��..������ ���*?8|��j2za�����2�O�I�$ed^.�c��>�7�n�`�{�aEF���-�u��*I��Q��U��_��.G�%�I#K���̈́�g�-��{����}{��&���_'�L:����q�d	/���W34�.�(GۊRn���W����ˡ|fGW����{�ߜ8�:����7�q��3Yz�Xi��5FFf�aם��,�MO8�5d����[���&�L8פ\���Iw�������2�"���q:�a)W8%>�Q���=:&O�B��yA�L�N`��*��JR5��&�㑢T��c�$_� ��}�����%w识�٬+�������0��e�|���+״]�[柼� ��-!�O\{F,\��}�vn�?@{���/�؅�X����a��hp��NSCg��������8�\<.==��>��<��BB��;<!���9��@z�-��sB�P�~��K�rҡ@3vYe���g���n��Q�m�ۈ$F�h�IW�n�*��m|߶ª~$3B��" �����SN�0�aéQ��T�>R���1ď�a���,���Bn�T��`l�������F ��ZR�!��w��BMQ,�O"њP����:�������A�/A�B���N�]�5� �P�s�	h�|�Â�?�ҡb����ioTS��Ȏ���`P�߰��;��<����;�;���k���[|<vx�e��-7�;��������ͣ�4��$9��`�\�U\~�k �
9��J��Y�V�8ƈߌ��ݬȳ�S�Q3u���Z��@Q���s����/	xN9 �m����=�!7r���Ѵ'�*}s�I�K�%�_@���Xh��o�h�͵)�s��eڝv�'8�]:j�{swE��l��e6��+e�c��O���	a-�ݛ�dfZ�I�8#�bU���Z�INȠ��A��7^���M,
)��Z���:�@n���U}������f�"�.�7뷺��!�d��@�:�J-�
��_`�JQ�q�h�3�Q|G��/�2a�^�j��t��0�0%�!���ج񀧿� ��tp`M��K5�?[	5�)Vd��`�
���V���V{����(��V�r� �Bt��`��~V�y��A])��q��h�\I������0��,'�WC׼f�������X���[J;<ov��^;��D1�L���� ����u�_�P�i��D�����z�i�	(�5~�������(�BBҌFp2���<�tO�su�ad�b�J��)������9T��:��Y���GlIݱ�����҂U��<l g�ǲ\�B�}9(y�L�R�?qu�B҆�ӓ�U�)����w6$�$1T�Z�:�WoOA�5R�Й���7��5v���mC;b�&���n��U�p4��N���J���t�IkJ�%7��LV&_���lb����K��4��!����K[KE�p`�r=����|�f)>䌖���O�=ך�����q0 ��hG�����[���2�5#˒]��6Q�O�Si��s�����]�jȑ�wU��	�9���B���=�N�s�1�O���y��M��*r彏�@J�ǡ2�o�:�4*r����ˇ<�?�e^�h��cU���9�S��?�H�����m�Xwǝ�~//1?&�[S_l(�>CW�º�P$������}"�v�mn���������|�^L�_t� 뚎k����&��͆�[fx�4 ��.t�8m-}��ߡ���F����7[dЉG
�$%{w�?�RK&��R&�]���I AM�HZ �!���Jm�5xd�n��$��X��w��&E�qN�Ӄs��G"��'�}`~>6>~5�2jg>\i��6��ϴݾ[�WSKq�����ؿ�K<���/�����E�Í���hm��?�,d������U��?\�P��[w ��],:�:ƹ�6W\;�$�㩅d�1�%�<,T��ц����֑4;�r.^w��� �`����|+d􀸙��@��m�;P�4g ����;v�c��/���$�VE�����sDV:صW��	:jX6���2�g�����n|THa�����l���w]@|;W�k����f��.H�f�ʌ�8[#�?_Ȝ����VnsV`A�o�����,P< �Q��c�B|�Ed;��!N��e[ސ��Rk���V0oMK�A�1����}����ߤeA�o�!���@�v|����ホ��T�$�pN��R��3��w}�K����Mύ��@��g*��Ɇ�_l���Qt�>����4��l���P�,��L���H�L�.�#�[r�/��-	
f�@�th�~���&��ה\<f`F�_ג��������t��t�A7y�����G�����u��ұuQ��8�e��]�7�-��Y���]��k��	�j��/L�LHHS}��诤�(@Z��T���Ô"�@ۂ��B�o���oH'B݅
S�#����W��i�OJ����e��M�7��Ŋ�4>o�L�K�(�"��.O��0'E</:C1i�ܘ��	Orcq$����G��U�o�E+��.=j�L�^��/U�0�&��U��*Z�j5&:�*Q��5U���"��=��
�e�g�x��sX���)�,D�(ٺ�T�y���y�\K��n�3��`Q�pl�4�����k�ޥ��Vx��*f�z��!��/�Æ��/>��Ua���g]'Cv���Mˣ=#��H���H��v����pb��[�`�v��2!k�l�-���e�v�Լ�]��PU�"?�tqr:�7��8��t�x[��i���������؊��Ҥ�_�
WϺ�ǅ�����ޣ�]���h�l�>2d5�!�C/�|*���_��A]`6Sm1`N��\�vݟ�F[��N7���_v��I������7�d'���:X�[��
������*.�
I��^��.����G����z�5H�%�Q+�iغG�
��':|M��+fɅ};���yC�fO�?�����ȑ�Y�>�/�x�ƙ�7��
�e�:-��rl8D%9/C;���7�SޙyI�����Y��F���r�mw���KA�������K$�s���Aɔ��j�86�AS�O�s)ȃ�h����,�iKJ�	��4.�+j�^\>��%��F��)�h�:�'��9ܱ���n�܊��Vp.���
���Ū��d;��`���?W�GJ׾���坹���Z��Du!M�� �0l/X�_հ���tla�!C�7Z%�R�y��$���4�o��΁8���^����[���:�0)�+�ӱ��ƚbf�q�5��P��Uk^9\ ��MҕT8�5�B���;9;X?e#���끂�8U�b̮e��:������O�OT��	�J���9�O��;k�,�$獒0|�E�2�c4GF�`��q+?��
"�����nFx��`uV�U�Ç��Zm�L����Y1���4D�@�|ݩ��o���q��fS��,�٫�>�|٧�C�MT?r/8��̛w`�m��t�����P={"A����F&&�4e�W[�%��N��Y����#o���X%Uw�������I��&�(l�"�jӚ�Hǒ�aϕ����Ld���05�O!<P��~}(���k��]���5*��ᾚ�����,X8}8_p�G"]|�vX�|�V�C�W4F3Ո!�N�d�A�����<9���΋��Tzݾ�2���Y/���ް���ۣE��c��������W�|����*J��M���������(kT�M�����S�ϛ��3���J֥=gR�B�Am�7[�e6	�Y~\�c�`���s%���9�nj�[_���)SA+
�^�c�L-�ꈡ��KVV-А�Mr3�3P���נ���G��,93����`���W��ͽ��
�p�'֦�ưkz�;9���D0Iy]l'�?{�s���z31���8w��/a���W�_[��Y��S�����a����pC1�(LP���/Jq�������f0�scE��<���ݒ$<v#�c�IM�1��-�����O��Z^�|O~�S�ܸ@r���+��T���ф�p%�;�3T�.u���;G�!��﫳A+���
���;�'�[:����\�&\T�������.�TsBU�]�w��N/��}�_��54$5�u����z�&P���\.���ԧ��d4p{G� QMMm{/U����su�+ ���U������3����Q�$ik�UP�=Ϫ��p�ԬK�"��i�B�����5��u��M�bbPm���Z��.>w`�nEヺ�@����5FRR�7�R�ombj�	t�a�x|^�,,�j�6�ə���z�����Ð��0g^���cvgk�Q�o[���L���(�9���W�[�Dq���֣7�\ӷGi���ʴၜ���0�W�˅#nA[� ��A�ik�'�����4�n F��v7�Wcw�"�v>�U{{��Z������kJ.oB�8d�fhRS�Ya*?�C���,ǽ�ay�8u�.�*��;�382�B���dժ>/�����D�>)�B"`Z�0y���U���ֳB5Uoj[�`�A�Rܓ���]wS��?���W�[���&�QB_��:eV�.~+7ѳi@���4^@��5f#I��c���u�/���<A��냡M�`�����Ѻ�YG�o���nH�������|-���ҟ�#UDf,�p����ө^P�(xx�Jv�� �L(���.H���^��$2"L�8��T�0]��+mQ�Ѕ¨�h4d�Mj�y����DKM���!�iι��Rt�l����q
���ƕ����1K'�V .>���n[P����&�"P�@>��B��f�w��k�l����j���`�\$���r�� ���Z�g���S!KV���PL6]�24�*Q͍�;�5��|
e��/L\�U�=��u-� O�e �>koy})����$M��jğ 7���`�Ex?8��t�A�~
����Myi�rM�X�^��<T�$#��*�YM�M�K�wx�F��la��a����A�'փI]E(�Y� ��??�RXM� pFw�J�����L�H0���ܧ�Qk���N�X��#���A8�&5�!�h�?��{ra�D$�ʤ���v��qxU�l]w�Ó� <bZ9Ct��p.o��j�N���n$�}:^)����؊�%!�8kw�	�&�����0��s��&nJr������û�H�\P��=Ǎz��؞쳓E&�c�؄�f|�YE%�Z�|<o���'���9k����٘����i/5��P�1�Ú+1�ϣam��wNNN���e���m�s@}g������saBԴV�����O�dxtɺz$�V�tJ �ԧ��t#���/!�F*$ �ZQ#5ð��BCˮ��&Z�P(�bY?�K�Xc�܉���W[Y@��E+Vu*Ҡ_2hhhiL�0\N�
'-�>πH,��/��?��V4�ϊ���v�П�X{9b{EBPbb:�X��~�߁�T�(�h�^w:蓲=��>3��1+��0B-<�D=�L��Mf��w]u�Ҵ��h	��;��(8"}O�ʞ��C?��LS�����hM��RAx+7I6?Tׅ�9��V~��ގe#�^î�P�{QӏlK!Ş=?e�HB���n�p �b�q����{�_zI%��NPt��oh��h�k����Pk ��t�ep���&�"�|�C:,AC��F���Նo.#_�>�췫� �[�ȧ�1��Z
ÿ�=���<���>�~��&Ў9]y���Ep0,iS�BEI)�4�f�D^���͂�����}H�A=ڥ���Aq���0�]*8�y��555�����8:>�����:�OG��	8bu:6��7}UP����)4
V�	�V�7K$�V_�w����;*��-
p�?햒P�A��2�N���E�������b0����vZ�h���^�v�EE����Ͽ ����2�Uh���Q3G�]Һ$�VP7����w,�҈���A��-M؜��ˡ`�;�+�̪6}$b��9��x�8J8C-t�h�է�g��w��'�*B�� K�/�]�o�>���6�=�����T�7T>� �Z��go����y";ɒ�_-�X�q��[�{z�'�ky�4X��&�˺;�.��5�!�0�Vs�a!$�3��^Br4���N�����1�Z_Ө?��*�h��Q�$T��E��D�qA�k�J#������c�Q2jt>/��M�S�q$Ta�x�|��/�����n�!�~�e���?��y�J�:-F�[�
��C"yy89��y�t01�ݻFU�HO��!V��0%��2��P��s�+6|=������+�����|ޗ[�Ġ�E#��WIAq�_��X~L��D�3���=��=���>:ſ�&4r�^���q�\�u@Z����w_v����Dn��8�A��9��JR��7�:�Ԅ����z�oV�|y8�ȮDM"��9,�]M:�^�Ɔ�x�,ܑ���!}��>o�p��1�o��Dny�X���� �D&�;u@��2�"�#7��5�D[K:�]�F�%�6����7�{���T�՘���_r)4��M!�ߞ�I�*��+q"d���?ȍ8�䕉���HO�Z��]��!�T�k�oh����c�l]�	N�����J��`��b�	�״�p,G�osc4�7�ָ�{A���J�ٵ��:*aD�;�L���@�*V1u����Ӟ�q���V_�%�@�DjOʨP=��ﺹTH&oB���|�A����s��WنG��^+�yu8)�gr�oD`��u&�~-��AU�BM�mMJiy_JCy���3����z�:�������J��(�� ���iw2m�z˔K@�8�!xâ""�ٮ����A��oj�Ȋ@9kZ��:������ߜS�<_k�G�cժVxKs $����k����{?��\��?�2��ea}�-��1/�V�N�8��XDʊQ�8J"Y�v�t��J��D.��R�_{'[.�h�� �@��,9��8�ߠ���>�n�,��F�7��UJ��R��ޥs�����u�W��$At��'�Yԩ��+��O�Ң��ɛv=Zz�~6+~y��B|�c���H΍p�j���q|�3�'{�̖���Hv�V��oH���z"� ���g������xX59H5��q!QsÄO`�%�6�F#���B�3�>*g��,�O�*��`�O�
��!��*(97>��!�=7^U�\���3�e��w�J_�����w�>��z#<�����)��R�i���`�P����88Ӿ5��z����50�BX�A=�J]��ʈ=�;W��q��ĳ��il������T�z�	��������&��� h��2R��^���)�HH�y��p��du��mQQ1PՃ"�F1�yD�ȏ;�� s;�Rd�`#�_v���J��J3��^������'���1���zᘾ����^p�_Sy�2u<nGntw�ۃJ�A�_�����L@�Ts{��1�����ק�������q2�os��Sn<xԽ}��\���"�/!f3cb�Y0N�}d�[�A�5�J������i�%�q�Ι�V`u���RvJVx�,p/�H��IG�b_q-۰������,̥z�TEP#���.�n��t������N�X�A�i�z� m`��b|+FA�VJtܯ��(�Va�8�c�/�|ѽ ����X��l\�۶m�
�O�Dl�	���}�pQ;<��gZnI���Ċ���F�E�l����g����"����_��D��79~��y�T�ױ-�<qAm��Jy�7�Jr����ub𿙡��Z���pl��!���K�˃��u�&ڷ�7|����W:A\�1��/�V�	UL�P��u����8j���Q&?�������9F��#+g	[� {R�XA�.�p��-*���Ѹn�uH'�x
e�?����~ކ�����SϚ�&##3�=Y�t����;�C�Jm����{(
W�rŶb.���`�a�����_߅ʰ���V����M�����Bn�^�~�AJ��-}}l2g�w�#�yk�e}3DMtR�'RX�(Q�S��>O/�*�(6�rC��F|DP�%b����@n����������d�)��K!��)Ͱ!����\�W�)H䝼{:�8RDK�d�E��3���|t�Ө}�i�d���`�m'����i=i��@��D�'nY�@BҞ���+�{��o���𳸻kO`���q����_zMW_2�G��8�����o�H����3o�ix�����s�B����5ٟ?��m	�j7!��2A���H��	B댇�?�/>,�\v��@�������*�5\�	��Pq�fE�.���P����q�2��p
���6(Z��"��9p����DZ)��[4<�pE��r��}cHӸ��a��wf-Xs<���k�q�I�TD2<<4=|��P=��h,=@�Љ���Ρx]�5.̫�UTS�݁����\Y\�}��V��u]x�]G�v�����!^)��tK޺�^|���x��K�H�����/�V����H�;]GD ������u�Q�� ��X�n��?��sk�tƭ��^��y4Em���r"���{f�d��=U��u���l����hk3�*gC�~?���r�f�ɺ�1�i�a1@���Q��G�z����غ��0���ƽ�~������*���=�z�Go*Ko��Oa�c˽�d�}D�]ڪ��oy9o�.���_��C�P}�JM t���a�?H�����ф�.8����U��U@��ڬ�P�>���(��q���z@-b�"J����!-���Ԋz�'}�O�rhB^�+M�n��T��C�@ �kE�����f�s>Qc���0Ɩ�InP�_���Sz���h���0��aaJw�?-:�te*�qʫ)�P�0Tx�%�P.�d��j"U+Is2����+�TV>Z�t��2RJ��z�j�y���b��
���pb`7�?����������Y�i+��>CȦdXڡy孋"���*7�qe/�osT����ũP�<y�3���w�C�$,	J��
>��r֏�0�}g�Ұ���K����]]'t5w�� be���B����u�3f�]BAo\��!�I���K�c��F�-b
Q�|#���)}�v]&9��Ɲ����
A�q+y� p����
������Vե�j$Ө��"�`���&&dO?�a�|ߜ���ݿ2���Y���9"~�W̊P��h�}�W]�8���[n��=i{�1�V�\�M(x�a
!���P�C��B4�R����Ys�@H�����]&�4Z����N��Y�����e)6}ШɵCa�|Xx����ۜ+:�Ӗ���?����k���"��lOD�l�bU��M��5z��S"�J��qj��`�/�mn:�U���mEEr�>_����b��T��f�: Y���H�ʾX����LA��+*�ܛ�������x�O�ѝ�>��+�H�l[��G�����&]�;t��쟇�̱cV�[ʍ��e��즺��ݼ:������,Xn����v��	�_</_Ms-`-�� ����:��t֟��d�<&j7�b��?����(�HMj�jo�G��/�Ϡ��.4B���F}��&ga� �0�����p"Q���)�v�����˄�� �uL�m�hs {=���D�L�:I �e��4���C/GO�XY#pb�XM��,^�����"ȋQ�8�#��Ԁ��T�E�T1��.�Zȡ[�GP[�jb������U� �h�2P��t����둌�L�v�\6�s��mg0�v�����1#b �oLP�ωK����O�Z쿺y�Hc�fȐ'�|Z��h%�g�^g���r+�?'�H�}�u���z��H'q�u�p��4jX��!��Ǎ��L�Οa���	S�x��$T� �z'���;�������4y�m�	+��v��;ެ�nh����yf9�ʵ(�rc+�(r!�F&2� y�Z
����yЦ ?@;sV;^���9h'%'g����~b�eYO�������[��W&�	ᑞ� �E�us��8~��d�w��8��q�ӄ��ZrΥ��xs����:�g�Zƍl��s@���Z0%x_~#j�7��,��8%Ꮜ��Y��pב�(P���tPQ��z膡��F�AJ������n������Q������w�k,ל���]��X !ᡫ=��C��F���\�D�ϕ%QBE�����RT}�� �iJ�X�,��y�u}�4i]Ya`�P�,�.�{�<f��(C	B�?�;�.����nlIb0/����a���*�t���+:�����%���������,���ߝ���Ƥ{�v��������|}\bs�B�:��:>	I����������W��_.ǁ�o*D��A���)�龙ڛ��!"�t����G��L��k	�j�0f�Có=+�����fHMOw��?+[�L�L���D53f���7�a�m!�����p5T����y~a��!�-�3�5�7V:ѝ�����nk~���B۩����6��]���K��"2�t#MN�."�(�\o���;�q�w`��mn�%"�g���ӹ�~�ӎ�ڗ��H~���7t���m�^z���$;=�Ec�?m�Pt�6�?a��&��a��'�D0�ň�2�ql��
>� 
�H@��[������\�K���f���b?��D�y��h~�l���	���H�?�p�*�,�yJuto��D�V�.�}�P$y��
m���gz�.PQQyC ��T��(�Ro�Z���f�z��r$�!)]c;����E��Z$eڭ��t�~a�����l��u{�Z�~�Q��}>a�@��=��{�bZ��F?U��&�S�`WaB�d6a��phB\�<����^��9�ܝ���Q�~H��ڌ���#V>Ca@@@��z!��������>��>LݯȐ��.������R�:M�܈����ʫ��C�o@H��W!��d�1nC�al�X���pW�KgH{vM|a$�$�>s�&���ܶ�K���Y���h'�t�� �{"��a���-a�F2Hr;~>�z���%��;ѩ�B�����<f�!�`�h*)N�}i���E_s�ׇ���]E Dnv̳�)�%Ox��}6���0�!���B���w9��I���3�2е^oq[�����Ct��p��k�4� �H%@	Xu���>#S&����ȹYSȞ��$��1!]��^��,/ZH�Odq��=���6�5-�dGq�qQ֦ڶ�.�fڱv�����|�:- 9��/'��yYo�#�\s���| �R\��A5������ǃ�e���	O.�k4�2����{>tPWM:���-�UsſB[����;�����MF*^��7$�������]�?�c�4ZRa�D�q�F�d?W43�FQD�����Nw�[IU�*�-��C�W�d���l>;��B..����)��3��ϓ~�o��h {>?���4e���ԅ)iՏz͂��������˂(�Ӗ�ǝ�h.��!����l����iQ�+Ur��h o��2/)��y�$�s����DU�o�yP�u��(���{�J%,��s=�g�'o���*���bX�ޟ|+���^�B����
)��I�z4k�L�r
]D�����CE�)�Ib�`�6��<1��'r�~�DY��V/�.R��n�ѝ�Lަ6~�c�,W}<��@x�bF���b�۠Z������Ao`�z#��;��=�FV�?�5ol��g���'ZJz�ԅ�`�5�uP��w9rA���QU�f�S[	Ms�N� d�,��Wa�d�S��?�S�j�����>|��H�6���%��#����̚����(ɀ=o�/m:᷌�(;�������'/�=���o��d�_B��6�ssIE�^��6z:&]BBB���}s�d��>�ؒ16�'�X�΅j-�lQ��Z�ә<a�<B�-8�p�n���Gy�q��L� gs�`v���������Q��g�?���7���8N&|�}6j�֯�����#�eI��{�K'�5��)�@�����M����D^]_C�" ���|?�u}��B"�A��'3$��z� M�lۼ/�8=Ou���)X��/�E��H�����S>����n����]�Lr�0dy�X��!��� �i��nW<U8W�q-&��x ��磖nFT��.|c�ye��bG�,t��}'�Tx�dX��J�Kssk�v�J�9CC���沥]��(��&�B������`Iһ䞒o�Ǘ����8V�+�T#=j,�aUmwΚ_���o$��i\����Yb�g̿���z�h3�A�)5��N����6�`�-�e�D\���p��6���I�B�
é�0�+�D�S%�N�b��=�i��j��ф��z/%��Y$�y��ݤ�k���9��$+����܍C�!��P���&+�w,�����*�؜�|]��wj��N�aJ�`��ط{a;�{��C]P���H��p�"�O�m?���BI�L�;0�D���&���(�A�T�KE����xO=j��ꛐ𘕥��0���՟�K�$�)T����~81y���$�m�s�}�hӇfVju��z��Q�F��S��x���2J.��ղG��'9�c����������a�Tl^5 ش����5
o����el��^۶	r�>}?H�A����@�RΡD���^<�@�Eˢ�~��x��\��|�~�_���#�tw�=�����y�	ZP<�W��?������ d�EFi�Y�؛�c�;� �h?�Zz����)�ŷ@S��y:3"̄�5�Z�[gAOL�yJ��xt�7�}��2�f�Xe�Ȫ�<���2y��7�D��Lfh�2��Y����N���(W�':*�ǐ7��Lܷ{C��	�M/���~?��>1��'^�
W�Ĵ1I�r��")n�Q"��n20N��匿�%��x���\���D;[�9ӈQ�0=���Q��)V��=�4'�$p�TW�K�j#٨����|��;t��=�~� �G�;
-f$�Ԗ���=*F��)V��\���"*rOT㽵���Ʒ�J��H��:/{��3C5��'P����x�'�G
��&�GW��f�Y�k�n�s�+��54��w⽯wk�m�n%�T'�]��>�him�;<ߝy?�u������%�rٸX2�ɿ��Ӳ�%xO�vߨ�V�V�����3�o�4s�������	���T�Vy�k[^5G�2�O�r.e�>t�7�~��S�S�����J���g\U���ۜ��4�^ȅ�6�#|x���TR��Ǣ����g�W�յ�c����O���re�����z� ��D��o<��P(0�a�ml�ޘMy�<�TW� ���7@��p�V��{���J���;u����ؑA'�������i�$�o�:' pS���<��SZ�=�-䮏�c���2)�F]���(��������G����<�@^p��|��������9�ؗi�p�U�=��	uC��ly��HV�-��1�RC0�V�Ş����/UΪaL�埪�lȶ�^Q̹nCbj��/l,t�$
�K����������v��!ae�=���w�������/o]����}�܎HD���Ftq�#%l4My�_LO��B�DbG��b+G'��U�Y��C��V�y'S2�gyyY��r�D�Ǔ-�Q��9����$.A$�Ax��̣��;K	�JҮ7�U�#A4�ur��TQ�7�n�\�*���O�h��]��f෵��hJ�t����g�V���17�Q����|�56����6�4��t��$e�t�V��,d?�HF���v��y��F@� ��.��'��s�G�gO�1��\�����q^��A1�o��kV��1M6�k�h�}O�k��^Q��o��i�<V�X��7]���)@J��遬y��l�b��;)g����D��z\{X�'��Bi{:0�-�+=(u�\E��t��#�炂¶m�_�-�����p�_=b~p9w�"�jzi�A�+��9����o�o���p�*/Y�,\�=��`Sg?�?m�p�Ć�֍1��t� w�����"����L>�P$]`r��y�P[��ۋ��}&���*B�s���~
�Uːy��{�z�K/�.KUj��1i{0��U ߂��� �8'�)H,6��C�nl�J�v��=��p�:��n�3h�w�j���� i�vH���3Y���0���ď �?��d��EW'�8à�[��M.�^NT��[�ǩWOaf��C����Z�ӵ�$��X`W�a�h4"&i�S�#"�Yg��=�����K�$ap'\���o@�^Ks��缸v��<B�&�z"z;Y�����v94n��)z�6m����=}��/���^�VR�#�f�BN$X�1�h��_�/f���zH�c�����V�"�=K���*)@Ib11
��ɾjnxD�ݪ���J��F�Ks����-�4��IE�^�S��������%A���������Yf~_�,�N���V�L<[&t�sv���#�)Lg����:�N�)�N8��>��<�������Oȸ�U��	�����k�s{h�T�V����x��l5����D� �h���|�ӰxI��@2��	J0�[+�0��+�Ņ����t��pI��g�޶��$�)�S|C�Oaڵ�8r��5T�]�(O�1��8�
=�(`�A"�f��R�ޟq���r���F�ti#���"�VI���"A�ѽ�m2��6��䤋�H��:$�{{&X�S�)�
E��0���Q��7�ѣ�(�����7��.�v8�!�"�;��L�?��y���{0�W>�m\+�]*:������m��㤐���PPT�n��_n��#4ט�ۆ���(��u_��a'
���/���x��ZF�%�9m��[O��_�~)}�|[�9﬜��.p��)�ߔ J|�D���d/�Я��y�Э����9�pm����#i����s�%�Ǔ)e�;�3;Ƚ~N�U7���n=|��s�mƧv}Jd��1P�lkP��\hϼ��@�����eج]c4�0?��{�*(Q�2M��zx����=���u��6����=JX�2d��r��4��E��QP@��ӆ��)99]&�666.r�$�4�g�*++9�iQ�C�8-�}��?<=a��i׌��!]<$0��K �/N�Ft��m�%�K��u��d�l@�
�+��ŗw�9����jM���݇���+�mc���e��λ�I#v	X��ۥ��h�b$Ah���v5x�3�Z�wB,��*!
�b-?�ό���L�DQy�]$�5�F����~^�O`
��Xsse4�m�:�{?�/��m�ҍ�?ɩ.���xB^�pFΗy�����͜"�׆��F�8�gX��) �R��=�S���f��1|-�b�Y���,y^Zʏ}�����
�1��T����9q���^F�Kɀ����p͏�3k�f��pSC��?�*�8�H�x���Kr4t%H�q2�B)X�9�E}>��f\��˵�N�
�Q��ܙ����M`���M���9]���E>� ��Ų�-�c���{���B�~`A���(Q	}_^[��xe�Pq��V}.���).��$�RRQ}���@��yz��|��D.��/,�d�~� <�Zް]�xL9����qnKw�u}�n����ſZ��#�sMF��N�<�l��_÷�4��PЏp0��-�/Ɣ��G�〘u҅��/h����/͞�h����;	 ������rȯ_��k���R^>(XX��A���Ϙ=�g���q1V
����
�v��P�ɫש������c:A�\<�e{�3ֹ�;q`�Yr����*hmq��tM����1��$��k�������H�L�V������2�_�k��1�Ii��nVD"֑0"XN�OO�?yJ��1Q*�`~y0�/���\��g���e��ֵa:�C�Z���G�W��yl���`��7������Rc�X�1����j*b�gusN+�.�yC����@ϒY�6�c{`*,�h�����{ǲ��ΕV���E����A���{}�O��,͛o� 93tWP�0��[���.	��Ԓ���ئ�ּ?	w&���2I��l
�H��u�i��0����$��-c�_�yS1˶-��9�.�后x�X7u�űqcWEaW  3��yP%�k��?��X:b!	��q�3�5'�ȒA����]n�{���T\\_�\=R�����)~����?r�E_N���;��%�aF���^���+��F���lx	%%,<���0�=���N�!`�D��zmYSֆ�LhXte�&{<l�n�]�	)��M�|������tp�(�D��AN*����^�X��Tv����#�돜��w$�9!a��DCq�P35I��I���1唔>���`R|��jQ�!���ї��hZmmm7?U���P���/q�Z�yW@�h�W�2xU(�Q�K�E�Ӱ��{t׶��ʋ�m��ä́�JЪ4`�4��:љצ�����I�WO��nh2F�3��}�
 �7�B�L�k��1Ԏ
)\nI��uu
�����_M����[ɨ��N�l6�y��"������� �]�Ӓ4���zr�c:�r�#_bY���%*��������(
ȕ,�����װ��,E��fff0]�����*�q_k0��0Fy#�B���|t�m�\�H\��~��#تq��+u���ױ���t�SE�^������iA��cd�ۑ-
�kjR���[���^x�aڎ��U,a��("¡��{����kw�@%ɑ�:)�B]�'���)^8���:��q�h5M%X�	`cc[n�#T��G�о+���3 K��Pg����ίL�fⳋ�F�OL6�[@�'�KQ�s�U�ڳa��$�NHR>�(����U����L�Fv�5k��05 u�qaHX�LL(�����,�J�
e���l���}�3�V�>�S"ވƨ���|�c+0n��K��j��q4���/)����k��qiX�;�5Q2�6aC��z��f�����Y{L�Ͽ]� �*��Bj��f�P�Ï�k���a���@{z��WL'������(��N��;4 ��g�p������s3^��Nv�<16��H�e��]�ɢb-�̈��S�/An��\�5/'����y�m�H�	�����N-���jis�mV.�"M;޶��}�%D�{��zy�w��P}��X6���G`��"�m��n�\#x���=!ݼ�|�.1eM?��f���*å%��B��m����7za�8m��+�G���[��K��9+�H�st�ʋ����(�c���$���fa��}C�^ԛ�kة,�긋����7����{���K|D�
���QG?O�q��m���s n��ڶA7��-�%ln�N%Cb�u��aPf����zv�]�����w�:��B--�p�����"�:��J��0�_nҵZ�pY'�mi�����5�������+MjzZ��DHB)�cJjjРU/����d���r�8���������x��A{s98L�WpF��?�h�[2��#=�����ě`�� J��(�?���aPP��M�H��2`���;�c��}��'	�R@~�]gF?O9$��]��S���g��R�	�-����;��(�!(�H���#��D_g����)���0��n��
 ޴�:p}#��;�1�Vk�*����<�y%�`E%6��������!��I�
�<3��U=+�j^/K�z'w��*$w�x�6�L����=�3,<Js��r�k`<vD�I����@�����L(�� ��+��\�ތ���	8�F��̈w��_Oj:����\dC�"�}�.�?�u�s�G�G��siX�h��_!�F���C�e�,��UiG\�C��������?s��^��ގ���3��{�j3��'���G� ��${��L�i|&AK�l�����&�����~�nUs��^c�T�ק[h����΀T�7��'5C�j/Ѐ��9Y\afc�C?�Zh�C3�w�-�E�ui&_�Q�13(`��c�K��"
Z�"�9�bsn�U��w�UZ=j��R1���X���';y}���φ"�]�:}� �B�����0�vtd�{����Ã��WXX���Z
n
zԘ��Ԭ���f'E�S��L�CC���]�%��9����@�'�B&r�F:�����6���a�_I� �i�"�M��Ő*��+�����Y�ŃM��Wq{���Ƒ�8"A���}�Ʋ�ޮM���'�����2�J��4�XE�9*��d�mA�O���X�n��F���V��Ixy������t����c.��*ͳ%�C��\u)�!�FC~��D�>#�3FaQ��Z\�\��Ͽ\������-�$Y�PS�}�x��X\�mo绹�1��ԥ��ę:���!�g?/uy�	�e�2n�R�d�D�;�s��r#��Jhb��r�t���,�3}l�=��F�������	z~�	�qgZ�0m�jkX�����"�G�cA�7�P#�b���5�?cZ�`�1 �ݾ�N6��0?�i�z��%�<b��\�l����7f@�Wg=ƥ��� �a��ywz����|���z!Vr�Ӆ&�B,�]%==k[�����	��F�Ñ���

��&B �j�g�W�;c�H��;;�����䘥C����:���j��FI�Ā��/]��HKD��$H�*�>�]�L�>��z
�e�k��!3�gץkȗ��Xi�S�}�Ԙ�9<!?����_W� ��*(*Jik,��a������'N� �	EM��$���0��C��fz{�O�Ve���Esy9��ˡT��O��:�T��"���-�uH��9����Vw �$�9���
��2תľ�
�TD����~���,��ЛG�le�E���t������H���й�g��AB��/.�D8ȡշ@�4޲�w�c�x@�d��з|$��Ga���¾�΁��쓟����
>w��ǧ��\�����L��	��Ż�/S-�1^s$Ȅ����P��cy��%�����<ۥ���C<��?`�bP�6��5�UAqQ�Dm�q�&a�^^ݱSܪ��~J��7"�]V�;�����_���|����?2��J1�B�A�yK�P� �#x40p�hW<���k�э��T!�fI���vՖ�x6�e6�ނ��im�	�wj/�L�4x�9o�3���:�Q��%�e�;E�9��4��C �>�xC�k`���AIh�($ s?@��>�>erh�F��X��6#���n���EzL9����B0��OO�+.Hd0TIM�\��Ȗ�h���!ľY���*a��9x/ �u�����>{���WV+�>7Q�Y��dN!_�Bf;|.��}s�̃�#q��ֈ�:��m��i	-�����V��ф�v8�%9!""6ZϒC�o���XI��{Gs�DE6��Q rGO$������R������5Y~ǉ��ݗ�`k;���|��i�c��_����\#�Ϡ�UƷ�pE��Y[�\����p�W��'�y�۫�ܸbd����8��#���OR��'�H:0�ĝ�> �v8�ȟ|��� MKԘz*��N6=��s��h���͐w���#��u���$A��#t���/�w������C�����&�P7Nt���������ސ]�'XxC�~-'��ɳk�e����������Ãt�� cd@��Ei8IRs��m�����>���XjmߛI[�Z��3�r���(�?���f�O`n���S��*<R7�S _�"����_n��PB���*K	֬�� /B�޿�ZBB��J�豜E~�an�=��V*����'�d��u꒩�*��J���L�u��
��z���G��^����q�q��s�ؖ���ϱ��b����9��G֯Y�ML��>�(%� ��|No/lQ�C��m$R��t����>�;$��X�o���>�H	|���ݪ�
�S�&�����KX?��T�P�~b���(�G� k*�Z�İ�Z
qX_�,��h�^~�|d���G�!�S��E�5Bq�@va��ĐJH��So���׷����XZ5�;��,"�"WTT�&��{}�SRS� 񬩭��tf�?˕���@3���^����� k8��>���4J �!<�q!"�q_x{��K��B�Κ�|@�o����I�=�O��N5Q���2ܣw,��M�s7a5=�p�_�f���7��ɂK?�H�d�'+�ٜ�n%Ƃ��t	me��%�2�ЗZ?@B"�%���+�u@q�@[7�,�9�d����k`�E�R]hi�Bl���և���N]�ύ"�}!÷���Vx�Os���$��3$/S��EL�����
����W=1`n����w�dG���s�F م_ƭ�}ղ��w;�ܷ3��=E--��O�p��msڠ�}�����}���'gpS!��J>�;@lu�p7�=l�rn4��U2癌�?���͞"�ɛS�Z��!����ED!�o��������Kޙ�>�߿@Ro t��+ݙ�DQ��z-�:����^��uum��ᆻ<>=��2���>����RQ�;������#!�6��E�
�ۆ�[ժL������Y�"����r��N)�2V.P�l��Ig�U�G���r�`����_��5�͉アdn"�5���d��K�}X#i�ˇ)�|�$@E	luFՖ}ޮc��A+�/�$������䢱P��Z+Y!�3=A������8B8$,�p�2��x� e��ӕ��/��*y����p�����]+� B�W�0��p7�[�H��Y z�@��=��ca��=|:ĭ�$qD[���2?;F�� ?�2�2��r�xK�$Ǔֱ�	p6ڋ  ��k��"�߳��w³O�&��.ka��P������LNC&�}����a���i�F�Q?76^��w��>m�3�W�ϐT0��@�?����D�� _K?�8I�&�6T�,�N��hk���uS���*�7�ڧ���w��g���\H�Sص���~7e<��rys�y+�$ɩ�f!����U�;$W�}�偀h�V������&Ȥ 18����-(�<���N��1oA�fy �u�y��x��`��m
���/�i�U�R$Iz�fM\>"	_�������k��� ]PĢx�$t������D7U64`�݃G�,��� 6� 	I��������f���*�*�P ��:t� T�UV2�	��C${��?��,� �9����؄
½u���OW�ZE��C���~���s.-s.)�v��.�?�)��k�<	���
	ݺ2Q��>�P�w2�m%����pL�t��m8��dB}���^״��)�0^�>���_n�QYe?$c�s^�vt��%���G5An4ZzzI�w���_>���	w8n͗�~��Ub6��HLOǇ�l�h�������+F)���J��U^���G3��$�ݳJE����GH0�sz4
�ԃg�i�۶Eiot�0�,`�K���e2���y���a�,�D�K<�Ν��l_�GN��`Q���X�[�w-�i�|�~ī~M{j*�iCD�Fܽu�G�60�Tv������SGXN�/��t�����m��b��"2�9�EM�����,��r,��O�.R��5jo�e}���Fw+�޾U}_\���DM����ߜ$U�M��,�Lu[g���ౠ��eR ����K��?�H���R9A����.�ttI��apI�ԧ�\��0��f�J��փ3.�Ȑe୎ͣ��B�Z$��P�J?Q�W;�&��L�P�e}��\?����������9�	C���������@*�
8�G��<�Y����}i^k؅���/�����D#�hz�8�@NqW�Gˡ��8$
�.~qzNa5��̉�&ǽ�s��d�

><'���@���M�ی�;���s�f������
:�Q��H<j?Zu����-P�u�rϱ�#���8��Ϳ(9�����;N8�!��A$�L���6�~��7:�IHD�C�4LLL�G@ff��	t*JJ@LLLtRE;����ښ�Å�£YA8���ca�[�d�C���c������(����B��|,�*ǥ�AxH�m�Z�b�թ�|����Za���n4uB��}X�N��<At!A�_�0��ķ���-�O���9�U&.�V�d������ߝI�u��L�om�9��X�j0�Z���y�#�6��O���p���<���i�`��肵�.��ty���s+\�� ��Hћ`�� ��|1��	�]��䨅�I�B��볩b���Xh�D��.�f��:N�j�8����p����q���m6xZ��Iu=;����:���K����!��3R0��w�w0�1-
x�W�D 6�#�u�v�/?���^�����^�B�tKd��[[�s�G�^��|47/�������q�ڗ?��!$#K�o$�����	��1��f�kӀ��`CUF�����߭� �aΥ�E_}m�n���#��J<�A2 ��s�c�SC������P$kπom^��ڶ�'���Wƌr��<F3"BdȮ�2�n>�o�}e�!���ym�$�M����w�&��88d�p�eee-���SC�4��\���[�ŋ�Lw�"��� �;�n��M$��e(ԮAȦ�I�ʷ&!t�v �[�=W�;����fr��!U�SFyI��c�����F�*�3>s#~�v6���oj��冷]�)|½�>\�vy.�{Qhp!G���.N��]���0���v�^L�����`�/![�x��y�1%������=���q�'�p�x��'n���� 2"_36m�b�6a/�Ԫ��z1�irʖ�i[^ܲ#������� �I�ٹKEq� �̐����_XS�w��-7:�mf`y^KD��eW:%D��M����Ws ��Nk�T���	�]A�1��4��`)�?}��&���f�oP!���m��/�Dluuu�i�%4��B��~���E�����	�{�Fbp��XW���dX	h��!���E1����/��"r����fZ^%&�eC�.��M�����z|'_$����{p�Ė���n��D,7����hܹ���;�X�iW�ƀ-��3�C�撳�;p�?k�q�^���D6Kf�����O�z5�V2�C���jq��a Q���� Ձ��	���MN��v۷��XS�}R��R74d����]�E)O�~��6���� quulL2����ٰ��K����1N-Z0�;��4���t��u� J��8�&z�� !����i?/��X�F|=�G@iw�w�mN-͸�b}��&����<o�t��ā\���*���J;�;�@ؓf�]��'`z>k�2꒱�et�Є������ �9<�M�ˇa^��xs���g[��-�wC_��:�>i�%N;�}���xJm1�'��>����� ��Y��S���U|��N<�\�_ rÞ��.��o�ǳ�NAh #x�����Uq��S�r��f�����$D5r���Z`�M��Y"c+�a.E�T�F�;,z���o{���ϟaaHX�G�%���T��Fhy`dd{У��8���8��0�����c������q�����Vҕ���!�{C��5�y����lU�6��?�7Q��l��.�d��\���� ��*�Wg�%���_ )z�#�k�Z�H �Z	�=Q���^
���/����<��,����}I	^��^hΕ@C�j���[Ξ�:(�Ë���=y�E��;w����!����Y�r����_����{CWףizdl,*�o���m��p�G>EC���F?[ʓ��SA�I�׹L``�87����\��""9	��υ��U�W���hRy�|�jV��t�Y�|���-r%�CbE�|�3&T�&]��W�~
BD����޴_��r^`E�JF4"Y#7R�xO=�*^~X�_d3l;�4}e	9���1I�ڿ���������n95�t��fKP&Fx�'N��F������kP��tg�NؖS�X(��oo\�k<�u��~����ӹK����E�b�n� ȝ!%�'J�E,B���١�\��;�QM4i��wm�}-J��"�s{��?A��&�{��,ض�)(HB�"����>JK�,�iT}������Q32J@#|O�Ą���gF$,,<U F��������׫�+h����"5�B${SE7
��g��|�Z��M��|f�U�-���BΞ���'\:��i��A�Q�eH��� �����t���>1��0d�+��)�m>ȱp��_��бˍ}"�A���f"A%	hN�h�	#�v��	���*�(��O��� �y��DhJ��/�����d�ڴ���k�㱱a���:�����A?^!����E������� �Ty|lc%�_�����+L���mΓ��"�~�@}�E F4��i���L�����B�M�U�Ga㙇��&�"��p�NjF�`�7��*;k��e����e}z}(�F1V��p��`���]��K���`����Tf�;*��3n�X)���z�;�Y�����oV�P�U���Ƌ/�E��E���큒�Azx�l�)>�&'�	� ie�M������}�s�:�b,r�QS�6;,������]��?�J��b�
��`�������#�>Ά4�&�k ����8g��x��˨��f�u7)̡[�����P�uz��u�����
��Z��(l�8dx@WW���tDC�v�nHx8�-N���k<����槪T�����u��T__�ZI~�2�Ù���8N�1�9%�_��VQ���S76~?Ǌ����q��>-$�7�u��y�a%��ky��m�`����}����I����M�&~��fd����]o&��օ.��k��;���yV�w��ε2�s�J�y�rk�Cy\��@z�B�ȝ�{���&�z�o'K�@8�Pa��҇�������wh'�c������c>B��������#���J�ˋ;t�l�͛A�+-��>1!������܌c=��$5�"��l��_�PD����A��o�����/�����6U�DB���� ����f�}�es ] �K	$�ih�w���� /i�}�o|ݹ��^�h�QOֻW���2��}�L���n�!�?A��'3�C��J�~I	!֏���{�mm��*�c�U5��g���~r���aIkVi�+�qM�,����K?�]j0߮O�0��7�F��@$=.�Ý~�4�	U�i��E��y���O"oy,�bx�!=�h��G��=A޸�֌��P�L@t���@�ʽ��χ�N�p�fЂ�/�/��q$����j_4^x���a>�H�O���d���ejjXlll�?u5�`&�B�����}0���3������z���r�O��s�)�{�����O�`E����o��K���=�~{��}�#�Od��(5�KF�ާ�g�2x�E�Zy���YM\w�Ҷ�+��E��g�|u	�a&�6����806�]�_倠<և����lL�;9E�AMg�_u;*+F��4�i�^M��W,�Z䡔�VP7�|w&��K����F�G�O��R\R�MF���_`iY��B�b���ӓ�m����������0�RR�
��ggҶ��3��p�
t���d�)�a�� �	D9R�YQ�6J�!���@��D��J��׆}�=���/��OK ����#qk���l��o� ��_g�}�%�W�����Bv�"L\`����TS	?�� ;�Ѕ��o�{�g�Ѓa+�}�y���F�{5�~!�_�ij�,����Ib��=S6p�$���B{\�ftgN��lX#6J�y5��-%��p\�X�4Z��-/60NfSȈ��b��`�� �9����Hgs��ȕ���*Y+�x-Ņ�T=���ڎ3�j�۶0�g��3$�G	�t�[��Pb���g��m���QN5y����Srrb_^^&+xԴMp��7}<TVV��$|}������E9��tu)���!�zI�ʨd����A%�@��������#�>�jhY<�b��\�����N��-i��䓟�4����`"gy���j\�PI�u+���Nj����j�g�O�<�����u4�Q͎�*?��	'��q��5�L3�6^����F�/�����O�4C[<*�O�P���8%{훜�I�oB��$�=�Y��C�
5� /S;���o�z���n����qqR�����0*w�=����B�3g���!9����z�����_������EV�tn9��kƊ\���I*��c�p$��C��F#�)����w�T:UY����z���k�on�Hj�7	�{.��+��ܠ���D���)MNB=U.����.}L���.������ag_�Z�Hͅ���D d��W�ٗ5��E���d;6���5�'��t�������_ob����u����G���s�7�`�b��5H�-Yk=�#� ��a;IB��0�mZ�藧X��B@1N/�zǻӡF��
o�>����"��մq*����\�9�ow��#��l�,J�� lPة�D�.4��'��g>@c?���,��-�;����t�	�"�{wwZ?}x8
$�a%�6��A�/� JZZv&������!�v@�ã�P깽���Z�AYr&J�=)�M�c��$��Щ��TZ\�qo�����G�"�~>�-\������<�e�H�q6l�8s���#߶�4J�^�\���ٿ����Y�T{��*G��-*8�*Xq�Wb��mp18�����3��^����+���h���Cq)ZܽP�Xqwww���Ŋ{p����P �����{�e��a&�I��g���9�9�¾�$��K���Su�i�9��mw�><Z����wcNO����,��!�����9lư`!��u��i�ւ~|VT��LD$��9+�z:lĐ�P
��TVV�nh��.���-�l�W:F�5���Z?'uk�|5��~"(3�_D���hi�©W���ĢND��.	&�WI`u4crj�x�]o�v@/¸)��!+
��ny
-?����5��ó����}v�T��T�fGƒF�4��nW�����X�l4�֯�A��QѼ��;�m��ɦ���T�5��=z2ª�aX�Σ�`Y{l�½4	37�EՐ��w؞�?�K=����p� �j�y� ��������Y��B��[
yjV}l	Y��������h3�*�B	���L�i[ר���s�#;]w�FE��3!2Q�#��WM�����ڏ����h
�<�X�
�����6F�Ʈ�QW�X���EDD �����ӻ_z������BYKU����
���%��������%tL~����k)#5�B]&lk68��̖g'����D�9���V�#��.�N��fzckq���r�~��oA[$D	�/�Օ��ukP���������!�	B?�g,�0�R Yb��{�z@���q�"Hf��f#+�+[H�B�s|���q��������\c �t��;���3������~���E�e�,�LI�kkk{7o%sV��1$!RSSo�i�DL������Hzx�|���w `�@~��D�;�"��0��_S�I�Ss�d���0��)�ǂ�QZZ����f�������M`k��y1��il4�T��}g�Va����J�-*�G��h|��+Grp��������퍹�f��tPH���1��֧�I��ͅQL�g+����c�"�����G��E���U���/��6�@ay���;��Ȱ���7���K�q��-vn�5�4t�#��$�V���j�@��s6+���V[}�2��ƣy��́�|Jf\|e�]��n�n�Х�w�ۢNѰ�c�q�96�-�C�4y$�Z�g�[�]ȘJ�\.��/�Tk��O���?����nwoo��������]�{^�r���9����sZW���w��� ��?CC0��d <�.�H�{"2C��o߀��;�Z����Sn����*�]c/'.ܗf����K�#��Z��4H6��t�zQF�.4�ާ�s"~�X�-�����Kla&���[�� ���}+*^��ʘ���9��L0��ծIZb�L\��fz���@�{ܞ����do�Ϣ���q���7����=�W�"~KYPD�֎I`���a89�����}������D���п�AJ�
 +� ����))�QQ���B�`����������R�l�#~;	���z?>x,G�hO���F��V)��	��M �ۂ��`w뙼���f���ˉ�\��x�ݜ_�]�he���B/+g�фW��>�$�4�vW@����9�5�r��_i��G�w�R�A����[�;�8*��c?�+:�k@'L�?;@�}K�Lca98�75�-��X�Y��4�&����G?{�5
1�Xq���ޭ��ϋ��VՐ���e5'LR�QXB^�lz~g�-O�_��
[1�~c�<��Q jA+��*�����s|lE�|&\�K@��#�Z�0o̍<�[����k�l���L�Q&5"�D�z>t"b����5ڪ��Aw�A�/��|����4�8�9Ò���lF�ipe������Ko	?:���X�-�Y�\_\��)ii��i���@GO1�hZ O��=1������&maA�S�w�������6ؘ�w#�V%�5l��)��N��Y�v� y��DE��}�Hf�I[�ӕ�y<]2�1kÒ��"�_(��"����B�n@P)�9ա�mm������X�y����Z�ryf��l������iy�{ԅ1������6C.�Q�ަ�Qfk1ӝ?9��3��:>臆~;͋�ߡ݃�#0��@�rnM��"��ظL�`��:�g�E[K�33���# Ԙ�HO/��'����=''~\�e%�����D�u�'�W��@��6��α`�t�\����S�}n��de�~w݄�."�P&���VT��/���ܳSa����Ք^!O�|�e�v!X���͂�'�`%65���!�s�rt/kMч�N�������bP{�-���=��S�s���y?W�29U@�j��{YSғ�axDsd��8*�m�;7!-�lhP�3�������{�T8�kC?J<�i-�,��,B��{@ś;nV�@`]#���~M\���@����g���1�E��t�K�$Ⱥ�u{�+m����t0�j�#l�_�UQ3�w�ܨ�:���}�j�_��8� �%j��+uA�҂��z:pyE �(===���>tCj;�w����蟉	i77�啛��Á�Q�����<�j@��70ݿ�_��!(�������r�~�9��Qs>����o��V��=.}e�����|ʸ�~����l"J��K����Ra��D,�dZ�M�[�d�ɯA��w���ĝ����}��+��_Qo��KQ�̤?���X�[ ߜ��_�;|�k�k��U�Ir�»ԑ^��}�]�a���x������{W��|b��h�F�$ad/8��x�
nб��o1GG6YYY%���m��sC�������+��06��s\*X<l��+pJ���ޒ���vӣ�hP����g�9$,��κ��6�p��^'����y#HD����ݍQ3!Wԙ{�o���)����"?��o��-�-޳R������U�e������z>uMiE���C�?m�w
�6���(z�w�9i������w-@df��1���.�q��П��c`AZ�� �`����&ŝ*���{�	�����,z�A���axk&�l������c�$>d��[�lBm��.F1�n����@�/�:��m���^�S����m��L�v�f�wX���w��ac��]������>��N����2�@Pj����2����"��FnF�d��B���! ���p�����a���֔0(7���(������������$�	�-��y*�	��q��	���IF�6�$�ϣ�nf��'�+��_Gg^��f{R�_[��@u�w%p3�v&y��iS�3F��m����3鬖��>�{7��R��KE�c�X(~b��K�ѣ���
�3����68)�|�ٙLNG�mDX���*��@�'�u��`����_�yA�2k+�(�)������������,�{�_*�A�����`B?d��9������N=}�x�i���gnm-���ZIee�Y�������������PU����,䖎x0��/���ƒH�U5���ɫ����:��t���/Tm|�H������A�6�C�	q��w첛�鸐$"�z˚rq���f��;YnGpd�aK	�:��|�|��T��Tۓ4�[��|��/06g�g�x��I]�����+�̚���F��w��R�ښ���:~ϬL�.��I��h���Azȃ�y%���%�u?�!p"��&r��I���� ��G�����0�/���4��O��wё�XH�Gp�X�-�m2;4���[�k���L���`�Ps�á��ʘ�C�H�u:L7�W#7������p)�����(Z�쾡�ݬ�>���C����`�ͻ�����U�V1(g�+��r�FS��(hi!|yy����Ǆ�=Tkk$����0�6����e���GGG@�''��9�g�w�/ �����
g/́�l�8A�!l����|����ka�L����[g5���?3�:�-/��G��Єy��߿үv��j	w*�8�iC5�	�>C0'Ͽ�'?O#�GY��_�����lBj�����-� nO��NJ���8��Ofc����+��p�z�)1��1)P/��O
  W���/�=�.I6ؘ���{h���-X��.


8i�LM���)kkGH}��R���*����9W����^��Ro>>>���U�_��y���՚��İ(�疞��ٔ��%}*8����	a����#�t���R��z9��������3i8�����-*`�G�K����.��"�-7�-uٗ������f�Ami���M�R�B�msǆs�	���u��ǳB.�����TS/g�_�_15�B#zan�+\&t�����5OR�7.�e���1e���8rH����уW�_�r0��J��ф��$���C� m��Ϫ���Fs�g4���>m$.����r{��68X�r��ℰU��@���BB]��$Od����A��:��PC�I�v
m�E��qp�����v���	6U�%%t�x�KK��������;������p�2%��wVwt�Z5\��p��"��҂����������<���U���MI_�����{rrXL�'N�gۻV�vbX9?Mr��<�r��Ha���כ���=�8ιc��w=�f������࿻��<���x�,T���wn*[���[�P+�
|��`#4��D
�PRd|RR,��g�)+�t.Ϳc��]�{[s�Z��9h5.S�z�'��8��l�`��j�w򬂈�hYeĉ���Kط�u��A5���u�vY����uL�x��a��*t�C�!	��Hխ2\6\D*\	 $�@��LV��E�N��7�3[��O���OO⚗Rӟӛ9(�&�k\]�ڤ���_g_e�/����g��8(�G�V�<޼OOޟ���[<�KKK���?j�	��-��V��²~�25�����k�d����*H�ψ��:f�~���Spr”�,U���ھ%��[^���q�<��	���φi3t��˛�:l�'�	��P�6<H��V��)��h"�W���/! �4�Eez�ڟ(�!=^2&�g��i߈�?q޴;C�ߌ��X6`��?⯝�'���sti裩�O��`Ŏ��+)bo���R��,A?�\���o�M�D�?h��P���hm}���bii�Xإ[y�x��X�8G��Ug�m����)dt<�ފ�N^'���\�0��V��9�R�u2�|�:�Wӊ{�<ew35�����ÿX�tGS~�Dp��M�w�o�c'��(C�G
**�*S2�뽿�]SX���H���`AD@Н-��>��@��7C�v�;+���hU�� ��SRB�a_:/�0$����3ɞ4��kǍV��1���=��*Ԭ������EEi//���|]���P�x��`<�����خE�GE���i6�u�Q���Z��]������c�ܠ���)�������W�A׻S����QgxP�v¯/,��F��8W��^a��[���?m#Fn!f*F9��陸:x<ox�r����t6��2.n�W*��?yu�����qv�
]w"��>/��#x���D��d���ң
I�8���,��64@�NQSW7�}7��t��2��=���$�`o8�D-����޺�к�OF�r6��棟Hœ�U+g.g�҃0����.��Ѕρ.K�B)V��J�*\�@TV6�&���fɦ��TTW����jrv��
���38e�<�ډ�vf	<�m�шC
Y�F%ל>j-d���A�/l�h�sDLR~�@牦�F7�v\ׂ4�K�k�
"��F'7�؆��f1�� i^ܱ�b�����=3hы8�������k��h��_3�A�Q�酘��K���SP�i����ws�p)z{R��4�ի���*=�v/�������`} ��ۚ�rj4Ə�h�aH��%7֖��F�b�����|�x#A�k���+ݚH;$c�N*t������Z�p��Y��g���P�lvni�$M%
[���)�R��y|?)��|�OMIyO�XP:�������foo�.���+��w��P��'k|hu��A,���:|��iM�zY����o|Y�L#=�"Sr���r22�S1� �0�����=�Ė08R����O�
;��-ؖ�L�1�uR��
���ͷ���	;����g�o���G���_�6?~�}qW�K�*>4I��
����2��&|z�����cѸ����p�V脌�Ѯ�m��P)Qz�Wq3�y���u��f���t;0m�"<X�t��)2rH:sl��Z� ��郚��)��'WdRt�������S��
�]�|���&P}�:�����x�1���e�����f�w�?��֧�u�7�&���(6�+���nl��e�ph�Gufy��o.�OU�^�I���}*��)��1x�S�A�,u�6nԋ�8��(�T�_i��֠��I�)I�'���5�\Y��L�vy:iA��v�7#���r(����&�󏦏��`Wt���x�z��P(�ݹ�W6���ӂ���-98Š����ds����f
����{Š�Ϥ�b�	������Y�˸>%ac-)�b��Q�߄U#��85��p<��t�slU� ��Ĉ�#��-��ŵ���@��?��jjs&�չ���?�c��W�F�\����~���쬁��!���"�,��ͥ���]��"��ͤ���=���AՅ�B�9�i�}��v�������#��O����"C�1�ruޗq�x���d<�(=��n+'}<?^EN�>J(��+D�X�b��C�@��[Jg���o{ e`�,���&���J������p)񐡢���|����l����<��X:�3dE&�A�U��ڭG8��-5���4}��d�z3�N�=w0�}�xir�K:&JVV���I_�n+@Φ3%##���7?7���3�^P�\�WV������z��&B�RA
��s�hU38W5p�Z���"U������ݹ�qs�.=��w�H�kʴ~~�F������
е� ��PL0��Q�/B�z#�d��]*�M��(�`�ud�c	��Jd��]��g#�qŲ����V����@R�1�Z<��.#8Oj�n<�
�H V+a�o^$��;Z�2�ZnwRR�-��;����#S�Q�y�`��!9[�ln�
f1�p���t����F��K*V�3��^q��۲�Pv�٢|<�D.1htDQ�|�b�uB�77[c�ЬI,m	�L��⢢`��Cly��C,��s{�v1=�(��
���7�T��|��yߴ�l�Y�S�0�1C�~6A O_���x���?�n ؋P�@Ǭ:�XP��{9X�2�0~�gӳH�ʄe�T-�,�Æ��6��i�o�[��@Z�0W�(Z�މd:֪����IrB�o5�b�:( t��Ё����#�Lٶ00k�4�C�ti-����@Hٌ��?;){����>T�_��N�$�)�0�i�jX���utb��?��I��5
Ԓ�R>q�oim�����7�ol�on&P(�X��gB�d:N� � �i�������$ �a�:F�m��TP3lvg}.ȡ����y1!+!�)�s> ���u��Y�z�]�Ԁ 3��5�	5���F���i�|u^�l@�\!�$S���@�
פ/���.�	x~�u[}ٴC��q3lҢP��������5��O�\叚�'�I����ݷx���r��7�c�'��?�|-O���c���>n���+H�艒P�n-��!�G�p���S��_J����J$���@Kk6�W���btt���,�v=����#	<--���i�4���;g0��ĝ������4�]�����Qg��h�a���:���ET�yx�Jԡtz�ͳ�2��u �V��y�z�%�Lqi�A�T;E�	2�A}��~~����>���T`�nha/O��W�p����!���NNlL��>���)m��c���YXX���Bxv6���5���V�͓�?Q��L>��l$����L�镶�e��*��O��JK�	���2��a%��/,�!Քq��TA�Cd�#�P{o����~3�4����D?k�]0��B� 8.?�n��RD�#&`y�t3Ʋ.{��'��`���A���3����:�$���N�u�3���kW��3o�	31o����F{�Ω6RG6܀����&c$�O�'7^�au�l�.-m:���1PJ9�짹�)�?țs�|X;L�O-';{X����>��1�0᎘ĝo�*(���<|�"��I���
�����&�]G�L	ה~���e���\��<�6��I_]�p�r�C�<j�ӄ`�4�g�^����2�#\��DR��NY'k�)W��'B��Zs�$��;:�����������ۋ��%�U� �X��]�!�H/��j ���`8ܲ�$�t��Y�mi�����d���g�
�����������R!~�pq�)M�,#�r�*p�B��t��fP��ة:�.�[��J2�ĸ��~@��'x�
�y)lD`�<I&b7A9x�-��� �r�W�Z _�H���Y�6��u��/s���Y:]�__���������5�u��8�l��]��i$�u����*�j�t�Q��$Or��ȅ	���p��t����*��7����&�b �U��~?|Qt��P<�0�u0G�
Ā� &n��$�=���y�b��������ox>B및��21	��t\]#</�)e�J��V<ې:=c�V���0X�r������J8�F+C��nz�Z�H���x�"sxfS�8�)o�xm�(P��2�I(K���R��e���D��7[��س;h�S�:lQ6��A��%c��T$���_yq#�g�S߀v4��oa0�f�.�^���01����8�l$��㔵K���y���(��<�,0�%�^5�Sac>�N�i���38���yv��xޓ�?ti�<K�*�v���&zO4�-��J;�K�ݷVR�
'���t��d��V�Y��UX�}�ě�U��o[5B�^w�=\�z��6��ld��������ll?&�C�C V�f����ݬ�+��,��y�2t|J�,r��.C4�%O>B�� ����IvMD ��z��`GE�< �n�/P͗,����.��^�1dM�5R�z>;��C�\���U��Y)qn��UY0�F����*$����7$f4���G+��}
��X��c����,�gG�,�8��C��A%z�Y?�$1!X%F7t�v b1b�qb�b�ab�٧`��!\J�B�U��p�"�S=�[� 1�9u2v�t��������k�����)��5k��8�#p�:U�7w�A���zT��@$g�Z3.�D~�3�������R�,ƅk(������yR�3]���NȪ�ߎ�f�x?B�-�6�`;Af�^�m���UP�uO���<��g�b�3�b>����`$��$dz�Y��6+Bߡ�8!�u��h��a�5�_Vv��f���l��V�J@��%�}o����t꿇-��B+
��N��6���D� ݗ�T%v8���̏ �9�1<7�hΜM�EE�	��|-:�uDdp��e��%���yԖk����H#�P����upZS���\}�Z�hN.�E��k���h$��.m�kk�2+�b�_�z��; ��܎�~k{xÔ_���T	��$��gp~��w�=�^葋��N|�̃4�y/]���q������N��M��N�E0����J����A��9��9JH� �8tH��s��?P�P%B?���}!A-FG�I
�����
��vԕ`Y�y{~Z��ݤ�����؈y
Aؿ�[ᦏ��b�.�sC�8�FɁ���z�����>����C��7��Wf:�8 �!�oo@خ(���9A��"�e�P�&�ݮ�1�H���֢
ƹk@p��5ϑ%[x���ß-�> ���s�$�Fx���6~��v'�Y��r��D|g�rc�d<�[Z�%33l/kB�O�:X�~ ���]��,.B�xd��X��Խ��^����run��H��_���rsH0g�����U	�~n���s�/K|�q����q�;�p���C{�hO����*�'�P��T?�r��4�BP�^)"���S=_�^#�:,�P� (��4��w�k�qϔ�@N:�O�����m��"���HZ�y��kG�GS�v��gFl^8O҅��1 zkB��__Uv�5J*3��%�6�]򈞉�cb�Uh����\�#�hD��y���=
���Z'�w������|�n��C�t�u@e`W,�Z��=��I�_�zik!�5浮��ƭ��Ds�K����J�gdBZڻ�i�_�T-�i�e��7����B�0�]�a!���$��2�?��#Tu��v���}=.�P~c�Ȗ��^�B���K�`j��%V���5Xu�I,�Պ����lw����bU
��Ԣ�4��/
�=�Gɬ�2���N�XAc��N��@tPѺ���ҏC�Q�V�'�6��)&
��p����r)鐺V����l$��T�Z�ɐ� ���\e ��A�����y.o�
���E6��Ŀ�iTM$�+����'	�
�T�X�|��=J���"A珪"�r@ԋ����F����/Vm;,����	J�7�?jQ���7a�Î@�G�Jx�!�#�y��&�
̊������s����l,m~�'x]�UzY�0�%^��_SL�+�?��<�>O q�-]�=��М�:��Ǫ�Tc��5?�����A��Ѿ�6�!~�7p.����9�y�Vg�_�!���b/~Irf[F�Q�����u���+4���3��K�m�2^`!�vc���I�N'�	������?�_���E?sH��>s���D�haC���bd�W�� �������؈8����OFs�Qs0�o+,_I5/�3���{���l<Y@�R2V=�?R���e�+b��-�f���8r�\"4�h���^��-�0;� ���h�i�!�	C�>�α�C!v��R	�~��T.E06U��h�_��zRp�.� �uܭ�������]��)i�,�jür4ګ�]1!*[�O�ŃA�p'|����E�+�ghN���2|as���`�A�a���F�$�L+�G`����:�>��H�W7�o�Xju��G�� X�p��q���O��������|���v]@Vl����|Ou�����4'(���O j<Y�'����F�i^�w�Ӹ� LɅ�"u���AB�U_�Xv_�q��0����6� l�i/+݊���b�q벨�<\�C�t;.S�����f��?���(���K|�$	��MGz/T���+�d�$�<��wZ".��ؒH���~��L�N6Cd��N�6:��  �z)����m���d`���J�Mʢ2��y�8�����W���L��H�oB0r��vr=�>/���z��t���Jpdf۷�50ǳ:]p�h&�8��5�1L�3␥mi�8x��E
��q��5)����I�tω1� �$�]���?8E�A`{��J��mepk����+�K&�K��k���\H����[��}C�D�_p��ii�[�Ƹ�O��뽷I�����۴�1�g�EbC�~�:���Y�\����[�Л�1��3����mB0���	&���ن��E	�1Y��V��#e��ѵ�l�������+��S�V�9	C��i�s���u�(�/2�<yA�*=��A�v2���uAQ���̈�}���U����NY�/���Y$;�����i�}�압���ޔ�1}�~5b���ۀ��d��d*��ۚ��6�H�D�S���z���9wL����r}�(��]�^�2Q�������F�!:�V���"Z�+����j����]��?)�`z��"�yܸӡ�n�[C��E�������D��i�_�Ʈ���1.�G��JF�wU���w_(k���>����%Ѩ6��P��u���\K�AqK�����a��{䒖���&0QM6ȼ�B΃�Ѷ#�*	Z�Ȥ��T�=��9�7v&���G��|'C7�� ���d���b��` �X�PM����(භ�*�� �;)�BHM�%��(A	��}�S���ڎb���A�p�@��_J��{XPZd�-�d�{����`��~~�JK��-��4���-p�P�,�|w5��F�A�A�!N�ګ�����#�9�Vq�{��&���C�F�v��5FM'B�R;:�z�n� f�e�7��'.�-��c2�m�8�2���F�_v 
*�	<�%gT���Hr����G�[)JT.�MFn�\�A�� :�E�Z��NO�����CXT�YnPQ_�����k{
�2П����j!�: ��F�dc��՜?�F�!��G������$�,�~�C!{�W8�!J�<"�:'{"����r@�i���/�}!21�������.i�֟�&�y7���������K_�։�י�Z���ը?-,aby]��w��k�h`�X����*I�mK��e��T���8��Q��&Na�����"[I�N��Z깩��b��f�B<ڃŷa�	��$
b^#�)m�;$�� �e�p�W���ڂ�P9��	�8�,P_��;�a�������q�)ЛWn��=���q�R�s��U眲#��`MET�n��R\A70�/�E�*?r���H\VيȄ�����dA�&u�c5C��qd�[�]�)��)��Z�a�[��s߭G�]^��X��n֡i�g��?��������&���k�8��~/�6��J����#K�m[�R�*��jJ�:���9+��\����ۨ!���iŝG�J�R�ǬC��}Tzya�{�>����k���y���iG[~����)ܾ% ����J����i�n��^��=����S�4�6iYf7���d~o������~R��Ŷs
�tQ�|MTn�����h=�x<����.��)��/��%�z!����ۉ��돰�Ȅ`�z��و�˓p4��J\��
`"E��B𿱤p�[��m��2z��z���N:6���6�"C�}��:c����A���pO���*��0����D�Z.:�}p�q�Z����z�엟f�#�O����V&NN�r����$�o>��,wkpU�5b��39R^^-6;��E96�뀎����rRP�$�������� �=8μf(�Z�+F�$�bs�)xL�Uf�+3�'�ֳ7�Y��.R��q����N���L+�z�;���qU�~�����*?�3�ImN�ɲ���Кz3~�j%V��u �����Lx��x�t�.��r�Ai�)~?�Y������/�)ډ��1.,uM)C%X�xSM�%��?Z����6���o�6�6fn=�Xe��)xke�r��ͤ��9즌�ki���:`W�a ˪%�h��X�7�!�_)�]���`�ú�����k"b3�,����D3݉~/��AO�Q!��+y#B��#�f�;p=E{=C��qf��1ԖrX�[�4?k���>�XȬB���j!�Kp�뭍Ó?h�>?�����YĿ�$k6�q#��}���1����O�j��/�9�H�
������`%���L�	�!h}��E<=]!���1)����&k0�������j
Y�m>��z�y�
Q�o1�N��7oa�O��KH4�M��S�s��kO-�tE�/�z�N%$7Y#�!��яq�Y���Һ���ɚ�+�<���N�� �9>l�	Sjm���^��H5B�'v���	
�#�o�:]��t#���s]O��i�w*Ո5�?��G�#F�6���������ڈJ�#%,=�y?�U�]���Q���Ih��(Z��5O&D*�����; ¾ۇ#)'VW��4^mq[9�H�6��I��u���.����i�>b;��8u���j�#�(pvѼ�@q�����]��7fPѸ��xIp�ޫƻ��Tg�#O~Q�tu�A��w���i@���rzk"e��x�%Y�_	����ʒ�@�;#��&[tG��=���ct��U�s2��Uߑ�1���ɺ��������$e�I.�>�t�N� V��+Bu��a=��+�T�Q���/�����t�o��g�P�6�yl��N�<�{�qhW�	��/<!T0�}�u��o��?َK��w�/r��`k>�V��({}/7����6 #�ߺ[�Ẻ���x�����B}�њ���h5�
b�eG���#��j:�J����nx��76��a��U��fq��A2�4��֢X�%oE=qآG _Ä�ȶ�R�B��Љ�D����k�x�Z�)Ԫz��w�tv�llL�*�A�`���lĩ+���>󌤷�-nkka��8FC�|k����Z���ml˅����������ڐ��.6v�'���(̿�V�����r�����kr���|,�����O��Dޔ��.%Y�ڈ�?#����g��-�EFI�%�w�F��A���y8K���t
�Y�M.:� �,Ѓ��C�L��[S�d���+@�����N�s���WS2o}]'w�N��P2_���m��;�Jpf��xCs)�M��͓����KY�jW����e���h/]� n#�� ߷^w��G �Y��-yg�pQ·���_�7Y�m�Z��UA7����D3)��f=o����d��I�Q�>tH�ӝ޶��t�>���*9jQH��r���~�'-CQ�vP~��[����p��ka�W��v ��5��3y��;�QPY���drU]��!c��+����������8���S��Q�Ѫp^IdLf����nM��v��������)����ӟ� ��:��������x ����I�¯�������%�֋[�i���8�$)���!+��e4�X�W���a�U���I"���S��Y����K��(ފ���0�&j�A��HBOW�� �@��.A葠1:8�6�)V���8:>H��bp�����mǹK���/A�$�o%a4�q�c�+�M���,�&P[��O�e�Pc�ՒP}/-ow	�O-#r��Ǎ�e����KKɋї��#?Ѿ�y�L�J@!��j	A�L�Q�ן��6|�C�1��&'9o12�kX22b����� �p�;Xu�c�Gf� �8]5����l��bH����n��D�%:5,W!�b�~ 4���0��3��"�A�� h��Q�Ɠ����J'�����N^���'��H%nvlP���:���\��ڏ�CTg��	� ��|�$�?��q��f��Éܻ��aף������U�vU�TD�`O�l<8��v�Εbړ�&��|)���E�2�Y���hǐ�����1]�bD�n-V�<�*hr���E]��S�ς�	!��o#�E��u|.�6^(��G�>^�����p�?9}�U������ ��a"&J�C݄0�r���Nh�g���6.�����ߝ%g���q����ɱ�=��6>�Uv����)rF�h�:B�XH�,D�+!5\����B��օ�������-����e/H�s-O�p�C|�.��7����f����P��W5?�k3F�WX���gO�@�db�}�O#�N2�e}��ޯ
�f=�px%)OH�H��u��!�w�w� ��;��ݟ���|Hlk�J'�|u6�-��^�����P�#<`BC�W�:��ϳ���#0�x�q�.�M'A�,�]P9m���_�y�b����B}+��6�742�O3�Z��Ni�������L�����X���D���E����O"V���Z��/��{��6����{�:��AyOb�-&����2U�;�\>|�c�ʧ?���l%��4ֱ�#=Ϣ�c��k�A�=�K�.��YR;��2���ǉ�z�d�@o�2�,�����L�D�W�A�y��ք�d֨i�"$�ڊ:4�ĥ�]2H-��
�eu�����E��ݺ��'=p�����>����$o�T�ERr�*	H�2�U�o����̔�����VT�jO�?����Y��])��p�����D{KN5~��{e,4�o���]J�a>*�Qyk���wt��j���f��N�tJ���n�@�t��/㟉�<&Z�%��bm�!KܥR�TW�g��j�:�n3���+�S_��c�YqA�!����ѻw]+�H��C�U���3Y�1��^@��fW��E���Λ�:�k��	����ǒ����q�B��:�k�K��s(�'��)���UK��q^��<tm��}!�t�75�Ww���fd�ya4�/��4�x:z7)��V�-p��;ᶕ������?�fa��CH���2�r�z,�0b'�L|�6d�2 r�_ۦ����ν�ٶ	X�2��{�H �ϴ��;u�D' ~���j��5$
[8�qK�3fLb55�&���i��/�``�w���
�O>�п��TJG7��7�*��/����8���T��V��\��f�����ԙ�Lc%~��Xe�����&�u�O���Kn�9r�����L����S�����-��ښ�a ��	����������!�����w���>��թ��sf��^�V��Y8�$<c�R�V��\|�����;��Ư;5���Q��Dމ�����.��0�)5��m�@�����l���3^�Aw����skz�j���O_�lC��爭$�0�d.ͮ6�G7��{��xt#�d�x�Q��q����[�W�� %n�i�~)��|�ڨ�<���5�|ގ$d��^���P;�y~����{���"�}�)m��WZ�qи����y���e��oYO�4�J�z8o���0�C2w+K��8��;ɸ��Va!m��H짥%2�L�u�� &
��I:�=���y�Y� O�߬��`4ʽ��
��dɡ�Sv�͍�ؖH�_����(.nBQ�vH����=�)�� �4Az����[W�����F�o<+�������l��6Ӛ\�r�sf\��;�<XS��Q�*̈́�1��
ر��/�Uw"M���B��?���uֱzD;p:�k���1d�%����{�N%��å$�mJ���\ 5��<)ۨ<8*�S1S�G�2�����'Ŵ�3�l�m �B'E�u=n�� "������1��͓P����sd�����eߑgt	 {�ձΏu����<#�t�	��,��¸N�-����5;��~�����uHT�3�2�|�z��_�X���^$57�J�	vQ��[ѓ*��zq�}^/e���"�s��_��������t�VÏ��5���.ˉ?�������DF>\>�ܹˑ��:s"Y��N4���������Qdzʼ�V�Ks.���f��'��J�{��S�!p����&^㻟Jſ�crd~�V� ���i��z����H4C�����Fı��mp�n:��/�O�UАk�"��ͧ�95�.{"�q�T��*���P��P�\HS�����fI
}rm��']��Y3/�_�ꮰ��L�N��S Mt ��0ϾCA�$$�A>Yw1x]�Fm|~.�����@�{��=>!)��ƲL��$ѢUh`��a�$ή��D����`vqP�.��!_��+x;�jn��E�%!�m�ݭ��e�0F����A*���+��y��I�B��pf٬�(F|{O[5�(�`x���v����`� �-h���F�ߋ��U{C�5�\����m�k�C�����}�m�7�om�"�Z�q��a<�r��Y�:���m��;1�r��� �n r��s�'Тپ��@���K��FSSِG$3�v���*��P��I@��3
���Y�C��F���ti-Lp�I��[��$���5=���s���~�ϵ��(Va,AQ��Db�ݯ��ǋ�$��ˊ���7�1�.:�ܵ3�Ud�ئ�������]ܟ�	���4Uv��\�Ý�7�6�ѥ�/P����a<|����Ϥ�:����s���]�/
�4R~(E�*��U>@�ݸ[��K�[Y�ѐC�b{�-hO�P.�����غh�[R�-I�+�qwфi����vI�T��Խ�iQW��l�o_i�m���q7��=�d�=\b1�����jQ���*L��+�de"��dsr'��[��{L~�u~����{��Y�	9(ҝ����ʿ���k�*V�c�7���Nc@(� ��8��-�
-����R��Z�K:����h�0��b��^S�<�0N�5�M�Nq��2�*��A���p�뵚�g(1o�s�CD*U��'d8�H��h�^� ���2�G��z~}�@h�X������D\f��~%ˀi1k�3g���Ŭ���0:Y��Qf����A���_�KiOp�a�6�DAM���2�cq�`���i��V4P������D���g�-�>l�����.��÷��%n�{��%���5�mx�͎}��T#Rn��.�$&##����=��B�L�����X���6SVX��BT�M$����"J�쵐0�������`�|{gŐ�^�-��@����_^,���D�w��{�%z�a�x�����z]=RP�B=��ｲ+:Q���9�S�*t��+���VD��xL��Y�h���<��(i�J<�	5R�l�
���ݵ��^�_/�n��9��p������==�H������92pm�����|�!�
��>�_<,Dͭ����"C���A4�s��a�Jx���=��d� UO����>����+Z?�<�#+9z�7�&��E0g`܂rfar�<��V�ۤ)��6=��X�q{F���3F:vD]�|P{@ܦ�W�@~�,J���:�L�#O;�w�/�^�m��h����^o���2t͆�P���9���3N��8t/�)6��t�4�;(��r�yl��|��z����m�l��V�|�9�n���]��4&����o�����=���?�ق������R'!�t�U 
Wk]���a�,:>t��py�5.�����5�T����(�f�]����[�k�{1q�@�&�YN�HP��p��'{k�ɒ�m�K7��# ��U�R#D�aF:�$3A�j�es�?��\�P�p�C\:�#�%}���[>Q��<d�D��p��x����*���S�ո���c���dA�Pm��R$�z�L{V��U�k�0z�Sx�} �tS-}���q��~9�O��p�?��pMm�������-{d]��K۬�G�-qD� �KGcy1>I��ҁ�r3=9ͭ���L�)m>MP
��*������A:�ˠ0E�n���c�H��̓�"\E�����Kz~Z|�y�=�$o<6���P��WJ�Wp!�G�O���y�,R�`���
�a�x�ыG;=��{��~<[�����a#@.���ԗ�nt�w%�Cf�1c��w͌Q~*+��Q��"�����O��ǽ!}*���'Pn���X�$��[01Ќ�$�u�,h��PA�o��� _��E�Boi$��EEO2�+p���S���w�
�zD�;�j6ķ�*9��9���T�pp?Lo�d<�sMY�	�{N}s�n)77ôA���-$*�%�	�4C+r���x&T�#J����[��+������l�5r�,��~@U�|�{��,�dŽ���7�@&���-*�0�S}����t�S&H��&P�#��v|�GG��vm�<̥�i5�@"�Q����2�6��K@���W}Q�٭�H�Z�/²Te�ҡ��8�{k����]����&1I1$S��;YYdy����g�\}3���*�g��?�G���,&���k���V]�2| Q�6���:@�oJP�VO���T��ϸy7RV?>�ZU������GNW�ߧ�oۥ����Rd�~�Ut�R�ӟ���ۍ�E�ߣ|
��z�}GXbҸY��F�ʻyy�Af<��Vr�>D>��|����qL�]�'�?�п��H�k�"5.P��-�6Y�4��u��	P��A���Z�xp��h�G>	����*�{�3��ƽ�+F�ŵ���FL?����PA-:XҬ����i��=�bDu��r [RH�r�a�Y���R�0��0��27��<7����N�P��������|N�g�P�44"��sT�i�߆o�J�@��N9��A/�C�u�4f�?e��
�����i�/��Ӆ�2�W��Tѣ(����^Uaú1���2-Ӿ.ɝ�:��g���s�F��0�g5 ��|,�Oo=B���3	 ���(k.H*�z�%�9"N%]�WV�m$Γ2YϦ�YVSUI�O�L_��{�t~K�j�#�4���1�>�����E�P�鰑�dR�b1~T]���,{�"Ѹ/���xr������s��8��$0<�Ii�(��a�~R���r7=�	�I�$N���>��-tס�^6����2
x?�)C�U�a��]+�C:�����ɑ�SV�(�m�����y
����Ӭ���Jθ{0�z��@G)�X�l��p��|�loͤ�F�S��{eƾ|��0ȟ}����/����x�{�8>����=�l�5a��J�& �s������n��Y4��
.,N�?��� |��!�mS�p�����>�%��iv�����0t�ڗ�1��� ?-F�r�\n>� :�r�Q�^�hF-�C�Q��D8>���vS2�fZ��άP�`��7U�p����Žg�����!��^��]��ކ����҇6'�]��	����&��:��6���He��l��H�P��̗����r	�^�;;,�j��]M��;q�E0���M<���?�1q���ɝ�:�Imz���Yܑ*�Z��N�?��y���hF���W%[=��`�q��.j�?��b�I�6�.�)��+3��g��<��^���,\��4"�A_�I����H=�ǌ��U���aa�);��_���ViG�G���K1"�O����9Zy��c�\�S�]�>�mˢ���ڊ���d�?�ᰥ������e�������B�7$� b}V�x�.-��_U�X���O�ݏ��.�x#n-@m�R�v�&��K�W�3uFp��S��bT�K�j&�X�!gh�z�ɇ�ojs�)�!�i��]���C	:xА��bKd��Kr��M�n[q���#N�N�COͣ�Wz�d<�����s��\A�_�kd�rhݽ�ja�:�$^�y�"�L>l�d£����Ε�4�j�(zϗ��+PCK���E+�O��G^�)�9�b�kOm� ����rwߐӆM��x����=�����$lff�9��z3t#p��٦�����,拄
�-�ꙹ�2�l�(j֝>�~^�������\�ȩ�k�,͑�юR�'g�D�[�z��~cb�����?A�J�a ��
Vx븦�����h�5�3�t`�\q%�<͚7��qYcj 67m$F�-��0nP�K5�o@��񈷝�#�	�p�F����*cG嚁fk�?)�o.KC�yu�Q����,�gXPbG��x:l2���.�o���;52���4��%�9�!��OX���E]�.��mH��u^�Q9����0�}�&2U"�-�BN�Gk� -����y ��Zǋ�/ON���.��Z�@�ʺXW���ҹ��3��0>��:�O\��
~}g����ڿ�qP��2&k49q�x�m)p8�Ѓع�h�}Ub�Y�|Ȕ�wX�N�6�2��:ԃ�"W�S-�Kc
,(���5�t4Aj��E�4�s��iU�9�=�Y:%�t��s4�?/�*�k��~�_P'���RLڈԯ�RX�Ш:�s~ Wf�OG�+HF�/���Uh��B]��!U��`��\/Z���b�y�Ť���񥎝��{uf�-SH�<e}?������bȯ"�������z�iJ�p����(���y��#m���6s�z.���@ۃ/�#]�F'��`Aǜ�Tl��N�Tv�]u'�-�q����������_��\�>���ܺ� ��Eԝ._��,��o�<N^_j����D��w����\��`�U7�鐨a�8�#����g�A�v+���("z��w����۾/ć�y��E�t��/��s��Q� wq��uE�	��ώ�HV������¸��]a�� )���λ+����k�'����f��´m�~vλ������QB���Z���k�&�e�� ��kTHX�t���-������Dk���G�\��f׮��ź��a����IU��ǥ���T������ٌ�J����R��N�E����M�A���:����̠@�~gkB�'X�Oơuե]��xӊC�]u�5�`�l�
�(i�ݵ��Al��uĩGm#�|�R������4�g\'�:�rn~:� ����׺����6^
)q��oR>R@��]Ś�����#�?]��N��:s�Ѷ��{�|��}޿f8`��q�^�q��TP��e�M�x�;�I�P�9�Fؿ�������ɢ��D%D�uK���L	��`����˳*#�+Ӑ��3/�&���e�Qp��g�=t��
1��{��>ZV���������п�����I�ˑ��~��˛dTX8s�F�n߃ڸ�8l��4��Џ]��&qpRA�J��wD����
K�t���!�w�,ӎԱ��n.��zJ�=�i�
�%�c^�"ݧ�a-�v�k�O�`T�궷��9�j%�M^�eOq��[� �<�MT�-l��.֏�O��#"֜�3&�|��y������Z8f�譴�n����%�חD֧Z?z�x��A����_�]J��Xx��P�G㼟ԋ�D��N��cZ
k�d6��z꣖Av�E����)��IG:(�<��
�~��=?����i̠`��VC$�$DjB!룼o�Y��"��C����~�e�w��}�hv��(T����N�J�մu7Y��z��j�tZF>�`,'�,�9c��d�>�mڿR+y] �]��k���.O��5/n���[�v�����C0ռ.c��	_�dt+\
��x	�s]@� `U[_�ED��rVٝ'zX���� �������y��'������hv��������e>��:�i`'Dw���H�^�<�����l2�����e�/�������{�Y��	���<�+̋K�$+SX�C��b��:�,
��9���4�h<앝�SP����;�얈ڨ]�͓L�3�s�t�/z�Y F𠌶T�w��\�����U��C_y=민�f������ׇ��)���_�oֿY�}��K}�����=��0�I�:���
�	ඹI�l�{.̊��S��j{ڔ��Bo�z��w��ߛ����k���iwF��v	���V�<ș�y�{
�L|�^���.�_�&ޤ���Fw�����~9���ܴ{MK�0
���4%�]� H��:e��=SHT��GDy��QK{�ұ���1��/n�S�_p�n
�J��!�� ~]	��3���O��D6i�?Dw�d�=��;�^�:�;n<��b�I�3O�Ѱ����ڷN�?������n�i�ح�Hm�m��U�
�w)j����䱯�v�N8+3Ƶ-7[���U�E�K����v!���`e��S+��c5c�5�6Ųǃ�!9�Glt�GQ���E��g��k���S=_;�]���1��Sw�;w���Rv���A���Q��J����cMa��M��3�1���4��zZ.�/L�s*Ga�������i���<����:B֣s?��b�˄��\/��|B1���V�F����,�����:=�|@�KuM���	�����\����}y�D�	MIm���Y�7��M���`޷���|��wO��-D�8w�~j6��L�s��1�L�m�/���u��}�-Ʋm��[��4�@�R���N�~�X?��.�{^XM ύ����tl�_��g�'�,^�|PF�Hl1��/0WFx4ƥn�ל���^j��EB�{��xҢ^c4��v��f��=��j��)}s��Վ�6��@~h-����)˼�Z49�;к@��������MC�P[�>q�ʾ��t!S���|f[
�}_�� ����w��^���!���:��ܓglˑ��J����U�R��l����62β}Ln�&��?i��-L���/��y�lʦ�f�GԈ��%��*�J�\a�S-0�����|���vo�c?�a���*d��5#�O{s��1�i=���ӄ�^B१d%���1�+I��J���D�q�f8��RܙA��������=m�MA(��M����촜iB�yJ|Z4��"��e��֬L��bQ��I�,�I͵>JC�0q1Ġ'b0�r��1�m�Ww�Q��ګ�G��B��K�����g��5�`Aq�Vq�d����[1mtX�+�{���E���?��6'�u۸�.<^Ǳ�o������e������9ei�N��w�&X��e��-U�l��(��+��D�Vtn��a�>�8�}�Y����
�UIZ:|�m���.���	=j��Ғ�k
���19�u=�F�`���Y��E�z�ׄ8k�m/O7e��O������&���x:<��9�8^>��BwZ�8$�og��b��zپ1��O�A��i��m���[3l}�f��g����a�^Q��d1�t2S*Mإ$���k�X����g��jkꒅ=��S]?�����dRq���"$��tv�>Xh7��(G˼1��i_`�@"�K$_"-�N#�$P��ϧN��}�| ���т���=a�m���w1-��4� �鉟���v�m��!y��d�l�!�*߻e5��=�Ad#W�k82im.��s�r���&nE ו1l��zu�'��}�q���1��*I��.}�!��2o��\j���
�������В����<�Qot� ��%ѷ�ḯ�beʟjlk���:���s<+UK��S�����u�e�,���������B�av^�^i��7s������1��z֞�gt����u��lbpaUo������C�!�O��Y����!၎D�ZG�,ז&\�`a���(p�&���Q>�C�Vui6)�W�;E�T�Rb}���&�`�?��äv�}ϝ��F;'���=El-x|����#+��步�����!��D��밍'kߔ��6 ��%b�q͜�pՍ� ��J�"��B�v�|��3T�x���,�M<Tq���!Q�����4;6.V	���]�3������#�m�d�{�3�Y�7S\�b��'��s5\���L������"��wǶZ_�G���cL�sw����pk��>�nf��W��]륻�u'?��1�cD�.7��L�DS/�)�q�
<�C�/3$@���5G����r�T���fM�J�?�S��;)��t�k��I�.K�y']��;�����
&�7�@Y�ԗ�.9?4�wz\&���U�'xz����սX�,��<A�/mh5Z-���mR[I�&$�=����<��̖���,��C���_=*��|��CG:)v0o�^�/ǁV����^b�|�:,�ó�V�u���Y�����&��A���Ӷ���]>��H��u�m������N�h��$�[P�X��,�_�.�h�;E�z����}�_�M5�F��\�g��޿5���οf�<iq�F�V����l���z�ȸޘDK]��*%�#��Ȍ�F1_η����~�yx`
�<��R4��O��%H[��ڟ���B��&hu;�XPe��_��J��s���W֟%�[i	���n�C��xSs�D�W��h�dQ_���5�}�8�-�@3��R�]=�=��s&Yҟ��C?N���Z	��+�`i��r��!�!P�Qo_z�W��L�q�8�=7V�筓'	�m9�X�]Z�^|ڳ��Z(�)����ď�7���T�fX��*�J�)�� �aH���� �aV�.��h�r�m�mM1I髐e�c���ҡgLi\vh�&|b�q��]�Up���FA�7N��T��̵���}���T"竻�����cy�5n�L����4�������\���=�m�ӡ6�NF��b��W�c[���;��tވ��k�*/~X^-�ӳ��55������ҼC����ok\��V#�!:�+C���<5!���i3~�'Ĩ��@Qe}&N3f؊��^h��������xC�~�T��9�F��X�ϊ�{ӊ����9n_z��sN�N*�K����[��g��Cr]��W�U�'�}c��66����L�aE%dB�J��c�w��Hg�6�f�%�����(Qn�w:��d#5�g5Ĵ"H;=B�I1�|s�4
���0	w��nEyrm����`Hs�*�n�-RH�DLܺo�y�R�M��p�dv{�r�A�7�Z�ߥŴ��ݕ�L�8�|��`}���d�t��B���\�S����Z��V7����(t���4�?�6Ȃe���B���ծ��C������KA�C� �+�9�Ϟ�(k����Q��\=d��g��\��z3g��G��/K�"zC�ɸ�wq�z/����b�I�k�B�7���\����g�ab����Z��w��xM��է���K�?Y�t���mG�|.�ۥ?�^�
U�W�>֮,�{��`+��6�?�^� 5�j�k�����?~q���g��rI���'��$f��/��m��r��K�5o�\猫h�0;�	�|�����(�xxe��8:�=@��]\UБY���3�����5�^�����V�)�WF�_"'��Qȧ޻��=�cB+c�cm�XxY�n����:�Y�^af�t�| �j#���.z���[�W��O�z]h5尰�k�%仡՟ݪi�� {*C@D῞���ޔ��4��7i!�^A��s XM�S���?�4�ܲ�<��1�}�
5_u
@�e�dyG���8��+z���p[Ĕ���.(��T��L؃j�R��z-���G�~-E�i#V�̏תK@�P�/1��>�dwm��0Xއn�����՝,�/gꖶ��9�@��������)�}4����'Hv�u�Yv����Ϊ�u4�+����F=m/Yb��^�Lqv���}��Meb�{����-���
ʳ���E�x�6�������2��I���-��X�����|ML?����~�/����jJ�L�S�3We��3�@����H�)@�oX��/t����%�G�����Gd����xkw�:ݹ"^v�����$������^̀�X����r��$��ψ��\9��o��,!N�J��5��:c�;?:��8!Ѽ����\%�w�����A4�@(�h.��	��>Z<Ϣ��ŉ��,���_��P�R;':�Ӥ�@���cF<����j;;]}u�Io�-��ʳ�Qk�N�o7�v4�Pp�%>C#K �6c��r����s�-����t���'+� AC�q'�[N�E
�|�>���0%NOA�X�[���3�T�?Yj$��L����X�=�_����r��3ϵ�F6}мI=����>$��Ԟ���3<)3I�H�u㕑�������3���	d���B#5���������6�
&0�n\ �V��4B�/��?��DC=�����+̮C�Z��$��y��R��^���X'f&i���ZD��u��Y�N[��S�(w���]�k��z�3����p���ε���r�}���H�Ii4���IL���Q�y5V��7�]����M�� ��V��m��H��w׏�d���ឥf�Z0*�x��莅�`kg��DzᇲGWe�4:�2���;���ݑ�X[�%Y����̫�9UE4��[�ح�S6�T��ON@�u�b�x4Ѧ���Wf�@�,��#�W����)�[����r	SpB�l��!�he���_��qݽ2{km�mX�[�#�W���3�w��{�ӛ
��;��ҳ]0�Ա�j�oR�Z4�T>"sMn�N�l�Lv��3'9�e�_��=Dyѥɻ'�4�;�����E�9��[	c�S���#�0��R_E����~�K֞l�J���V�8m◚@�Eˆ�W��њ����@T��w6�D<�?�q��Ҧg�)C�+��F�|���5n�v?��P����F��D�HĠT�7o9,�#�rܺ"�-�E���]K%S�ڧp�&J�:*�ٶm|A�@���4����[x��\�Ygj��ݗ2��:���� YY�������.+�B^�������'(Hpu\ ����h�f\��
��p�'�/)�	�w���j����Rt�#�޶naY�t�m�re�����|6k���Z	���C�.X���!�q�$_	���9�R+�	�&"�8ƕ ��b��.o^�`�@`G�V��ha�,?Q+��x9}�k����pYn&�,E[c%.	K���d��)�<Z�^�"�E7���"�}�� �P,	lM���/�{+�V���}��:J#��z"��n�v	6��f%}5�=�k}�"6,��b<g"��U��8�nz�U3Z�y�	q_�w$�)��$I�%�=���+�g��zd/+�,���0"*��q�ʛ���w�씴4�+W� ��d��'���-XW�A�_�!�1�/�
����x�%q򓞳љ��[n;��\��zfd۟c~h�*R��N���Z����Ԋ ��NV�1�<K�	�;��ô�4x<�z �_>�B��cd(� c���8INk��5�6Z<�X.w$^��:�İ/���A�������N��%�B/矫Ul�%)+<n�4�
��&NL�ll2B�j5Z�^��k�\�S�����g=������ɉv����[��م�2�~�/λOK�ߗ�J3%!�e�Z3WT{�M`)�Mov9�(�*���H�d�n	ZP>���oc�����:*3s��|���VGo���|���	�p'QWY����ŋ%�_���#������,�-��]�R�l�~�E��L&�Zt'V�Io�U�"&b���6%�;� ���ɩ���7��B������{u�Z�O[�'���_F�vy�f�K���_Ӝ+_P��Xz�~�A�%�������2�$����'8
��o �?G�ͨ\�8���,����S�um4��D)��!��B��{�|������[�k��C´W�yю\���zt ���i�$CA�T������@�@���!V���䡺����V��:ӝ_\Ǿ*3`K���=+r9�g�ǧN��<��3Ԭ.{O-�dq��"^�����^����u�!9S�FIB�����:��vD�t������L�c,ˈ��_������`3�������|oP-~��0[����љ�����.�M^s�����4��nFq+�F�~�t�B�����{/8�K�"d�� *Y���D��C����i8Y�ϹMsᬨx���sr����B ��.�E�Zڅ���nk��y�NA��DC�]�3�e� $ëLT��[�yb���kPc��(~ѭ�Y�)!<G���B	d���2\UG�s�9�s��T���y7�.#�����������%�}�i��T�5�Ͼ���l���Ło.C����v�b��w�V"��9Hz��v�s۸B>����x�.n��?.9kj����=���3�W��S�&�W?��-|�$10s
%蕃m��gy/0,�o�|P��a�����v��_� ''���".�,��+!��Ͱ��ó�c�����3���)��wHL�jn IOvg��9�N�5��h^z�D�;���Tf�0�.}�ka��M&lP<�g���S�-���;<��eG���Ufo�ށ�0�D�\m����Q�Aur��r��ʝ�3��MuG<6�'z�S�R��\��[�5�Hf���#G�=;,�~ްPR�V;aۭ�S�I�I�}�B��S�e�2tj�2ؙM*7+�a:m*�@W���bۖT�w�Sb�Ɣ����q��{ʍ�*�	�/<
^ι�.����@t$�kڽG����14�B[	q3O�n��?�QZ��
�n��ܯV��R��;��/����C82^��.MEN�i�I�E�9.��'��gԡ|US_�8�
�w�X?��=��}��[��]đ�o!}�?[��~����W[?�:�r��].һ#�cu��-�f��*&$����>�>�d����f>���f�bE<f�I
��.`�'���� ���g����,t=�*ryL�9��R7�Q�j��8�Sߝf57&���z���O��f�"'���?�y&|ҊW��U�6�N,L�9���pJb�y�֐�%���?Ô�kv���t�|��>77�G�������],m�%�$�� �ȟ6�vӥ��)ޡ�OP�zVɁIo��E�)�W_i�H�2򣏩�@)��:�>s��y������1�L���ۏ��|��@x�����B���Mk:R�	�r3E/���\��Zw�������ۈ���n��H@Ѫ��֨ln:��fegΖ{s��C�~�¼sfE1���d�,����o��g����2`�H�\x��}��mc+B*�'�D{4d�s^'�8���7A5?[�+�|_���!�]G�}8{����§S?�m:�dSi�����v��f�h�wV�1\U������V�p�Ys�e+k�&�;!i�p}�,D\���n8p_Y��Ӆ.�pl��-0�t��J��[�́�=�`�����,�C]�";�%yuu�p��TgEV]F�G�հ��H'_mNE-��>�Y�G:1����~�[r�|3؛�A�`��钒`�2���7�����������ru�71	e�-�o�h�����r9;/�}N��q!���L�a��U��39T�� @�&���Sk��<�� 6�)��!�"d�j���6>��/mgsQ��]*�Iez�MlN��E�& �F��Q��{&E�nmJ�E�
�YvU�]��L�S���o̊��T=���<n>q ��
N����[�]�aN]��y�(��R���S�S��O-khwi:�v�T�g��g'���g +)�ƣ�q���&^��,wj�3�������ܲ�Ӻ^��*0[������+��n;�p�K���sL]<�ԖӢ	�;a$�*�n���Ȟ�vu���=��s̭|a�}�j"����އ�_���y@���B�5�Z���#&��%Ã\��T��6�%�ɯd%XuB�4�Ӥ���~�g���Y J���KH�{�j�n}\,U�X)`\g���d���Z���]^QAQ�-�տc����[Z���EJr���׮y���4�6�%|g�p�M{�ݔ�y'������i��,�Q�>b�N��Z�&���&�gѬSCJ�y�S(wP3d����E�%�وg���bԆ�������;��%Z��%�hNDSè�Z��H��'	�%5c�1���/��S�}Y ݐG� �c��v�݈I��1�6t[�h�%��Z�͹-EqC��vm�ra�H��Ojp��)S�V�!pR�6�N���cj��޷��'굽�I@Ϩ���.�J��}��Uf���k�F��J�}��)�G/K/�j*�OW��Sڻ�JH�q4H��T��i�'� ��� �㙼m��8���*�.5�{�:_�߈$8��`�ƪ��6X��.����@'Fv���A7x�������rg-u��\�j�c[DW��h�#cC�LV��ͩqhI;8��X�d!x ��A2�8*�����?E�'4�ǁ���J��j�!	Z���v�$�;���J;\:B��W�)�\�܆���gnSo̢���j�P,)��M��q�\o�9�blwo�۟E�N�ʏ�;��;\�b7�Q�?�z]&k��Y������)�ñ�uuTb��l��S����N�=�r�u:pL�I����ݮ<�._��R�)����m��o�sP���4��yt2qT�j:Obh:���I��dGƔ�[���t9,.�ͪ͝�Lo�T��q����M�F���5���=�a1�K�q�N&�+�f�:}ײ�����µ�HV��
9���"ȓ�d������s�XI�R?�������֓}��3G�3n���k��|����ReʻYw�b�r��fl�Z��Q�$D!�]��G�O1�,Y��xw��Հ��9�\�5��/�ػ ���Y�Iu��Ʃ)7UU�}k�S��Ѡ�n�>:B�Nd�����o�h�G�*3H��F�N�������|�*�y�w�����FjR�>�u9=Y�G�o<��qb�Ӥa�D`�dYx��V0�a�)��#���W�C��[j��jl@(�]�
��T��Z�N�X��� /y\dA#V�n��8}��
(����D�;��hE/��#nЭ��ɛ*�"�/s1�/_c�(v]�?��7���_�h��t6����`z~�fߎ{:�U�tag���s�E�m���Y[�7�E����_~+ٶ<��4�K�Q�u%h��VH3�@�S#v�a�����}/Ҷ(�K��Z�������mG`�K4꼔����+&�v&Qy�i��-LcIL�l�^Z�yZM'�����w�~p [���u":�O]A�x��QO���k��nօ7��&U���cM�f�Lu<c}c]�B鐘ji���5��L5yd!�1�N8]g�n}C����}NX%�Yi�|6+��h�_=��0�mgzkB�P\�b���h���M�
4�58nEU5ߤ*��p��}<�������2�(Ә��^kO:Н���g��vW�;�I�j����
n+�E�f[猗I@ׄ(�����6���*!W��3�e�n͋q�5f�t�.���%0��{Ά�!kQ�J��-�����	������E��J��)�!T+Z����� E�%E��V��S��������/%�&���լ-G����Cx��Ҋ@./Vv������*��T����9�;��1�i�6��G����I��pS��@5��sk@N)+-�,�ĭ��V��զ�:���x���K�C�g��2�5�6�K�+�M`�h}�P�K����ف�T�%֖�X�vo�]%#��:�mg
{3;��N�C�	����t�BQU��nW��G��k���g���������$-�O�j�?̌�!+6J�!�o�L�nzk��躰���/>�|ioz�f2���Z�y���s���rifQ��'���5�%p�W����e^�_����9I�֛���
#Dc����I@yM׎,�������������t� - ݹ��"�� ݽ�t�H7H�t�� ݰtw��._�<�>��ι�0w��n{�|�ˁoQ��w=�>^�ݰ_�SR�wU���f�)N��t_9���qʖ'�QU&��}ˠ}\���i5�Z�M�)^���tL3E/p����H�kJ���w���C��(f�8]���O�]	�}CM1m[ ��q[������&}�Fۃ>FBǻMQ�I X\Zw�Z���y�Mf��@+
ە�(���T���9�^�U��`!�M��Frcj�S1�§]�h�Z�C��Ϸ�\�4㿄Q�Մ)Q����.{�2,Ŀ���R�g�;7Uy/����y�.L�t�}�����?�N�n>xqX0����Ŵ���L�X����:#j��i�&���5���'|�{f]b���6��>��0!�]\�\�>
A���)H�ћ;����W"���փ�M�e��ބ}z�K�����09j�l9=��3U���"#%���t�p\�DG���C�Ƿf�,����z��R�����l�xRY�ds%�`�w��32g.�y��FԚ~�B&���;�Y�yF�.cӕ�KGOT�K^�ڳ���T���Q���N���}�v>_n�8-=�2~YY�*���+M�絛s�.
#q���se��2v� II�f��b�
���Tp�����`hQ��՝��e�cI�I��/a��D*��<����PO�p���d簵��7�TB�F��CR8�k�ŸC{W�� ��(m���Xxg�2c����3���"=�@�֔eD)OI�x�ʦ�֖�x�j��I�vc�!Ԗ��5ugT	�����
&��O�ug@��=Y�eC��m�zH��{��iB���K+,§?���9A�;�=���z��~ꀂ��iTԍ��y��T�,��Fa����0�^�9m��r��Z���<��\3�;�xo����K���8|�╺7��"W޹�d��ڥ!=X��+b#�W��+Ⓝ]|h��rX��e�"�=��#�Q8�i]5t9����o����J�䷱l.&1E�WG�`�r���S���}cȭ`��m�u�W�B7@�E�6%j�~�a�fpm� U�9�Di.-���ˤ.�q(O7�#��fjzM����#A��R7�'���?��D6Q�Z�5X�t6�@-�I������ɕ	�)Q�co7��e��r��
)�	�JI��O!5iu~��S��w��ѱ�*xQj7�)�?��U�o�Yڳ҃d�\ƒ2�w��&5U�L�IY_T�B�uxx��2<�dv��}��&'��q����0����D�p9v����^>35�s�{�������Ǫ,�$��b�WZ!���Z�)d-��V�;���JW�O�+�+��Rb$6*>T���no�������o���5cHCZ�3 �>�<JF'�oy����z$V�WJ��D��@���T���L��
�[��2���p�P>W��:~�'�T��TM����d���jVs���vJ��T1���\ݛY��CǛl����;�j6� +7`n]H�]���a^6ϯn���v�PZQ��cœ�~x[t����E �f4��z�dUۂ���EU����Nې��F/.%���S�����U���K��U��0��ġ=t�f�֚I��[���l7�^'m�'-�5�"�$zZh���c��Fi��!M&�1L΋Y�ȯ+�#��Ml##�FRko��&ص�ԃE�)��N��ͭ{IS(q/���>����!�W]͆7�~��O*|;:6:�ܥ����]pHTvH��/�zh������J�	˯=�N���D��N|V�R}�f�J�Z:����fW��[��*�F�S���kw�yx�/�&\7.ə�p>ю!;o�W�U`��K�7�<��瘯u��.�d���P���3f�Gb��r����(�vw$j�s�S��WݖtrY\dK�c9�=]��" ��`�n�7���:*�R�7x�1ӏwV�=_�&�M"
�����+ҢT�h<k߂�q��Gb!�#��P���K]U���AÄ���:9Mǈȭo�T����Ԥ��Q�߶-�Kn���Ro]��\�
�Í̌�b��&ˮ�����w��z�ZY���X>:Q�Ⰰfw�XϝnUÉW��NA:��Ǚ:X��JXH�7����(�bWU�ά��OF��T�葵� |"��vA,O�K4=��F�$w��SIH,��7�H[bo|Z�~^h+�H�UM��P)s3(�j\�B�U��o!g��HQ�h>0%+d�X�_���bR��0ӽfl䴏��dV�pρ����p�9�-q�$)V.sr}A��r�)A�׶�qJ􌠡o�>
!�{�'uA"�=(b��]-#��)�Q�^���c0�����D\h���hu����eƘo{ת��ڷzC���V�RH�&�R�5����IT��u>��r�� ��_t%����iզ�ˌ�UX'q�4��yQ���
V)��?�Ü��-W�|�Z�	��X>١�D�0����p����2�TmX��Xq�<�BO�nW[4��m{8�}7m��^�F-82^����3���FҢ�]�γ8rl��kMI�(�{�,�]�rNvY����[��$W��=�>>A�<Êvj�t^�N-~�Č���K�tM��1c�oA�4w#|�w�}�S�`��=�:@2�;�����7\ҍ���D�{s݃�T�1e%�ջ*��+k6�m&��G�*�ɞ�|"nǢ�4y	���a�>���~}��C�F$����m�p�d'�|��fP�V��+E�'r�����r�߬�B�JRP�YgS`Sn�%.�8m��g�[prP�0bJ�����״��������TY���ay[u�X�^۷�W����)R��l����~���~����cx]�E�bn�Osj	E��$��4]�ct��;����	��#����Ȼ��42�W��ڥ`����� ��,�S73m����-2 �L�z�>��4؛�J��t7�uy�t~�C&��+���T������|7�,��n�U#����.x��Q�d�?;�5��n��$F��'�0Ԛē�:��_�JAUڒz��b�ױ�������`�S��RH�3���١�L����o5�UC���]�����ާ'�ё`J�s>w���*~�� ��V`�
��A��M�잸~ѽ=]�v���P�ű~ܳ�j5�F�����c�H�Q���=����כs�Y���}4�l��Z�1R�{���:ͨ=N,~���\�`V �\�����<N�����>3�IpeFX�{��d�֍ϧ�!]��m_ޙ��?��r�]r5Վ�Y���-��$������΅�����`��ڞ�u�T=�y7y���x<!vjbU�\��~�B���{v��=��-� 7v͸noS����QD?mo��J�E�&t\����ʏ�N�����a���;��݀ݕ�k�E�ɉ�˰?'0�	��&�sD��qZ�Q�0g��ڭ�T�j�OD31�p�2l]�:�#7��d_۬lB7�+��rs�4D�m��R["�Z]�A�5R�w�N�jH�飱R���7�[+O�Mz�oC��	�
�1|s�	���b����eS=���;�s���L�&���H(��k��ڬ��;�+_)K��}����W'0ae���9kp�_�(��$=!���0Y$t�դBT�����x�]u�g)�9��t��2p#koAC-�� ���*�׃��/4�,P���p �ݶ�	M�m;���6I	��>/(,/�c�Pͷ��A���PJ�Phc�N��w�-kݞ�A+,�SL�7 �-�V�u���@�Z�9n�fH�W�.�PE*�����޵i5�_�3���i���J�2S3H�b>y"���~����As������[������&d@�
|W�C�~��H���>�n��ڣ�Zbw҉ �~K�FB�$|>�'�@�����M���߹Ѩ-�qwE����敱�����ꨶGa�|�a���u{��Ǌ(��S�%#p��F_"-�>�|Q�`ց=�=�&È���s�<�#�j"u)�)�
��s�ķꐍ:�C��dg$O�d��|��H���Ŭx�[Q�S�/���D��.�NG�U�3®g����}��
��l5S��9�'��njZӧ���U�x9�q3�ð�K'������._s}�Я�o��[���q%�*�8]5�bD�
c����IFk��h
�xY_퀘�,E��ɷ�D��|�l�-=<+`p�+�̸[��FkXc|q�zwsR6|}����A�k\�����=36��+�!6��dn���F�{�|���02�xL�4��៷�;��A�䨤y����8��}ٷv�<���M����譅�V�̩�Ŭ������~�p\�p���'S��g���pd(�5A��V��4יJ���lipr�=R�z�l����U�O@�WOdk�k~s���M(�n��fx@�\[r;
�žU�~t���������_}	�<��J�r����W(��nai��̎V���1�"./�r��gk�\�l���lJ߃;�[�ikE3���9�"������=�3��2��s�@��-.�x�2�K�d��w�iA5�}R�y������a?�\���s��	߲�_���@o@&�W
c��G�Y%��A�`�����M�Z+��'� �z�9K���g��C�,R�����{=����Dd���0�<~�;:OF��?/�#l�X�
��O=U�L-]��!��E�|c��gXݢY���0��G�~���1e���C��ޜO���	9 ���@��`�7Q���-�%��f;��3�+�͵ͺ黄�.n�;��Z�k���s�D���-n�/�яz�Ff�Q�$F�����L�T�/G�b����>���ĵ�k@��z9_���㍥�f��u�����6]�\Se�c��fz��4ʂ���.�_��3ͳl�O��U���W�1�	Y��Ь�6�6ˍH�����V���&~�G�N��8&��r>l@]׺�p����[���e�}7&�d�@�&='��4��$��l�C!x���~�϶ ��Rs���d�b�2;�.bl�H S;QIIFS\�ko�(�+Z�l���4�t�q�Ϗr�#A2�1�'���a@ZS���=�3����:>m �?�'��I"��H�����v���?�J۲�Ү4TW�m�78u�N@XS��v�[S�~kY9\��lp��F�����U#�K�۴A�6��1P,
U���h�^��Y�r��/� `��"(@���xW$Lh_��K~cDi��F�v΍��>��pD�����L��)+ȝ�*���]BY�1IS���~j�'u/�XA\6-�Pi\��r��^��9#,q�-/4r�rp1jKe�0^J�����qT2�
� �Hu'��*��C/�RÕ���� o�3���s`?`���-;�(�Ȭ6x����(�[��"�̘~���q�u.+�rf�D��"���mqN)K�nyS�`��G}�7��e���	��m 1���G*�Mg��aM���f���k�3ML�ey���QP�z�#1���ǂud���@�ɨٞ�=���v�j�RҌ�x�WT���R�t�UX��8PL��`h�dj+G8�_��yJ�l���r2u$=y�����3�>�*M�ʬdV�M.nX{���j�]H�6�e��i�t�>�����7��:"�(�\�۫��ZI�!�@�8�!!J��TM̯��3Z��
gؤj����O2Z}�Z[v�KRBw�G2���D�=�-��U�+��@�7�sv�Ǭ�\˖[sQw�����4竞0��;���=����[�/��KL{p�=�#����� rb��0�8��`�A���I�Y��R���� v_���x.�K)6��Melќ~#* V$�ȟ�m���-����l�gU�/K$[�D�0u/!�
V���"k��tБΰ]�%�gʙ���v�g���]���;\4��^�.~:�uh1��$^���޷���7��k��$a1\��������%;&1�����:Q�
�<1�X��ۭ�K_S�L!��˿��񄊜k{k�̟��<�wh�K�ug*��pk����N�LD����P�I���� �W���l>�\�2���^$p�5����7B�.�`U��:LD |r��cft�saK5n���-h��k�y�����c�-�,nv�$ef�<�2��Rz��T��}?3�??��|N�2�qUI�������CJv��s��ᆓi&T"��J ��,we�}���L�)����tA����IR������������v� ���^7&;$��V�̡��& m��S_�����c3[{^�g���Q�h�2��Zg"7n�_̻\|�k�½/dO�t/�/2~o��W�v���ƌ��Qwo3F,��g�k	l� ˠ���QD\�������%�������4�<�l9F��yP�M��,�"���fa������vq�f�͒1M۶&A����.?f�֝`�=E-a�����E�P���X���	\��{7�� ����X%�^~��[9��	��C��K,J�0ܾ�&��*M��^���Hב`��T�dZ	ѓ��2�S����w��a4[Wb��k��k�u:w����g<���\��	v��k�^Q���T	/�ϙ�ݖzU�+�p���aW.�`�QP��e=���h�\dD��/=�9�������R�P��ӊ���A�8x� ��}d\�ՂHo��W��8�f����&�r�F?���λ�;�EF��f�ظ�_��&m�2���<�#^�q֎]�l�q����}K�مA�*%bw��֓��w0�-q�T+u��{��طp�J�ϯ+���}	��
t=v7Y�9�@�&�@Jh�S���:��*b�{�nv��PS���Y�І�ڕ�sٗ:Ɇ�Aa!�Z�K�ŦlW`��~��\ޚ�'\k$�ͩ���9��{�����~ċbU��ŷ&h�C�EO�R�y�Rs��d�����S���鉮C>�n�#뺞��_NG�P�Ҩ�U�l�+�r���H�_�؃���=`}�@�>;�TZ�o��r�e��Y_9�����*��g�t��p��:��(�ؼ��CI�O�-ߏW��lN9���|�Ao΁��ē�|x4W��%o������m����-�.�zS�ˬo�m����y�"@����z<�3�羚�`}����J�\���)�ff��N��82��i�ms���B�s�a�f�t�F�b�Ma{�|Ç���cWD���F��}*���1�u��7B���MV"� ���5��u>�<���)W2o�sn�"�P�����x2���YF��>�;u�e���9l�pHH���z��By�w�H�uA�wDx\���#��ӳ_���ZWfp�~��%��%[�V�V��&X(SL���{��K���.����#����ZJ��{����}���'��Nw5	H��duM_� �}_+��׬u*8+�A�A^sn��)R%֘�_��}��^���0������WB� ��`r��<���b��W��>(u�k̽h3:��Ƿ$9�:h���N7ᤦ�\n��ߋ�c�]�'hO����SB�v�x��[�L�j�]��%5aq�3p2������By���U��u���wj��/�F�I!� �qf'�݃ܤ_��II"��Թ�`k�v���a�(�y涆��@{i��T�Օ��?u7�vϙ3"�<����c�d���>"��#Zuut �\��Y�Q��4�Y��?�'�x]vk"�m6k�S*;�[���Ļ'~v�%�<�J�f�A۲I��(x�3��56��:�9�vt��{z��.+o75
���y�͙�yW�8��z��V><z���jY.���O�;�87:����jxͽ�R��R�P���zc���r�z���'��n�&�`Ҟ� �s�=���=:[ѽI|���jYw��p�	�ep�5�K8�����Q�����+2�f!�������D�'ܶ�PN[��D��0+�O	X����Q�R��o�d��T��w*J��������v�AY=C�j�K��`5~��Cm��&2"�����g���u���
ߊ�Źw�X>��_�p��K+{i|���{���w&���dc�Oo�z��ْ]�wvZW/5c�=d���Z^C����}{}���w��(OC��֍�4�~�hՎP2���<@9:�����F�?����w�I\~���)��/p�+��H׫���pCZy?8��e�&<e��Shh��ܺ�I<&M�|m�=���E/�O2�
4m��c1�q����j�����ؙש���գ��,%�bځB�bt�ޭ�m���}���V�k���j��m�-�'0gٻ�MZ1�,�ڒ���Ҧ�*|
�'����1��A�/��c���j�c�-���iz�\z��h�K�ª��K�"3o/Q��z��hk���+_���4��-��Q�̪���j@0<ُu�K����Ƿy�JJ��KֿV�5�+PH��s5��y�=����gΘwz�kSjC1N�RӦ'7��(z�/c��T{�*DN�rr�� �z׌���K@�M�e�bbqf�ã���SWzi��Qf���4�B��Gy����hq��M�@j�Ms�qe��|���?ߪ����o?̹�:�kV�Yt��۫��N	�٧�'�i�Tsw�Ҩ٧�\���p�5�h�H)��:�Įt�*=NN��)p�"[���!_+�AK�W3�f��QG����s��֟����@����~��%l�O��'%{Ӿ��!��s�·`,�r�Y���}��\|A@�|��c�M�y�ڮgY�&��M��_�߰�}h�0&��j|D��Vc�*&&(^5i�-]nע�ҭ�$6��(�^)�����Ą���L�Э��C�[����;�Η�dϙiS$�%[9�K�J�~F�L	$"2�tp��H����EZy?$�V݂oa�^9
�� Ix�Z&���T0��� �y�/�x?��p�)�]��.�t�=x��\i��a�YV" O؝�.gf�@��}L�m�9 .�Y�������\����m�Su�J�w��Y�mdm߾/m�/���(l�V`�J�q�^��7C������t��[7�(�f� X>у��^L�E�ɏ����'Ad�>�"���c6��S(wY���&���3Ö���%��M�%������7$|�1$�:1ּ�E
jO#0�����d��rt�P�OS�6od���G��l���d�*2���ZN�-7o�B�N?M���ca�ߵ�2X߯)ǎ�he�����"%}��N�ď�_�d�[�V����z�i{٩h�h�L4eD����m�A�[	���WpQ��XGo`�>89�[�}B�O�H����<��<-���S���b;�}m�=do�Q�����Ef��|�ݔ��Fw˭���&$!A`U]4���$�B�XSOY�"U�o[�%:$�Sa�?�e4�=��BY�Lmh:��
];�?��<8�9���Yj���<G�nG�0���j)ω�A!�beA��x�#���[�ߔP����Y�,e��k"k���f���V�j-|�a&�:ҽ������J�D�����"qP���O�F��"��'���&N�u�0@,��.x�����ƨ�N[9�}���w��p|��|��j;�2�S��?̛|���Y�S�p�]�E%v������.�O�O���ǳ'b��� K��v<1�$D�|�F)�&Q��,\�G����|�{���l,�'{�������d,(��F���3ɓ��6�V�E
*P��R`�w_�]vE:�A�]1i	s��/ar��#{c�����z���fK���D���y@�	�!7T|�H�6�:�"b���t^���0>�,gY_�LnڲI%|Č��������6Y�LR:��Np*Ţ;��I>�l^�A�/���1���N�x��ݣ�K1;����m��{
�H��TĨ���}�,q�W�I �sQ?v��"���v�X�xG�*5E�0�~2?<�ʶ��|��W���CD�/ßu�~�Vs���9~��������7�0���+)�������Dx�W���p���Iy^���:�R����`�r��_R$�#N���-z��ц�H�\k�� Rh)
:	��;^��z2HYHDD�������ES��8���*�笉�k����#tle&Q
�_uA����ٶ:6#�񾇬�w���[AJ��/[@��P9�M󢠱�H�rd)�V� C)J�<�Q"_/�7�̋2^�_%&���\�����ÿ�lv�Jvl�ӑ�L^�;dΪ�[���j�/8���?ޚ��sw �����7h`yG��K}�
�O�����w��RJ��f���̯��hj..�jf�az�TVz>�y��Dgp��F�Z=�զ�0���`�x�?��Z��?�nwS��S�pD��.m,�lzD�\{����פ���&�[Ë8(1ȶKhg�h�����;��ٱ���;P�>w�
��o|�9@����Do����

�rx�E�_8����[�#��8�p*��<�vxb�?w+�(���Z�d�A�X����5���!,aa����HR���2(P�R(f��&�����OO��ݕ�FQ�)�~����\�����'$�q��\Y�
Ȗ�0~\5ͯ�$���u=�ζ��N=l�O�T߿��-��=i����r��%Կ�b�W�҉L�r������+����j�]����E�c�>1D�s�#����E\�yX�&5&����&�m��8,@��K����L���?���+�ڀ��V�GF,[��QADB���z�I̟�}ù^�n�7l)�����ǀ�z����b-90�j�J�jE~�;J�Ff[
�7=�[�H����ރ��9z����Gu�ǭ�~g�p8m� ���]�ё�V�#Q��8�@�Խ�7���.4��O)���?������"��X@�d�%=��D������`��ZwW�V��z(}$��0?\~O�?�|�4l_�3�>��ٜ~����C�Z�؞�d1r����r�Oa�؛��w~�nu` D8����2d��6��L,��~��Kء��Ygfj��'C��_��S�*>�߶������zl���ް\	b�F����.�!w��Ĉ�_��b�}m��2>�~�[dU�j��N/�?��Ό���F�ׇ�.�W�j_��,�.#&�1��]A-�^�u1���MMt�(��B��P�s����@����d��lu�n:6*m������P4��g��7m�X��e;8�b8�?32A�w,r���(ž�����x�|���3D��*6����d��%�*`p$5J�\�vP�;�CZQ��= �=��*+��Rw��� �;���~Lۉ���7�.kZ�YA7�9�A���ͮC�����@9���jU����Υ����f���C}��Ugo0a����ۦE�J{U���mj�V�m�t^U��pp$�ϱd�}���s<��;k�
�A@�\����rr0���
���Ev���b:*��5x�v|��`H�=j���'�!�T��?�R&/2�;��ӻ��\:͠=,!�e�&[!��]��@J�7u��Ɖ	,���]�c��rL4���_��h���x0�EƂ`�~}͈(d��8!4]�T�|���h�'���(+I����/���LU�_"���)�
���=O@Bby�	Y�a�� � MզA�qa1����{~�X�.�9¯�S�6ڤ1���(t����`��D�{����ƧW����)�I�K{��2��Υ�%�'��D�A���fq�cgD���g%����G�:5>�`�T���EdYS�����Wj�� �R�˫�jS�� �s�#��^V9�(thi�(����(FI��~���t[(�f�D-�{�V��Qe6)��>��ih+���\�ww��Z^����d���xߑ��|j����u�����bi�pSf��[���@���el~-�����2�̄\�<��Ie)\ �S8M�WC�fC���;�ĸj��?�����ѱ�����7��	�NE��@��"��y��v�B=�$	���� ��5��{�Kv��c��܄����v4�ߵ�ټ%��P�{���.HR�l cc�C0�]�(6Km������<��Whr�{��%�ۨN[�AEQ�]��e���_�}1i, �������,32=�+l�EOc<����_ڈ6%�H)D�X���A���L��?��w�S`��*�������y����v��0���],�Y�4��y� ��$R��(�������p?-ţ��5xa!2�u�/�*�m��Ve�WO�q��=�6�_�W�^��`�� ��C��_j�� �����7B���������%���2�4��2Ѻ��*e 'J����&�.}%rъ�n�]��>p�B����r��>�Κ�� "��(�|}D����w��������l���?���l�A$�L4`�6� �(���SW�y��^�����R]��ڛN����X�T���/c7����Uܭ���>}~=q��ֶܿ��F�����P��N�W��ҩ#q�*Luq�����[���Z�y�`ǥ����Xo +�ʍ��W���O��qfQ�=\�ˋ\Ә��k�.M��kӇ�=1�@�)�8��E}�o�T�����b�����tN֍����8>d�XrB	�HH�_ 
L\}ٹ�Ae��*�%���	�z�k�_�.D�J����þ�����	�4QA��q�D
�ۥ��F�vϖ��u+
��q?(ö��h�3����ז4��z�F���9����x�|�5O��G�Gz�и�~�����p�*��`�@e��љ4tJA$\ԏ��y�[s�F��G"���~�:j�,�.8G�M�x@�=��y�z��
Ĉǥ��Mf��}2�8.�T�Ӫ�����������t�1֮��G�~�Oond�_�������hd���Eov��E5 �uu�~m��O��;���3&;��Y	����\�{�c�I	]L����%B Ic;��D5�{@�.Y�;�^.��&�b���{���{�Io�px�pK���v�_�R��TUT�'Ar�����q	\�u���J���@OMs���nّn�lX�L���V7��e��`��D�M�G��:(5�t[U흻�gi����W)��%/���m�C��eW=�b/���G�#�B���֥�~��o�ם�~�MR��)��e�y��"����A%�A�<u�)�@��9�t��&{*Zױ{�oC�J���L��"!t��%����9���<��^��L&E%�X����~-��+����4`�WMo�|��śf+�ot�l	8{��F�aVR:�s�#o����?�$��X�7Αh:��@T�gTW���%�0���Q�T�x5��*SMaD�^�'�����[�;�`6�=��^6�mb
�;�;���a"0���/�����5Is9avr��~��6���}6m{-�ݏ����y��@��!�q�s�%a)��kט_/�3�:g_�R܄�[(�t��	�����|��|W�"���}nC�1
�	t��9Lm�q,Kj�Xi���������n��kyO���,�;[���O�.�.и��J?�`�)#{kr���2�� <�o�F�N*�}�c�9�ح�(>#O(�lk�#�n�����*]�ȃ4f[��H��c�"���gR�l���rt�O�R5<L��%Z�Hd��*�����+���o,�e��*[�Ta>�����~�m�ƍ���J9����uC)����Kk
��@�j�e}��?�r��+�-K'���C���h�k^���'�<�u~�(�IZ���n���@} �����C�~#�S���ac��	����&���z7�c��w���WNuՎ9��08��7��{o�U�;�I�0���_��G�<���<�����n�\���B	ԭQ��k���4��,/��w}H���Xۋ��X�� ڝ� �֙U�qq �}�=��`hqê����Վ���7| ���5�v�QB�l�E��ڋ<Uԥ�`D�&	q�˳Hg7h���K����;0�9r����~��Z�:��][�k��Mg��4�o
�)}�q�N[c��޹�D�Qrq�Uӑ�/e`�p��򸈹kޟ�����}$�A�
l?g�h׽S��o��~�t�n�3_H��p��Pq�sl�G��wY�`Cr���+I�p׹��9��-!0,:�j���ci���iq��~u}<�J�n"�:Z�Pt@m�҈i54�NӢ}����+�Ѯb�՟I��5��%6g/�7v�+Bx%){3V$�D.a�~�O�7I��D����Fq(�
�� 
eЍzPyuǣ���29�f��P�J	�� �ܗi�y�۟/r��5�i=Ј��h����� ��P� �X� O���g���c�hLĆd�GB�*�c*�5-U�0�]S�ATdB�U�,����h�v��D��u�/䬺���A�6gw	R�u�3]� x�9��Ad��n?6_�6k��v�wەI���w�#�j�A�~���~��%��՛�!�q����;����'!�_�ܲ�o`���}.�G���tt&���.'���68�6jo!<�2�5>F)
��z[I�]��x�	-��x�jK���"|0�D,?0M~�/��ϙ�5��Z�ۊ!�?o&F�æX�0(��Эo	���ە����X����9(�ȿ�b�G��;(�F��8Uq�#�@֚�E������Rl%��BLlXJ�4�)ġ��T	�]��dL���3FX����MڧKP �Σ�@'��2����@�sKd����܈��egMs�fMJ.^p����ݓ�JE�`hk��we�2�"��*�3�N��/M��R�&����m$x�����<���ʊ��et�������&�#�P�Q?���Ɵ
�y���I\��0n$�첞��s�����ic`ˢ��>s��u�,2.�����b���/(�Σ6��Y�߉�Ui<�k��S�\�Z6�k}n�[,+�x=WL@5��v�(yl���ˏ����[�Tv�Ͱ%٢oѮ��&֮����i���Q1�5�QR[�h��k��ξ�A�>��v���cI��M^U�oGD���4�m�#�*��\�FHQ?�DoJȑ/]�}��������:�f��AC[�q��X߳=+���[��8�����:A�#��iGvMR:D���O]����_*�𑇀�DX�v>~�����VU/ik��v��~b[P����wgf�D����ts&��c�c�+1���r[˰�N��?/�	��k�3)�2�?�M��d�������/�-?�>����Z����#3s���h�#`?o�쑓[?�oc��e�$m{�6�0!��oN�Кs����C��%���0� �ᦜj�wb�!r)&���Č���2ug�J8�wO�#a�X�~YK�1�M�����"��e��çem�MUt����9}g0�&[2��Ԩ��|ܚ��wN�A�����Q=ʳ�NR�.���آC?�I�Dwt�iV�7��cL.���b��z���7'��%V�m-N�oT�,qv�&���[�zL9��K�qsuG�}��\�Gl��ꬓ�m��So�k����M�+6�H"��.���,��$���@�;#d ��5�S�-���:���\����DV|��$JU�3����3X��Ԉ��vw?=��"2{˸�d8�PuM\u��$��ȥ�0ob1��Q�x��Li���ԁ�����i�&B/�}Mmm�ZSz���0⭍���*�r�Ɂ�"���M �����? �Xv6D�o�z�Yo�����TL�#����Y�l0�Z�#��%7�ƫ����͢�8�����7< P��<�?��z�2�,
\H�w�����V:�%�c���>h��T�Z?�tF1)�@�s<���h�ƻN�$�us��ncT��zHo}Pp���D�	�z��������h_�.7��u�/;<�_��Q �Q�^���d]�a���Z���$l�FM(�5���K��-�S������������;����^�0_�6W�����������S������K�f�IԆ�L���ڬ��^Ï�:i΁)NB�tM͘�X�[yQ�0���)���WV�d�8��`L����ȥ�t�c��x��赵~X"3�&�fn��*m��n]L��Ɋ�c�N%�)H�lg�xw��ϖjTe���?�ę�>�wŭ�*B�RyO�X�N�{�3���Q���� �(�+UI����z����vUk�����ؙJf��XO�ƕ��{=�0R@�!��L5�@�M��9��&9{w~����?}�#����8;t�@F�E&�|ּ���K�9<'U�Ci^���/v�OR�vY��@+�N���6<���N�D(�'~#h�k����E�G[�����7pb�����0�����������k��XpZ��L�'�q��
���U|���В�R���b�Y��c�@/�r��'��v��kp$E����dj�5�� ?�2R��dKT�aAG������Sݒ��. >o��Зe�?��9���Y�mۚضm۶m{bg��ض&v2�mk��o?�y����k�u]��꽺��Vi1&��%!�7QT�Ao+\O���/U�z]q�oW��`��ED�S�TWkNa�d�X
YQ��!4�K�m��'A�f���}�!��ĎE���Ʊ��q�2F͵��8�S�����D��@3�y­�h��el�b���萹����0Li����N��P˰��r�$��r��o�/	OKg��1�� �Ѡ��o�j:VX�µ�K��	ξW!�'�7*o68*n6��贮j:Ɏ�N\:��%t�{mC���`7cXa���n�K	=�7�H*�#�"�P�t�֘{��xR�dg_e�i�\̚v��#x/ZO&�#�=I���xZ���V�ߕɶ��|����`2B�ED24}e]��j&)�5�E�I:�	�xj�� �\�����cՓx��j��� �;wҚb%	��yn7i�o7��S�C\�Đ"6'0�6�|��x���M#M�C��c~g�ݐ�W�vS%(b<����]Ep��Ph	wg��0���AZX�3�U{��i;�]���1?�~�םA��Z��A�(�"~�T�n���gʤ0��럎_�I���������X�c��.n���>���\���/�d��x��s5���
��ԛ o��?�7&[$��e��Ms#6�R�����/h	s6$S?��U��Ri*���,Ïp�%-�a=��@O���v�ݾ�@x��]�rbͻx�&�9��_�!��&u�-�40@Y� #��j�e��bP��>��&�b��bAF%��bT>=2���:����	n�$wH��,�ԏ��
d���G�U�މ����݇�!�%R��ˆw���槷
:
E�|�}��H�F��\ x~pdO!lCwn{b��g6#������J�(�-N���.�-A_��}f�'W�K�7uB�s��e�����Z s���5I�`7Y1ں����0�Ըct��s�|N��}�2��$S6�d���߿����k'����vR廞\�I��r�}��7�O� t���������A���鋚�`
�z����4J��q]�n�)7dTE��9�s¯�A�E��\������%h�6 �?�?~^���&��ėIWGy�(�q�����c�L������;�o�R���ڈc���J]�/!��$�F��z�z�~���l��i:��$m��3:N3��-�!?�����X�6V�u L_�X�e;������1�_�M�n��#�P[O#���R�9��]iЂ'���zx)���ћ`�+�����#���'���DM,��x7u�ې:7���~Ժ� ����Y���Y�]�ޔ?����YrX��$M���F�P̭���!��-	|���E��� �I���kcq?!�1v{WA��pI���+$w�Ң�Ug1�&���g��?��Zu��/	����<��x�w��l�W��Q/X*�>�R����??FV<�B�1�jA `� �z�k���GV�TBKR��Ō����{T�'�ڏH%���,G�	f{j��%F�����t������_�'�4���n�i�< �Z������Hy4��c� )&�,`ʡ�����q�l�E/�PEa@A�K�z�Lv����<�I�%!T��~��^G�gG��;�J�A䐣�\-Q�=X]�D��L N`��Y^�J';y�+�������J��s�kh;ke�Q��Ş�͆������Eߚ����s̜�莲^�:��vWvWBXu��_��z����<���]��.�*�\ږy$y���(h�H�qb�(�c��ƹ�c<�� ����>�'#|W2�A0KZl�;2�8l7(E@S�	>T��uSm���& փy5R{
�%d���<N�ɑ�!z}�]%��q
kf��C|�Ą@�! �4>��E�e��DBCUw�o���1lK��oZ�{��
V�ޚ���4�ط�0S�k'9K�B���O����)��������o�w�$��L=`�E|Bkā�F�0�AL���rh	��xI�GT��r���p��W���p%?�k��PU�B����M���ӌX
��6#(��(���l��+�L�K�v�0��^r#@V��J2S&�(O�9'��(���4~��{yχ�4?�
�z|7̓���>�4�:Iֱ	Ĝ�ӷ��v�H��]v6J<)}C���oH�!�~�0���o��!l�ԑ�|;i�mI�c�F�I9S�K�����6��йq�љ�)��љ�\l G+��-:��7_xk�� \�q���)�Zbұ�N�Ҡ��9J{kpy@ 3�0���~�S�\?�# t3�jb���k+��脛�=�.�/9�,�5�a8�,�@�UR4��8o�֔��+��[�z�HhR�5S��9,�#{ ��DڸFQ4�Lk�-����<؅��Ǎ�D_}V�>��f1�!��P�+A�}���9j��{^o��V������#�c��5ˬ��dG&�A@[���Ȥ��P�wn�B�$����w��"�6e�Iy�"�.���~a����"ZiM��N:t��8�F��l`C.l��t��`�n���ֻdfV��y����#�
=&b���&�L��>t�	qi�'���Q�=���G���ke{�V��e�M�%�����b� z�>�?�D��;bfOR>��G�^��g����F�؟��#
0��A `Q0Aڍ�]�����I������fe&�Kr�U*x5}�75���x��T����6(�D�PW<�2�Bx��7��8tntu�l������BA�D�K����s��*�,�wg�����®��L"��gLs@��*iWctIՍ��`[��ѕ�߱6�fm@p����3�X\R�����,�'ux�X$Ԩ�̟k>b�֭�������f-��&�W�EZմ	|9�����juM'3��}q�Y��r�q�MG��U��k�ub��C����1�Q"06M�*�<��۶�U�wL̴C��qͿ��\,��\b�"]�}���k������h���$BA�
cg�	��e;V�Ad谻iF�y�{��(��m| ���*�"Ñ�|��)�!Q�������)���f24>=L�� 8���k���V�d}<��]}V��eD�S��/����`h8�b�D��Ƈ�����Cʒ�Ɉ��T�s!c�qvQ�y}�sJR��L]y(�/�l2:pǽ�JNf''�m�^�E ��hD�y)��/���]�B@�	d|�41c�Gv~B(�Ƞ-9�ر�».��VЌ�� �o��#R0k����Wǣڝo�ˎ�H��T#8�l�ӳ��ZB!x�����8��8�?��W�7�
�!JD��v��.�D--�V��	�b�a),��FP�l�Ƈ1V,�w���*0�Q"�$0��G��ۊ�.dSM��`������P�U�68��9�Q�7) �W9d��Ky#���{���?|�	�~���{��W��a#��?�]��/��T�����쀒�Q�8+}�#��j�`�<L�ro�Q��@ '
Oĉn,:ɍ��SH�F�h�w%aѤlѧc=[u��ϐ�Ĳ�e�Ze?�u�A|5٘m���`e���G�g� B(�t(��[N��ʀ����y���gfc,���I2(�������θI�"��QG� �eq�~�JȂ���P��1�9qh��߰��`�nxˮ�w-�(��#h��wwg�$A?}A+W�q��B�M��A��Wih��m�6��Z-���ԛH��T�}#�=3Y�$q�a[ͨ��q�R����R�-�ϗ�`d9� @?�^�hkJ%`:�X"���z?���l���)Ò��x�7<������R}���Y,�TB�Q3�����A�wwe�=������ʁ1<�Z8|�:+R�%4T�����6=H?��g�*��b����ZJru 8v���Ǎ������A� ��g�M!s<f̵ߚ����g�K�f���b���i�,�
;vZғ5�*C
�`}�<k���k�{�ب�^ ����\$�6�Û# �Ѵf��!�l�2�F�л�q�Y!�\��$���V(�p��yі&�Y!����,H��-(���M p%3����٣?��Hz�C���ʰQf�����ϫ�SvM��D��33c�ڹQ�LǦLX�@��������8U�W<4��4H��֏P�b�m%~�C��Sѷ=��B$�y3���/�R�yf�>�w:n�Xh����(B���A�@Q��YX� ��M������3�b��y��>&�ڸa�GG�Ŧ�����P��X��e6	�o��w�"�g�H�Ȗ\-���伎�g��,�ݿF ��7�D�7E!�F��/�?��@*�HO㑑+Dk��)�_�gt@N�qЋ<=e�	]ؓi��k`nux{�7��z��,��F�����yX�@\� ��R�l�G�Dt
���z4F���y$��Cm(_Aዳ��J�O���Q� �2|A�͟�H}?��V�ax0���TX���Ѿ"�I3zP��oف�z�a=b�_������&�>W��:ү:r��s����"���	�E%]qgn^��ד�3��[S	� ^�d���7�����!�1�a�qo&�Jw������X�j�>ߎK�>>j�/�^5��:M6K���1����`��vN����{�LiQ�+�NaI{R�����":ڌ"����I�x�2}��{L0^������@S�W���3ڸ jy�w����n�������w'ӻ�6f�;�<��\f�g^z����v2ʖ�QT��>�X��v/C�����L������I�U��y)�E�Ǌ	����_��^���`^ ܁w`T�~?+6Z��ȚNM�QZND\ک	�"m�Sh�4����c��+��
ا�D��F��]�����UW���;h�g���^Zߐ�5�IͻH#�̻��x���~WJU��hU����*a�O1�%ʊHW�>�I��aͩ�� ܙ>9�1�9����]��K�F�⚗�K���'-2�Nb�(J����?�������~U�2F2Ԁ�X\� �r-�~-�j5�[����C�_�U��y�B�c�#Ţ��ќC.�ܣ!�]�n>��b�}4��>����)����K+l8m�M(�=������=�;�^�	��^�(F�Ð���5��muˑ�ٱ�#t�S��������۲|6^���{�8�(+ڀm��[�Kf���I�f��L��Ĩu�7���?�?k��-V<�)8y%�Hӣ��:�}�,��}$��N�+p�̚�w�1)�Gnr|����(9�(p��T��g�;�%�	���u�8~�5Bfc�¨��:*
=s�$���g�TW���C10�K<>7�O&���I��/�z�#�- ��v�`.��x�8�%^��-��Ğ�fR���F�V`D��p�0��f:�[�8+�Tі�,z�ٍ�gT�xV��4Ÿe�-#=]S��s&���6[��4�����o�	ڞ��{���+�&"�[9�Y9��B�v��l������8��I������߆MxzӲ�~�����U(�6ma���}:b�Y��|����E�:]����/�~6�U��Y�6K�z,�ӟ�/��Ԋ,sˊ�9|iWw�j�1����=����g�F�ׁ^y�F�V ����J��tb�8��)%T��J*;b�.�j+��}lp48Na}�Uل{��#��o2��%����lȽk�]{���!���u{b+��J{�<>c�;��`�r�Je���>��V�c2�'+*�Z�O��f��HE�%jp��kF�-���6�ͩ-9�as�w�8�g��V���T^�NYG�Sa���iMo���F��_DC5�ER��YhF�S|������t�?z�(����ξ<n�Qz^]�����t���[C��G��, k[���re�,,����"���Fs��Ж�(���#�s_|B���z�5�K������0���@򪝧/)Cx�p�<wj��g�Ҟ��4�H����������|�ї��������*'� JL�E����)����O�v������a���=�����Ho�Q��1fI#�g���Wf?��?k�SB��sv.�U�0Κn�u�����A��g�କ�W��µ�+'|j��
:�� /�{�*Լ�1�e�j�_�o~~(��X/��{֒E}���	��miWpC�ʓl�\<R���d�n]xa抛?�D��/V㋄Â�t�M�X��-��D���8�-:�l3�/�݋�ϖ��u�N����v���e��EB��ySa�y(f�^ޞ�@z���{wO�zȼ.���wŶ]D�D��2�$~�)�?K�gZ;$�\��� ��/���˟_���;K�;'�s���,���
|3�)��]68��<��d�7��[��?S�u��,���ʷ��z��&~�B�'o�@�~�p��h��[�rZ�eaCj���>�>D3r@���	v�q��6o	JCDӽ�FG�S��:��-(�l9ai����A��2�+�Q������]0��ţA�A�:��唙� 0�@�ϼ3��1Ơ���VP��g�R"](\��$DIfMk��L}j���$p��2�σ��i��`w��w��}SĬ��:2}��3F�0X�}5 l�(����D�<�X�~~6�l	]���Iβ4��t5y�"4���%��NE������Iԕ�=/ؼ�������X�����u�Ñba�~�#�a��X�~|)K�G�W��+JBc��s�����J�f�{=(�����͑�� *q��!w���.â��\ZY��+mG���=V��}Cu�����o�G"!��RS����2�U��-����F����[�N�w�J����U��$!	oo�d�����kiBu�UƷ�0m��-�>�Bl�I��<_ʅ_O5ͽ-Q�[we��xW~��^�7=�N$�w�|�6̼�!(�U��Li-�r��J8��|T�M de��g�|l�_��N���^cfI��b��,v�a�\o��b���W��7B�-ZM�#��_5��Ӄ��?�R�aI3����/,�lb��:�N<p����"��
���Nĸ''�Rh�'o.��,s����&b���3Ҡ�E��G�������8���7�}���qv��q��Z����k���Tْ_v�B��<,��p>c@���3�̰)B�U΃`�"u�M���e�����N������ng	X�`r��R�
z�8��c��[��	W��,�7��{�o4���&����4�g��8���p�B�<�������YO@(5��7I9�-��\���j^���3� e�'*C,��3vX1���8` �U�8�)t��g��1�T���(��L�1^8����8�k͏^}^=��_�Z�6H��u�	oh���<�J�%��`˫>�����8,������޺�4:�#�x6�b��P�� ��t�}�}I���6��N,(�O?�Qx�Y�ힳl*�d��4��d�t;�J���{\����O��G�'ܺ��\9n鳦w���E؁wo��^�B^^ދ��u�ՇO�����.�i-�B/	5ԤGS�`eS7;_����^Y`h���c���v��)�t,�WGg5G	�o(+�Nt	����q`nC�_�L�Wf_��қSPM Rh�?b}1`�s8shA��2�G���3�f����j?!��Wmw�Ig �O:��b'7:m��"�Y�o]�hS��a;���x��*�j� @@��6P��}7�jn�4w�zv���H3��	���I�YcG�vuT0j���k��e/L��1���i����J�`�� ;����C�k^�݋C����|OX��uhvI����L3V����p��5���	�xل(r���]m��u��N���5�>H\�}��҇��+x']�U7��N��!K�;��3�v�4�\:�_E��|��]�B���2s?.6�!�� G���^��F���cg���.m��e�3���i����"}�T�Dm0�BȜ��mV�<V���cE���KTO;?'N ����+0�
�3��?Q� /.մT%&�R�V�ӴJ���J%�//���xǻ��WQ7R-񣇛1@��5�N.d��e-�ٹ���N����m.��{X�|�G�%L��N"P��VR�{�}�̠v�Ȃ|i�c��J�ܹ�m�I���w�2,9��*���Ih��(��������������N��h�D����M�[tU4<T����/:!6�-�'�Xٌ���j�~`RW\ɾ�.�{4i�󔀫 �԰V�gI����0�A��*�7�$We�z�Ǒ/JWNG�'T����a顋�uY���ؕq���"x���_Ϟ�gy_�nsTK;��/t�J݊�ĥ,Ol��P��9�����h��Td��v��SIG��u�^��,G%(lE��*'D_��Zr�~f:E��H3�<m���ٝEԅ&'�B��lD��i<)񔖞�z)�N>O
���'�~�����n���:�}��@l^a��yYFo-""	~a�[W�<2//p�|b�����l2i���Qo�sڙXj#dXN�J���3��w�DP�@kLA~���!o+[�3�$�LV40��'R_Wx 􉋿 5r��B#�����g�g13J�K600Z(���Y�6�	MSS��r�%%�T�"aN��R4zG`cf@�W��ٲ�n�2����X�+�ë��To���M���5*6.	�m�{ۦo%�;��m���@���Z#���	��!9N�ܟ?�fB��';q63�~��=�y��o. ���H q��;�x�&݆h�b:���q�۴��������U��d�XO�d�jB�dy�TW������!�]姺s���X��-�\�ᢌn8��s�(�3e���;�=&'�M��6,^�����Ĉ4m(~�(��S���h3����O}B���Vطy9?�8{���zd��������̝�iW����#������D�{9'�d��_ִ?����>�=V&��M���0���j�:����t��͂��~�ÙɅ��W_*R���VY�<Ϻ�gj[�z���K�L��������^L�<����M��Za*V�	,=<V�������G73/����u������Y�<O ���
,7��_pCa�,C4=����[�S/�����R�b6�����k��e����59ф[�.B~��mnn��(�N�Vh�K�Z+��k�͟�7�<��(���A�t����?o�b��2�t�u��S���F���A����F6����QyS"4��
��Z���C����,�%�yt��p��l�l̆�߀��Gm?�L�|��\�~�Y}}/����awW<�"��n�x���~"��҄u����*��.��}�vۜ�a ~��;����Ca����T/�A+;���	Eg�R��df*՞|�m�mu]~��AC
+Y\?ti2��{�ґ��k�.b
Mհ����Qccu5Ь�k��aً���1I���ٍ�p1?�����OpIh�'l�l]�uv��"�#��E���$���v��tX�q��b%DV~�y c;�Q�2��`$$,��kBj�]��:�U)���uvی�z�3)�_]�\�X���ţsVw�~=7�au����Iu~1k��i7Ǥ?@t�mm\D�6�2"��u+�����H�����f�Ӈ����ޞ��ֲ�o{7p��{{T:�M��s��A�'3Y��EB�Ϳ1g�vki��f�G�)�Oz_q�S��fڐ�4?��Mb����o!è�����=hDn�.����"~����y����l�����|���hf��L�#��>��:�TZL.Bo���r���l�'�k��hMݼb�����M ��@˵�s���}�%D�} �Y��}� �'��CV4N�-��آ0*�إ/z��(��4�GyE@|�������d[��84%6���..�'%�p��G�����^PW ٞ�w�(l���1�r��յp�I�S5��►zP/�TK;b>�+��ֆ?�ѿ?���!�݆�T�ʂ�PLU����=��c�M�0C�Y�����E�K{ 6��j�^V���|�̞��,��(�gY���G����d����OH{1}uagv8|���M2��(5i2Ƀ֝I����'��/++Q}���Z�cdl*�"�KQv}ÅS�5T�SH�*$\_׷�bh�\�96�\�oD�Bü�;�\M-G�� )¶���D",��pߍU����քa�$d��E+j(��٫������Ķ �C~��?^휀���������|��9p����6�����Hx�����a먩hD0}:�� 9�����J����N�z�'u��˷󝦯ޤ?�[|��a�U�5NA����G�*�:A��F�����B[��J�u��ȸ+��։���\�9b����xQK#jK1��Sy��L
�C[+? 1Sͅ�[�v窣�YWMBp�m<���Ш�X���-��W
�O�zO�@�猂>\�se����\V�.� ʿS?��q�ع�o�	�
0��yU} 7�5syIiK=DrH�Z[-!6U�x$Ο�����;��/�� ��I����Jb�`%��[ל{�Z�Y�\���`q�PO]8�ѝxI�����2�OB��~в�JCbe"J�J��=tG��2$��w?���F�J��c�q�������/���B��8!@��VAD��T,P�O�@�z_-��$j�N�����*��5������.��}y�^�������*-�Pz%ӥ%�~�:�n�^�! y�Sr�M��t}��Y��������� Z���Y��.�	W��V��Q���u��i�͒Er;����u����U}��42��1BI�Z���(�ߞ�SFo$��}���yy~�W=]�ˡ��j�U���*���t�KHHHɉ5����=�c�fU���iSnf���ǫ��@%O��u��ΰx5c=���Ƅ}�^'>�]���kC�8��sZ�R�l���ڕ���(`
rwj�Z��!6bc�M��~����dG4PLg����3���؝�v�	8u�4[s �����ʹ��TT�%$Bs6���[{�
"Ge�\,ij�sk��R70��Q��
����R%.%���N��㐫&��$�oK�����eC5�7��O17q��x`�y�ҝ��W��I�Q�d�$	��Mt���_�� �uZY[t[	1�9�y�^��r����N,�e�ن��	E?|ۯ������E�{e��a�+8�#]�W����Ɨ�?�^�3�)���h�i�ߔ�����bE��]�R����b��1IA�M5��S]3��c���6�咽��#�E���mm�(xg���a�a�U	��9
�\r�3��ޖ�����8)#�mwPx)2����Ԙ�5�U���Q�%͕�@4٪��������|^���įx��܊'��*U�|d���A¨��/� �-}�z��n����U�}R�݂<'��o�>�t�f��5̽�����[��|i���*�n@�Òb��F�̾ѽapyDQ�����̇�}2P�Z���N3�红6r3�vқOc���l�N�w�d��n��<�}o,�*h�W���Uc�Щ����{�9�ͪ�F��^�<	�&�8L����5z���$��g�8EJ/��x�A���&��y��Ϧ�>Q����"���;�P���1�������a���ȵ�� ˋ����-�.H�v&ShO�[��~����gٲ���&�奁Z�D¾��y�;��0����=7�&����bL3�M�D�g���Ű?��n�Ĥ�a��b�a"5U�@��Ba<��`�����a��0�۷�4l-K6Y�D�`+���B���q�X�Ţ�^/O�A{3I�N����̼�?q-�E@"{�y~���L�l�.לi�>\���*��@����n�_1^�B��M���x�N+/rqVW���N�m���@�و^W a%ԥ"����,�Ʊ|}1;�y��6��ǃ1�x.��ҋ�=t���8��/O3��8�R�����K�|�	��4�e��18jq;Z������7�o�����ev2Ar�ۏ#M3ɩHA�%*�V耰\�;!9�t�ϳ���gqR��2l��|e}r��X���Y	snv��6���r�CVz�E�N|?	rY	3�)CU��	˩���⩉��3��mEa��-zBk�ʰ�9�8�@��i=�Wzq�:焘v �}q�sޓ�K0����pV�����"�B�[����[8i29���h< �,(���zY��9m��w��7%�����wGdƙ���S��U�A�Lxۃ!t�_�����%��/��nv�6��/s�%)u�W�ٓ=�Zp�ºwS�[�M��<��u��e@c{��P�����ڎ}�7$����AjN֩Z�t��0��T���@�����U�$*�t ��e�����D�MNVgH�1^Vd��e�q���!��=Xe%��[��[a��HCy9&��x"sl�ݲ �B�!�%�d�T�*����-@l��Ya����Ů$�.���I�.���S���ol��7;a�E6n���I����1�Lǂm�o�f@���6�$~��h���N�"n4s!�O�$_�
�#ͨ����H%����2�~��@x��7}JE���`����Wm��#e��/�;x��ml��c0�.�CГ|���X	ܺ��'���
y㜉�=ϱ �8��̘B/A�_��'��XT��J�2�&��S\,�B�ۗ����2��&Ò��B_�/��u���{�,���w�ي��C�Swkzi��mw�e)3~�g�e�*�������I�â�3zq	Y�`�q�Ͻ\<�C���_v��X�:N�?tY�ե���`��A�Mǚ6�
���g��x��`LT5N��3���y����=���2<��!�����V�l�d�yʂnЌ��$�U��
��t�H�$uLr*�}�A׮n������d�t[_��� �� �䬭�N^+������i���,.mg��ʨl	|�S�`ȨQA}��R�L����u�z��b�PI�ƞ��D@B�[U�i󉾈m��Nm����t�
'�3SM�n�q��α�xA	Z�x7�ک����'4����+1��1�>��U���`+��1V�����G�����eE\��7?��lt�(d�k��T�IC�fJf��s������2|̋�o�b+,Ԋ2,k�n���O�U1(��VmL[k�l\n~Tb���_�QR��F��5�	����6>啔U�Z�0{-5)���%��Z�c_��y4��/�~;�l�Z���ռz�_Z㢃��ű����L@�a�+Dh��H��@s=Y�o�'�݉��MA6�h#�{��+�4�n�QYٽ�7��P��d��\U�>��Ʋ0�w<|�k��ӱ-��n$J����)$W� ��j�	�
�n>w��\q
޺�k[a6��=�@6�aUM5����� ;/��ץ�j��恨?�Y�o�\���71%��+X�td��<yf)S��Z�2�{�u%;O���e, gRR�-�
M;+P���XcG�ԫ �rq�+	F��g���G�;c��G��Wܩ�6�:����d�1�堖��ҫr��v�A�,�oWV,��J�]	������.���x��/UK-r�|Y	-��D��Kc*J�˾�{���c7�WZ|o`VH��ӾB�m�g����24���H���3�c%m�~Ko�8Mlv���\*�/���\����S����$%�sb�Η�g��W���0���w�ͥIf}����}=�턞J\����1�ԩS����데y/��� �vm\�aR�����vj����aj�Zd�CQW�.��+ ��MW� �����z�tx�&��fit�����/��58��'�r��&�0�t��O9��ϳN�-��痺����j�y�*�8Ŀ.j����Y�U�����ٗ����l�j�e�4��|�hg��.'��G�\����g- �9+{�'m�k
�����9xl]?���Lr~�/�6�̯
�ى�O*�:78���ݤ������M~<y�0�4Tԝ��޻��+X��h,�}�J���!|�Z����n�l8�cLiL�4��7\}��}m�%��*�vl���[��

�����4X�U\�:��E�˜���/�u4��Xߟ����n
��Ϟ���82v��K�{�|uG��������Ō�L� o�7�i�_�~/w]/3φ�����ޏ�|�ľ�v�w\*�gL�ϗ'E�,�q��V�%0��r�Jc"��@-NP���kG�����/8 "�R_n/�/��l��Lî?����{�W�[��/����Ld����J�۬�=Y�6G�x�x]��
��4x�������ʡ��@歵����ز�0�9��N�qcüo��@�]P2<7�7+,S:(IVS<���RӋ֓p�{�H��F���͞�2���呀'1c��@5ak[nm;����g`�Q*�+X�K����tB�~b9�� ���g x�|;x���'��ηI�ڲ���Хl��'��$�|'�,������F].�N7Լ��ɴԮ���=�f�&��G<0`�4�?&ry��_#/p�
�@!��4UTu�7Чէ���1�𸤇3}��Zo�0��{(6߿��"���'��������e�W秛��J=/SI%-]��5?k��W���n��Y�]`�̉��9��y�ˎ ߷g���7C6�R�z�Y��񝇷\��/���)7����%��s�/�:�� I)�GÌ'�Ԡ�dr�a��#B���������n�}�g�ֶ��<y��������?V��_�E��B�����Jg�1�A����7�@z��3��,xt����U�R�p����T�&��Tf��`�>^�y��
�߰^nb4�� )�}Y��H�r��_w�z�&�ecw<�fZ3tV��ٯ���Yti�gS�b��l+�/�f|�ي���x����`+A_N�c�˙��2�O��+ /���ewlQHmB���z!�nn��#odC��a������?�,U]N�K�j�,���)���k�y��<;���28;�R;ɟ_�~)^��h^���h��*5^2�X��^��2��Z���B�N�j���f���'.<���h����F�	M�'��������v��p����A:��ӄ�Β��(}p*�5���$�Ű>���������Q8��ʥߕ�����(�A(��C2
2�f���Z������<����0�����S�(������4����N��r���f�h�^��$�E8���e��)��U�����E�n����R	�\�p��Bn�Q�B��.>�����_�ܱ]�_�k��K�Ψ���k���Fm4���N u̹A�c̱��yg�$� `Q=�+�G#bc�!����]�!	���ԭ���ftU�����qt��/r�V*�1���M�i���:����T5�:-��	�x�-�lFTф�f*����Ϋ�֪rU��&]����TK���̝x�z'Hp�^��t�JÐ�/Y�Qx6��b�W�VR�ۊ�
F׌��i+Lg.<���'`�^xSu�(
����geCa���z��`}y?
�����=MD���>�R�*�G:3k̀�i������-=\㸢�NZ.��+���"��t�^�X���y�p�y}aR��d�]s�>��"��]-rB���DwP��K�S��#B�ys���+Y���4�FU���v:f;QO�,�<��:,���Ձ	G���H���\R� �t�"�.�s��_���爭)w� .��J֯�ʥ*�th�ن?�-+��o��s�9k$0�n��t���+�T����p|�oN�W�ø��#V�0d6���#u{�q��צ��I���$�K{�=^E4�[��͸��Q�'����w�N�! vN]L�(G��jb
+VB���B����O�Dl�/YY�wZ#g?���h|����5��G��Y��n�� �轟sJ1é}.�C���ϻA� �%���bf�]C���I^l)+	�v@��k�����{Ű''�ﮫ�c��딉��Ϧ�UJP�ǻ�o5�Z+���T�����\��I8z#�۠����I����)�_�EFQ:/���Lu?W��Ͻ&yy�T}�c��eVg-\��"DR�j:f>.��;���V�v�������|f�ud��v�o��a~���Fr�������?U�(��6O���#�����g��S�Z� 7���p���ۋjYp��b�TdgBe�gsÊOx��dOk��� 8���eUh[���w��VN��Yk�R�����̴`�JOL8�75�W�L�eT[����и���;$������-���;w���:�������?���v�=׷���m�1ݾ��I��� �t�zoi�梹xs�|Y1����@��x�|-L��ɸ��x���2W���ȯ�xX�*��R�I���]A9��շ޷�jq0F��V�j[���{Vr��[�1v�d�Y��6 �
��:��5�a�QVDA�������������Py��JW����{��Q��>�=6�-��F��阩�c���]��kP�M!�h׭�ʜA�!�����^�S�%��Mx
&�*f�r�4p�d�կFfAS�P�J�S(���p��|Q�gQ��5���F��}~-k�ϫ���E���^ �k̖��A��m��'_�'��7��]��dߓJ��/=v�p�9o�[������h~����e۩u��>ב)�گ��v~Z���~_$����{ӳ�s@��]w����>���+�)���3��?���2�Frd>�y컙zM�2>f��.?1b�����$I�:�����RA��z Qdt�)E�{��Ğ穳}�\r�f*lQ|,kO`�7t�b�;�"�K���h)[6�&vP��̭�HZj��|Ŏ$cIް�~ �U��l"-���q�<\cՁ:~Ю8n�a���W^���z�|l�'�˱�/#�mp����}:#D�k*��l�j�c-"{ &D��.�C���%�'?�����	�:j�Ͼ�:a�L�.fOܱ�|Y|��H��[-�A�|�@Y�i% �W�M ���>+��\{�u/�Mq?hB��4��ؐ��?U�R�b)x#��`�3[Tմ��ؼe�����9��0E�g��n�jq�Nzymkf�ێ1����Nw��e;���f
�SL�T��+Ļ>��X������jSץNL��GA��$�;�w�/'`��i;�&6�����G]����!��k.�^�ٔ_V��yR���~Ua�w{���1����1A�*mF��ǣ�Q���n=!��k������D��Kŗ�����ޯ­��o擼6}Ύ��l���>�*��կ:�T�\�l@�kH���h<Imq�ԡ�7c�Ǿg��e��ja,����Q��>������=�2N�$�������Nx�RR�A��Z;޳�p{��:���l�6���z9{�ǧ��� ��J��	�脸ۏݽ1�/^��U���Hk�NE�V��lZ�ZU���b�s��}"��+|׺m��"�Ҷ�&;������b%e�n!N�?�O�?�(U�w�ٟX��3��y���8t.�)��	�G��"hӓj�Ӟj�N�o+��\[tN��X�<}�>s��ڎ�p�i�п)��_��su�	��obD>]�2Ny4c���l}�a�wR�b�o���-1�+\D���l��S��ZFGh�	�/��#� �b��S6a׸c-tnIdGO�X��k����폿[A�8�M܁*���/;Pը&GHj��ͽ��\3�頬����B�p�'&A�3�K�T/��f�Ƹ����l�!j�N���=�"*�?x)�ٝa���՝�R�+�gbj]�Х�gq݁���KM�eE���Ò���X�2]J� �Bx�K'yi�;rҬ�{h`Ғm���A�U�>M � ��n��GRڌф�խS�u�������a��,�����Gۙc������:�R�"��d�-��E��TL�'�̂wb��m��IOm�!L��x�����9�Qۼ2����,�����L����k�D�kr�z�;k�1��rZ�Bzf�Mx���~Z�Z+���j�/��7_YB�Bw�u�~P+���cߧ�� �����X�!�n[�?j��?�`�lс[�Q�!�ַ��ok)>�/me���2�Ϊ^��[���4�o��(����ǷGI�?��97p��Td�	!7H>j��BO��d�!�	!S�2��������J����:\|K=�1g���chK"���?&�=�}��ɚ�'�2+\nXi֜���ًA
�i*3Not�@yφK�a��>d�nAF���6a�26��紷G��KBv6����;. >]�UpP���Bp���0���ɿ�1&�d�Jhʫ�z#dq���9��|�E5pIyU�Y�8i��k˛a9e=�P��ܰ0�6\�`�ظ��i��m�d5�60Kp�PCK�[��i�ͪ����^=͞���[)j\Q��k>Y1���?�څZ|�g���q��r�U{�)!!݁�<��8@d��,��Q��A�Ҽ�p�#��� ��w�Z�݇>z�Yߙˡj�GKJ&�3Ȓ�`�fV�;�I�jh8�NV,ץ5i{bqͅ$g�*+!�ڜ�XpV��2�+�q�k	+|@d�.�C�?L��[�
��L��5%$��OU�r��:��P��F���Y�ˤ_\�=��w__#:���D:X4���(����tF�OTT�f����#EEYk�IU���ɲ_��Eо��N�γ4����;\��>�y�s�7�ԭTx���:��k>�c~d��D|�̖�[���~����g�%���㻥�ݬ�_��E�|~��zP����o˲�����].3}����q7M�����yD���U�h	=T:��E�L��1��_^_�I��*�q�Ơ V�V�I�)���9��(3i��͝	�����b�Z̅�'\��9���/9�S�������B��<F��lN�{G��̫�藽K�f<��G������"�k
����y\ü��ᄛ�x2�@������ц��|+t�A�D�.z�~[G�b�s��=S3�Д*�k���^�э���c�yL1��e�!'�7�ըm�h���a�߹����¦)���a�y��P���ب��,[��z�-V�otE��!��M���9�����7Vac7p�% C�<o�OA'k��cQ�CH��a�/3�(��e?]R��A�K�m�"߉��G���5���zo$��9�#n���6�J��a����$��-ؘ.8�;o ��sN��&�$n��>�;� U^N��i�;á2��o׻�Y�l�i��e��w.T����xMs��	^�A��U�}R�YŰ*�3Hh���]Ml���?n�E����o��$�齐7��O�[fo�I�@�~�X�\x�@మ��a��@h"~Z�5�c�C�T-�z;����䉸��2�j62>�a�;]m-��Y*����o�k����1�H� N�w�e?���t9��_-�Tƻ?�L5�)>��S�C^h>w�Tw�yw=o;���.ύ�����7�T�����6�}�?�8ݭ��Kiy��/ׯ�<\l�c�ۊ��D�֧����c��p?�Ǿ�ې�5*Me�rYC��=a^u9'F7�"O #�8|9�u��kk�hӇTsn8��D)�Q89L��U��#z\�$�R�g� �F���s��jO��?/���@�i%��6�A:�9=Nm�~u]x���zS|zo8F�[ka�l���������Mp{C��C�㰴��kk���������&����S�~�,��`�������r�$�ڲ�<t��f/��q��s�1�S;j�Ϋ�5I���
:�I��ڕ�}�8��$��p3 x���1%Ԙ���~׃�['�V�����1���9j�O9@b�o������eRRe7��.�A6y@�1+�
���AI��e��D�UWC���sb�q^�������R:���o��l��\�='NJ�>��6}�a�ٹ�z;p������lϢ�G�v)I;�,��*GX�IS�"tH�s˟Y�����.tA�]�o��k䂏)uk�oח�Q��{�ۖQ����AM)�"����Z����@7�S���yK�,�:6�~���N�ن�*Xڥą��q"/0�,K�����Y���K�T�*���޾���/��#����9��# �;<� �cOzj��8�q�e�, ��D--�f��ާ$��>��x��s�[��j��,���Z?+u��������UeU�睎|K<Z��^&/���"#�i���n1���Ԏ������"�Kg]�L��;i���~��L��:_d�l���'e՛;�]�k�Q�*\�l@ӱ��ߦ�����2|���|%�ґ�(�yHb3:���pF��0��1d���XZ����+�cC���4.���-�~87 ���)�=�Dڇ�yr�Tp\�_��@�5^B�)��h����*�W�n������Q���H�Ѐ�U�����r)#�N��B�� ;mV�ff}7��X��ǌd���7�C��D���N�a���3
��TS�6�T�-�xE�����-������?%M��W�}n�����q�?��{�É�]���w$�aSH�����i�6l���H=����u��|{.��/�U֚�T������ve���7��F`��e�Ѿf��ǎx��%�n��L)�H�f3x�*��M(�Q{��0P�=͎ۂ0��=5�r4������ܾD��7�]{�u��#�+����H���n6Ჲ��ETq}�����Φ�dvlTB��qN"���	vS�ۇ}�k
���}�>����i���ȸ u}y� ��4����u��⛢��̢�*1�]\B�p"3�5,�ϴ���,+�������r��u��Z�nń R��\Ѵ��Iބ�Ĉ�"w�pu�l���1��{�/u��-�P�C���R�$|(�3�7H�B�(m��Ą�1d��񙬕����/�/���ti��ȄzPVq�Ӟk�f�2�ڱ#��kF���ta�sV:�V�	��9"�Z=Fh;d�c�89-��7���M��R�xv\wO�+�������!�Z��c�-_���������+��d�m���<8��u��j��������U�̦�����y�2DR��Vt�����m�I�&[P�?�t�z*Hg㝊��Jk<��T�ԍ��p�#�����`���zO�n�);6o�[� s9O�9�g#YHXF@�U��k�}����K��M�P�\x�̪�ӏ���������^4���O�L�3I۵@c?��:/ "MQ��eiSh��q�b3��r�yˊ�EC$�|��Zy36E��-Y��Q�0���z W���&k��?˖����ɸ���O}<|�Y� �?U�ݘ�xb���P,���
�0�!RT�tzlB��~O�2z\F\�sT�����(.OlD��Q�V�¹���n�=i����Y�D����܁�t��t���$��Sv�z����I�Jm�U\@��Ǡa��rzl�@SZ}Au	1�c3ԇ�A�Y��8���Q@�Di�4Z sN��2��U��Q��dB�gƲ�i��nEI���U�1e!C�]�$Ń��IM�͢���!�)����5�����*�QƐ��s<_�qn�u�2��^���4T���AF�O&�s��e,SkJ 3��6˻M�Y�ǽ���iq�������W�T_�?n�Mr�-\Xo�}bq�+1XJ�$9oX�2!5/�(ɥ��s=l�x��)LE;��.�p�Ͻ�z��,��V�Y�}�o��G0�B;����_7�`�-9�ʍ�^�m��m8��6�c�3Cȕ.[i?�-	�d�R!����� �XX���� �2{ㅮ��m��K�sAy�[��NUv�u?�	��t��[x#�-���Ru�ED=H�+�tOR$	zf�Ѭ�(6��ͽ�!͖�����J�Ё��E��%<m�"TS�:i�K;{f��kEA}\7or%e!K��K��``�F����R�̮?Eߟ����L��<��p,�^��̹|�S�bR�`��ʷأ㩦�_�>�l؋�����t�q�v\JC��4�Jr�)��v^�9W�k*��ܻ@�n�C��^I��3�:!qbt05.Lgx�h�GO�3{��qT�3b��$��iq��Ip"6\�PFW���W��b%���2�eX��3�Wx�9J�B>؜^��S3<˔�L'�WO�IFh��e>d3���D�|X `g��;'�J��U:عa��] h�>�����9+T 0��TurZ��0F���	<*Z��20&�+H����2�T�H8�'���+�@���h���ZW3���[7���S���
����@o:��Ӯ�zoy$�B��-<j�~�<VH�1O87>�����u��u�����+>e�z��DJ�_�$Pi����3�ϸ]�^[O)�^LU�L1��W���=��(�b����$�B��s`��^%��<���R�C�b.�{���@���!������/�z�	�<ڮ�"�t��[t3�SZ[�!EU����-%c戏��=���ql�6�=p��M9/{�
��G��Gp������e�H�.����g4�f��͘&T��z0���&�ZҜ��78a����0c�u3�Y3[AQD(�����M|3�RP�^Eiz�%(e�����ڈ^�W��n��u�m	�8&��ڪ���R�榛�@vhH�yi��(��KCW�3g+.s�qJ�V1]��t�PD XX%㓂�e��'@Q��#'I�,������]�I�&���'Ƨ�:�~���=�2��1�5���Z	��<>�����`r�)2m@j��}Z�|'S�ٓ�J��իi͒D�5:�z�ݚ貭���{),fݼ�]ҍ���/��kf�	$��&G���2����΃��K?���_��Ċ�¨������)��s�ܖ���յ�jp,�j\!��)"Y��*?�q�����`�7Y"�����k:�M�}�Է���y56G_yt����씻��U��������}z�ۿ�ߌ�V�a�j��B']5�3n�m� ������� �*H[��������)�:-³�^�}K�\\e��1�T�1[V������ٰ.�n����vY5�ޱ�Ղ@�&�8����M!��?�����0'�ʴaz��y�{L�%��C�FER��T
{�h��/^D�ߏ@9o�!*h��iHM0¿D��<��]��f�R���Mq̬�F�q��z2g�,'��n�W�������͞l~ʴ���ꗮ"L{99��ʆ�x2]���f˧a,I����]�mW�ͤZ��4�����4��x��Z��Jo@��^I*7�����3t&���<�9�;����&�ytaak؅�*�9e.'a��`�w��w@�˃Pn\�P�P��?��xa)E� q�����J�|�C�p�,��|���k�{�]�h$�mS��V�=��׌���e"	�g�iq,�Qow�'v�#S�����	*���U�S<r��5�|�8�*��T�sus��&�ʨB��ʦ�(��XT�������Nx�z�Y J�ڶ��nh���>Ota�jZ=���� �Eb�J�e�����z���nu���m#n}**dM�0�?El�2&x�\����:m��G�Y$ۊ�w1Y�Ss Nq������%^{��>�f�@���:3�^�f�ճ��;=(:h�\J�!6��[��%y�Gq��y�y��H'�X���t�'��ׅ^͑l�������+lh�gƬVƙ��G�� �%�
�����z[-�w��{?��f��)י�&w�(<����|��/�������,��!�=�����6��0�������kw��1��A�>�L�WVq4_��F��ΜS�Nў8��5�d� #ۢb��K_P��&����,�c�r��s���(��`�b��i��i &D��7egmf�IU9�|���ƒv=@��q���9��!G�K��텂��e��?3^���u��~�uhy�w�]���:Gs�IA!%s�2����p��2��kx��U�C�9�ٽ�Yu8`���KG�Q/�����4L�b2)�^A���8�b��B���7���ݎy"�{�3b��&O@0�	��R��=���D���|s�*~��mG��Um�1���nn���@��Eg	������]-{4�#м�ˋ}}X=�+�Љ��i \O��~@$����a��e��cN�·1�� �%���2�3y)8������3�K���;�H��l�'Y�WS�%��ds�j@��܇�������^�hmN`Z�il;(ͷ�*Dg;���(v.$������Jlq��!����*��� �8��&I�h\� J�Go���k�%�S��X�����lԖ����=z}��
�^��4^�L�U��kp��&vzm�l�Xz\�I���tQ*=6�<n&y�h�B|��sr��bKif ywp�0��F��Z��j���:l��Y���J��>�L�9����� 	�Y��9�?���-*VخݭCx!/�����O�D]�Z+�O��Ffr�����寢�o��]���I��fi����v[�jk�]D�H�,L���X�D�YLl��_��P��-�<��Z>QcE��ލ�]:�"*�D�V�2=�ҟ��5J�ϗ���g��L/��'i��5�"��H)Ke"�1�ʇf����?��u	���-m]�iJ0|�H^���[Q��O����vD�-UGurT!@����gz佧&?_IX8��mlg@�������|��DY�]��A�q�ό���9�u�+�7�Q�r@��~}_f0�7LG�!��o+l�MѶ@+�ڠ���'	�y�bv�����%>V����gF=�%=�^ۇ�h1������U����#}�A�8&�E
7?���mQ�F���iɨj��X�Y�;�mf�~��J_MV�I�e��:��\gҟ����`��C���w��rT�
8�~�N�o��X�$�~�<����¶hN̰5t�{��u�s�^�'7�/��!�ڏF���A�����	"{�ޮB�����O��
��b��}�n��71����`�l��;TZ�7��+�=ކ)��Ud�����w�y5%L�M&h���>`��G]�z��ǰ��龜@���(ڐ��&��w�[�*%��7�r¤���t���m����p���M-Xbv|��O�j�-���[�a�f�w6s�����'޸g�ZȐ,kK�θП���'�U�,����𛹮n��	~��4���Oë�4x�x�Vp
�='EU!&�����c�dfn�X�@��m$��L��4��\\�|��=�x���L�9��Y�Wb�W�-�y�L)��縩���d���"¿��a�-�;۬@�/�v�3qS�@��b?֐��]���"(/���m#9Aw\_0�aAB�")B|1@	)`a3|�EPt �u4��g�#q�\c���f�!�1�b��x�����;�P��W :߂�g�ay��0������EK*�3W�A�ߊ�iV�̰�ƫ%��=TN������
'q�h��F�8�GA�JQ4t���>�]~�2x\���v��n�L��<ֲ)\����[t �s�/���u����
c�gG4��Rާ ��7-� ��L(7��7nR.��n�-��m�c�����t3�1�0�^�G�e�~��������Ix#q��w�TǹIk٩�.��wq#�q���d z�֡
�Ad�kO�k����Uh�+�{[�� ��@�\�����2�hm��x�P�v��0�h�.d;j�9\Xj�{�1�n�%$B������6��B0�֟��N�F[�RyJ����.���P���bN��k���&~��'rs)OZ��	�\B����!L�6;��Ez���7�(A�0j؉'c�	P������F�$�����~�c�����2�*4�V������HX2�dɀ'����x�!��6S����'��W~�l�(�x@���hr9��	-�_�	L�Q9I*lG$��İ�A�燀��Q��D]ġ��w.��Q9H�Fɚtc�|�	����?�����c���#��8�X���C����D�Y*1����B��9��g� �m�+�}�n��[;�s`ƭ���M�r%1�m�L8��-n��r�����[u��]6N�����яqX5vV?�]`Xz�&E��/t�3��*i
Ыv�����8q,s���\�S���Q;Sw3��rYpNR9�L�
]�����?*S*��A�9kE�_�j�=ń�����VE��b<�����@nm�h�st�k�ߩ�5�3NKn~A�����hFƒP�
cվy�hNV�c�\`��܃`i}�� ����ˡV��g����fJ��Vt)��	��w��0�k�E'�3\��;)���[A!��	kA;A�����'d���8mI&��p��tt�8��q������'�1Iy����E�f`�����>�$�KM�������qH<��/a��S�I0#9�N^�X,&'�����({t�R]����J��D_䢚@��h8��s�3���G�s�̜<Y���c�oΤ�^_3� =��OJ&�������]At�O]�;�
|��|�e�ؾw��<HmF5����W�[�Fd`����.$�ՠL��g�w{�)���m�~��f9�u���ז�݀��f`D�������h���Ƕ��}?�*&���=���)�k�ę&Y�K��jҩEi��23��v2��/b�<�'����61"�����K���lA�!����L��n������K���:�x;p�iU2sRfBh����p�^��)I穢f�=�-�gz�b�>v���{�l��Z�c:��s�g�k��Pq�(:�[	ǟ'�ڷ�w�s��^��i���"��~I���d���P�"���&�΀�k�g}�9� ��Ku`iF3Bl��sm�����N����XQ6��&Uᔞt�����s�8�V�)����	/�� !t��غ�Ѩ2�f�
;-���L��+�G�jk�2@sX�Tu��b�^�l<h7��_L��R)�:��p\!����閭ߜ��h+J����/�g�}���T�Ie�O��N����D�}+�"�rSF1OT��*�Y�{m �$|t��Z�+q�I!'�)^66�8�h	;ؖ	�L`8�"H� ��������j�����z@�9��wp�-��2�+^��	�ن+�l"�նƼ�+j�t�=��f׬`im"���l���ӯ�:B; �y?�%��,�Vo�.���I��28�n��M �y4���7J��JCL4d�G[���,��qm�UXՠq>̃X��E�g�Z�jbR�2�S=�+0�d�f�x��ޣ���>TȤ�<�X�gDש��Z+8vI�=j��	{��j�Z~�����>FE;�d���"̇9O���)^�ݑU�n[A��Po��ԗ��W�o����Կ8��C�'�9"��Uw?�m%З"�z�{X�H���/�=�mkARE��Jއv?���Y����u2v2�=g���}[��̉tv)Ɇ�4���աa(wf�O�"�� ���
O*�U�VQÊ��+���S�)����RzN�7�M��Vf��Z�?�i��_\�H���Ea�r-i�RP��!l�ܘ������y��\i��ap��?؋����1��!�~�*�a�4���~�bJ�K=��#��ZˉV��wD@������*s�{b�"�@�/#�x:-u	� �P;�*l cn_`�$�]#��D"�	@�Q6@2®FP���[���|#nx�?��ʜ�3�dr�kyA� �����Q
\v�����S��Rm]��{+t)�5)�6�l���(TsA�E��9��G��ؘ������������h���	Zf�YfT��˪8��:G|�+��0��Wu(�jL٘��**����~��?�"0!�'�Oo����F3���_��3����l'� �d��#B5�"���DB"�P/t�̰�Ř��H������Ź7��\>��ւ�~B`�IYҙNϋ����N�����LT�����`������7��%iS蠆��Az�S��M������1\Td�����xpG]���k�2x�h�/U��ݞ��z���*��[%b�}�xQz��_�$����g�A�b��Y��0@��L��!TY!-p�w�YEm�e�)����0��)õ���1���f��Ǝ�H�y~s-�v�T~w)�:wt�Х���#��g��1f:j���.�q��**SDJ������M����T�:�/��"h�j�N�4a��z�7�ܦ�ʷ,GS��"���p'|v�A�	��u�|��Y�0�w3��g��="���̃~XF��y�)�w>����P�Ɉ�kjk6�!�x��R�.����'���B�:�x��V��Ut��C���!�*�]�:$��7�s�y���|Aw+zH���?-'��B���(M�J�E�ߡ�P�1�#�-4\�h�!����u�Q�c��B�S �!^�4Fn��Vn����o�v�G�?PS�ӽ;�n�������s���}oF�;�H����s;Ɋ��n���g��a�<��F;-�;���w��y�;�����W�q��%��aAT���L��DZOA�b��	J'r�������E�h��`�秳�
^Л�O)��̐+�A(QQ����r�Aݯ����O�������·P�ҷ�����IQ^	��a�z7�x�m�I�bDS���6,�G[{�!4n�������Lm�7��u���%�����!j2]��,�Td���w&��^3h�͸�������/]੔�Gl��(�c��f�뗕��CY7��T�&�V�����9~4��_}V�n�u��[�g�W������G�X!|}@�%�4�n���I�D���H�tQV>����:`�&��e�]�W�\p0��8�Z}��0�w���MY�+Q�E� #|�����i^�\�F#����Z8P��^h֒1yn�J*�+�X��8e�o\s9�"��x��| 2sbã�W祲�?k�w.�]s�?�U*���S��K����-�K�����q�U�Q������.�0�y�ɘ]Z�*Z,Yi��.�{ПS�d�z8 *)��r�N��k�a���d���+���,�Gn1o��#�p��&�X���[�&���2�����!%b�#;G��R63%�WP�{����R��B�Su�h���&�,'@�b��3��I%w��A�y>�x�ؘ�gÁ�v�6&{Zk6I�W@!����xGƢ/�"1�2oц	��,���<�� ;N��� �8�����i�����s���b���N���_��>>-�}%n�\��5,��{���7KC��@C�pm�ӊ:��	�i���MhG�.�&Z��X
�B�/�=�Y����o�=�)Z�a���:��Ϩ���x�w�p��e>���'��+<�����Ȇ^�j��;<�X!1�W_�)�#=���Jpq�Z���4����B��"�ӥ��^��ܳ��2X,�=�ֳqd2ۂ�ѯ���Lj��M����j��G���I�/�#���8� E��ᒥו�[K|>S����fG9@�h���j�y5��~(H�+ϔڲd��%H��G�׸ہ����)=l�0���g`
�y=�Q>,o�e�e�D��J���v� P��\P��+��!�L���pnI����+2ϯ�`��U�>�a��	;M2�����^��g����	�;o+�}�R�]��p��A���9�]D`yف��|�RE����:�)�r��Ή���s�ʋD��fJ��T��� K��������>�'x�q�����l
���B�S9<�����6��� c��Q�qIo��^���1TQ��>	�U1�jz7Vw�m�Ɠ1��0�)#D?����.�^����RXq}�f_I<D×vK"q��P(MJf�b>I �x(6L�Pz��\�^e��}XE���U���(�N�_ş�h�l�DLw���e;e�w��y�p'VkF���F�������s-d���=��2���59-���)C��JG/I��4y��"s�9ƣm���	J�^��Z8	�.��Sm��?{�i~�֔n>����]w�W5��b�zQ�ۛI�5�� �4t�ZY^%�=U�����W����;�=�&� j�Z�g�Ƚ&s��.;�XV�k��C���q�M�������,w�ʥb1e�'����|A�1FB��SS&9�~e.�z_R3��g�O��a��������-� 6Z�`�����zY3�-9�����ꂤ�� 
˚ȑq�ed�яڍl���5�����\��W�Ӷ����ݕ:�}��K������|yo�H�-�G�-��CDѵ�/a�m���󮐿=�o�:��R���\���R���2�#�n.�۽�������$8�jn�����g�ƣ�L��c��m��d*�� ����9*��㰵)��Somi'%������KI'xc��{b�9���b(�<?�v䧷T��{�p�V�:}��(���p�aj�BuG�ˆ-���h�=�P�_��R�ߜq��9�^c,
�z-���4�n�Ou,V�x^x�,8���ǥ�'��������V2C&��-ItF!�׮�|'"T�����Cd#�@@�t'��ʽ+��1*�%FT�VR�}Ky�ʛ���Zhg�A�*����hd|U����2%���gS�C@1�x�|�ȍ+��c��4�.��P��^!:��R~��n'gp�˖�[G?�ۛ�=�3��W�~~�UA��W�X�.�:��04vZ%��������\~٥?d<��~���ϡ���oh粩l���� `no0��J��	�h��Z���i;@0��s���N���A��V��sC]�Vp��p��/�lξR%���7��3{H�v��Ϲ�U÷0�.�i��`9��ާ}q���l`.������3w!��$�(�~�A���ۛ]2ׯ���M��+i�	9��X���3�A]P���xL�T�q���2�'����Fոs��i1�������)��u��H��9֔��N�^�Tz�?�MR��rh�ц�M]�0�ե;�.���"�`�ޮ�Cs<�L�Ӵ���s��.9�e��3����՝X��Ex�G����B�W@���u�yd��r��6�*�p��|�|p�9�C�4����������G:t�h��}�Z��vR�D�b��z�6_�����|:�T�1��kL]�<Y�3A`��l���T�9�/�6M�7��m*��)/� 2^�W�E'��q����Hc`��e6@1z��)���6�0�+�S��'�{����������k'�c�|�?�;\!��M���K�Qo;��vi�T��$M{�'`���b�a5*vL��9L�-�J�g�b�f�Ԇ���B,�t5N��_&U�q�J�E��x"#�H���O�w񂝨�9&/�_�}� ��!F`a�����:č#�@���	�7v
�bm�ݬ�u��멎v�z6,_�������t�рd������R�}/$��G�ӫ��*�w�� ��htݡ�b�[�-��5gk�l�G4w��|��b���f�9 ��_^����,�N��A��5,@���:?�^HX�ky3�.���J�
�SC�xuP����VbF�� &仟1Bxx����H���T�JL��@�e����C�It��O+f�x�{����^�b�(d"Y�S����%��2�����m'Nۙ�WЛe����(}?�BP��	�������"
��☄�%�og�����A�D�=G��7�Y�� ��|�Kq�9�����7	���b	����.�f�M�;.��O ��Thb�S~g:�FD^��+�m���k�/�F�a ڭ�WA7zG>��Ԣ�I�KC�\?���Ԁޡ����I�q�� ��h�V����;���F�x!Dr{��\x�;̿=�4�aN0����1����5��ݜ�RZ>�YqZ���8�{B����f2�ʮ�ǲ�Ɇkm�(M)�1��pu�7�zLA�M�2}Q��p�Y["w����o�y�`�㉫��D#�cK��\�p#�o �M�=I��{,jl7'^t��W��:od��n=�P�V���A�m�B#�}�!��=�xt�^�z��İd�O���=��)G�$�sS1�~��ߝ�ȣ��okl��)�!�ymA�?���V��zwl2�q&�/S�X�*�� ���s酵C���Bt<'|`@E(���ݨ/o��@��'�T����b�������&�SN���Մ��6%�y3>w�§Џ=\i�sP����	x���/\Bt��$2T
h|����O����7�M���"�37�j�4l@�sO�S4�:Ө!o�*���X*�ޥ{�l�]ZJ�@J8��� �����f��,���#9�G�R���YA��!w�%>��U����r=� ~�U�/���_
#Z�#J"�	�v�xnW�tX�O��r�j��&@y����=0��@�]�?ZH���C�N����>�At|^XcD�y���*�kZF̠O���Gሸe4��y��]6�X9/�����óf��L�;'(��8?���V[�i0�y�/�.f��p<�P�� z[�y����fF�+��C��]^(,��jDҦ���S��҉.�[���H�.�,����a�[�M����o,&���o��iߎm۶�l���N6�mol;�${b�����}/�NM��u�L�}����"�N���}���J��
q��oaĪ\S�j��������f��3�m�v5��D�0kg�E�kt!�V��?�
㗟����j,uB�/�C�s�#�/+��VcUh�T�̎���/J�|W��_�QG�m)5+;~7�����Y�����^�1��|p���@�k����j:���Bߨ���|w[4�s��O����.���k�p7T����}&A��w-M%�]�O�m�*�QkT�|N'��>�?I��ęE��#t�� t�s6\�����$�Eϻ
g3}�+eٯ�g���w�iK�Ed-��2Ζ��b�y�V��<$��c�� �|c��R����󆔋��2����ݦv���s��l����ݺ�F?���uXK�UҌ_����i����z?�O�-ݒ��g*Gcgm�=�;�{O��e�f
[��Ǥ���P�1TF���^�l��b�}���v��U�7�	����ǽ��׏U]c���ZZ0%�x��9_���DJٲ����='��<%F�ߊ� ������A���o�A���� �a,<�t�f�ָ(��e1��u>��串J��dq��r�r�����pJx�>�!x��c�2��D=���3�������ۍ�hR	�k��|�R�{�q��%2�~ȝ�Ć�I�<*�w}�D`��ak�;��z�7ax��&8���[7oH[�q-�#`5�H��Ɠ������}m:�<d�+N@o�&|��IO���ɵ%��,��H>�mq��������k(�@Ƭ�B-�?6��◻t|�H���"щ-`����kMQB�y��� �1��&|�7=l��If.�I��+�I:����ieO��:���n��à��-0�^�e8fu�4� Y���6�x�j�Ր���d�@x��)?'��wm+)|��'�o\�W�xa)���!R����0w+�1g�g�u�Ĺoo�k?؍��B=�4�~u��Y�uV�Ԋ�F�m��� iZ�;6�{�(�¥��7���E�*�_�؊�ZA%���e,�:\�5ꏗ���c�k� ])�G�{���M����'�����P�̐�rm��a$3����~^�y3��+(�䠠N]t`�u��� �6y��dtԂ�Kh�	"���5d�	B�+|�%5�}1!��El��)7����D�F��gx�̊��4���&A>X'��a���t��2n.������}jgXˠo
RK�:�7͗��$�����q��9��������OX��<t�fz!d	ś5[���IT��L�\�-C,{,֑]/�\&:#��"��B���.�BWʷ�<��蕱�#j� zU}F:�9g�j�"+XI�f��m�!�7�2���[����B�;���Ϯ��"CSy����9z�F+Ǐ��S���X���X���w?�O��GPw�+�r�u� ��(��G.Ф�DA5_Į� ~��ԅd*�����5�%���º��7���C�#I8�2�W�鑽U�Ovb�ѨAil�s}-��ܫ?�1x�JR���')���]�L�H�=*����F?��>�@�N�w�.؁h���qkYg���|]&�J0���t],�W���s`���P9Y�L���;�߉4�h_�Wn�M�u8Y�������%�%����+��~y5|iw q�D?�����H!�gD�����Km}���~<�X�z��n�$�������@J|�X�E�����'� Aj2�5�2dÎ��m��2�8�NO�tB�~Ǒ��/,ZI�>⩊� S���3����2Qo��kk�6-����/�jw4�\ 2�3|Q_Y|��@��Pe)����v�BD]��f�T�D�4�Ĩ�84�� ?���r�V@�>.r9���ÜO�9����&S�� B�a�9�*e���w��:��;�w�3|:���� ʹ�Y�s�1��.�ҹ߼��V{L��sscm;5긻�v{Gx=%�ZAJ���oP[R�x���ZT�2��h2T��f��I��0#�� ��������'���ĔM(CJ���^+���q��b� ڏB��E���:��������/>���q�����Q�dQ�,��c����b m[�9����W��{�n�o��"�U,�"H ����a�Aų�(KO�]�v Ǻ-��%ɺ��a����U���r�$�x��L23�
�7~=��^?��I��y��n���A�!�d�����!p��\\�7o@��xX�ܢ������Kε����QVZ���J��`�wd�)x�ZK����>P����ώ�O%ċ�ſ�e�e����;�����z�,�d�`���][͕I.�[���7
y]�~[�ebn����s�Z�[�ǖ�J���o�G���܉�_Oß������/|2 ��谘>����RI��ЙxǮۉ=5�y����'9�:�U2E�;ՒP��E�ǟ�W,�K�Ł�"fۺ9�s�6۔�] ��^	Y~��b w̾[c�W��o�F�2LƜGl��F7�@��rq�Bg ����,M���t˧`+$gyw<���+��N>�7�˵�aŃFq���?��
���E}��l,:s�4E��X��],�iT��v�`=��!X@��cV�iA����<O���'����I�LcHR5��_f�Ȕ�HaD��K l�9H�rI20>����v<����I�WFIwd��g&T�L�:��j�-�H}1�m��Çty���+!,TB9�	h�[��c��H=c�L� �
}F�����rZ'��D�;�Gp�C䢮Y��g ��2+��T~K��m�����6�q�p�xz=@���`R�N��C�ݵ�%t��O��U��W���`��q�c�;��,�vQ׬7��~=KT)D8*�Q0���`U�Xk)d����R?PF�j��n�\�C��Fߟ�Fö �?��j��l�n�����E"�T��1�3$(2�<z�ҷ��}=��wlTe��c NL�/$Y�ӕ��џ�S/��1�,�8���`Wj��tҪA�2��G	,B��i�\����!�K�w!�:Imƙ��[zUڧ�a2�mvፍ����&	��v��ȸ�YF�{~O#�x���m�����m��FƉ�R5�O��Y7��7�|�)o�������e���a��۷:���דH�+Z!j�u�K��+��{g��rYW+ŮL�q��XnK��4dP���N�#k�̫;��/*XgZ]o��X2��u�_&����,�$+�{�u`C�K mU���]�_�!;C�fF���F�aJ���1
�?5�V`$6Au�����^��9����)�Áza+�ڂIxy&�p��lӅY���
��ީv��=���N>���=�ܐ Z?SkɁ��C+K��ꊑ۶�{;6A�f[��nD:��zd�AB��e,�x#�D�Ƿ�����7C����u!H�j�n�^��L�)��Z��q��;�W\G�ͩ���� 3�	V����+�3_�^��*0�����6�<�,�7���.ND.ȮD��������PE򃞎Z��&$�i��@�����X�*ȥ:>v~��\���^������^�Q��һl|
b�ww/"x��fY�YB��{����n�vŦ"o�^d���HH-��T�$���?�BVD[b>�+Ky��t<	 7iA��9�Jۤ	v����/{��@?D�/�%����U�����)�^��-�:�zB�Zz��}�b�2��6��t��UI�6�=���A�����;bᩤn��ȑc����)}��a���^˅�ǹ���>�	"7"{5]G�O*99�/���}_iVi�uD�z��X>��,���C�>J��T*y�{��:WF>)U�'�l���p�����<�M��~���Lr5M���
��>�L�>�r��ybQ�l��u��6D�B�ʀ��*�#=��O)����*-{o���P{@\��!��Z�\�7�o�˾�1��{�Ѐ)�֜o�e0��$�:��#��M����@�;�%��G M`�k��Q�NB�}�l ]�r"p�q�3ő�t�M��SZ�́{�]�ȫ!��_R��)��)\�3�z��sk�FU�c����	H)�����j���F���mX�a�e'��
��zn<=y�w���Έ�����-}��A�{T,��ʕq�Ȋ]�Cm[9���4u�並i�����;����,�g��J�mfЖ���#�0Ta������,�NC�8�c֝��V�́���I���W禍�[���_B'8@� q�ٱ�b1'�^M�O/8 N�E�O���N}�I��Q���'߃ �\_C�Q���)�]��Bu^H�C���b��y���n��Ī����O�l����� �yO�Z
�G�f_� �K��⃏H^,폰�|����H\!�N�Q@ �����Vs1$���i��ߤ�.hM�����DQ��]�8k�d>����L��rw��̃��e��⪚?đ�X�A��;���	Sl-��}���z4� ���^;r���,J�B�/�Y�&�F�VB
��e����]�i�����&�g���%l�"vrs�Sݞ�vd#~�?%��A{,���[B| [���ojΈ�O�FbX��b!��7s�$Vx�	l��N͕��|�*.�OK�5i�W�KJ�e�\%�*���g�+c�eX��zz�n���d�_mǥ�[Q�.[LtwtkBP�*m��@�S�� d�z�Ը�&�rH`�,�R��gl|4�$��r[2T�KHo��'�Ք�-��,ࠏ3yR$�!pxӆ�B���]�e&mM����kߡ:��Ȧu����-��U��6��I`z���yyy���M���7֖(��`=�����p�A��ra��@�_O�]TO59���VDY�� �z���r��Ф1�tZ��Ua�zOk����c�ߛ��GJ�v[��=!�D�*1h��p�����F�����=� ���D����)��
�2k6:���p��_�|������c�hрe�B����lWrծ����n��|Ѹ�p��@�5{������V��H��[ޣmO`�ϜP:0��UW�$o���G����i�0tg~Uo��U��fI7������0����1�0���)IJm0.A��	���[A��ඖ�Ɨ"=����}�����c���X.����Y�H���
f��l�P����(��J��eS�zr��[�g~D��X�����No�|Fb��q�X��Ǌ�28�sRםh���G4�YH���4s�a�6�fɣ$��-mrH/�%������e+�R
,���DR>)�����R[�,a���snUr���T��U���e�egn�9���;S$$�ec��%�s���N�:T,>� ��~Mf�	�������[8	cS��yz���8Z+����*p�f�ش]YH�����ޘ<�o���� ޛB��2��GV�~�/��/!r�e-�?^��́��8������8P	�Hs8�!����2=d2N��7�)��k��vg��S~������,��,�_�C�18:dm�v~&)j��rT3/D3���?�G��ߗ`8`C"���횈���2��µ��x��j�Bh��<��U&d~0Y����Q�4v�n�Qb��|�vY��:>&I����u|�*t�!�:�,���}�Цx7�~�u�yw��\akPux�Y�ͧu!6���� ��ʘ5�S#��x���=>W\x�ۑ����uC�
=<��0w�����֖�'����jk�%�t}i�ٓ�qQ5�f���b�0rr~g%��:����@�>��8�iOΚn��A�><]��u��4���"��(2kAu���<Z\�Tb�9}򷮧:0�	����7<��%��<������J�Ь|XU�����Fr06��!3�U��?��Iy� ��6���9�k�k`�ć���řC�ߋA����;�KJJQ�/�� Gi��kh�Ԯk2�^��^���_�n�n^y�VC����~+������!��ק`���4(���1�C�Hr���鶳�Ė11\�p�'nhvdd�"Ͷ�	6����1�$��9W'V��+o$��d��c\_:fވa=������'��E�3n���);y��Z���>�ڇ&\�u?˶��	��T�l�����9���槟-y�cs~#�݈�d�:\��/}RT'��=}}�M�w��԰�]-5y��a�w�B�>���z��==;����~t�R���������g49�4�(A���,5��d a�r�� �R��4�k#Fv=��~��t� }RX��1�Ġ�# �/�%y'���A~��莢���/���|(�J*p���d"�����q�sۏ�K��R��ɴ|�k�(1	���SLX+&��
M�8�������؇Hj$B���~�yJEW�S��Ќ����%bbn��QI��\J���F���D�kS�4ݪ�TKt�8���>�\|Wd�k�G�"\���+}Y�?Y���E[ߣ�U���@����d�KwL�UL�\�~J��s�l#���Q*\Fڲp���nk�!�Vҁ���ɪc1hi9���j�b3���;d)l����"��V~{/Q�G���D�0���U��������8��m|<O	�6�Ud*a%��K����]L��TK����	�x��m6)���pQ1L�
D�ۖ�:�,<x;Q7R�*L�b  ��Ϟ"�m��f���w6��K��U/�3�������ǝ�,���5"�J�w_��6��Q����W 6�5���!��3���{��֧��fjo�n�;�x��b~5c�F.S�4>�WA��$]�w{�T9���(?��r�X��J]�q�ۮ�8�5]�z����/�o~tq-��鴼��h�Aco�(vvL�'z?K���y ��}�?�>*�L\<\U�70ړ(]�o�'"����3����������d����w���{q�NR\T1���K�������%Έ���z���R�Z�ͷ��rR�:�^�j�W?9�#TRPp�^$^u�l�|�4��E{L6��el������)��H��-���x'���	bs�7�w9
Tm����"@��=N�9����c��R����|��]�e��������3%n8^;G�D�N��H������Ū?J�0�D�l\'Օ�^�����F=;R�t���B��Ɨ�y�����Sp�E��i�X� �� ���7[�J��$��Vs��ѳp�����-nI�{/��U5���6��* ��5��C�,:J�u�yUlu�bȭ��١�� �y�ƀ��v�!�u&��닧�p�4Hw�RL���7=6��V��!���U��B>PM��ԁ���M�{��"���ʕ�b�B�������dG�c�n��M������3[O��?�&>�F�]�%F�k�"jM�\�/�T��l�U���C�#��SB�R�^E���o}(���H5,۞o+�{��������4c�6-�9� +��a�l|vO�C;ly��(��5�W}ҧ�(Z'�6,C�Kw?*K�:�C������Q�p�_m�_-F�"_LE�{�D��A{�@~�߂�6R�
[Ä��E�~]� z�G(��i�fi�������׫х�XN�׬0i~�l�?�FG��T�RRP��N���e�/
���*���7��	�S$������K�fϷ��$�
p1�=�2�tP�㛧����V�"B�'9�8Yn7a��/�-����m�p�|���j�J���"�ו�ݒr=A�7��*_�i����@���Z;�у��G�<Q�츟�F2iQ���o0�f5M��у����{kps;|J�B$z���l����K�����!j4���ƞek m��oc�N�e�ٽۿ���P"��臱?������k�-�)O�9�Ֆ��
��zI���Ĉ�G�5h-]p�ȴP��Ѻĭ�bH�˪*��%hﻗ�7+/�YN��oi�)6MVk�zհդ?.X2��o�p;o��������x�,n~��Y���C:�!X�p�:��P���	0~id'��Z�Jư�#��{4��2`v4łm�ΟQM7�"�Sh��NAI����A��
#Vh-�~�}�G�������C�z�5��E���W�sgZ�{�ǡܳ@ᾝ�܏pSx�z���%���,iP?�'�Ϡ#�G�)AjД�چ��Û$���<'����{�k6�I�h��ا&� ������b�P� ��?b��/��E�į�w��0a1���\fl����C�P�q��>�U0iJ{>U���b�E���	٠n�|����T��E�ڎ�jQ��Κ���سVeb���ۄT�V�v�^�+o8�&���~N}�ޟ3�������ī`�e�!�GӞWjR�RX�]�`bJ�u3l[����S�F�d9��q�%���<��:�zI�6�GG�G�Ю6#3���P��͘�|6��睗�%2Ha�|��&�Jm�$h�xIU+�\7r�[j"��cQ-H-��i��N���B���Q��$�LB����U�:���Z�[�(�vsw���)����s<-�	��OV3��̔�JcR۴��I�#��
�Bm�ľ�* 7�B�}��i�B?���F1���`��2��s���I5S�!��=���~K�F�k�ϡH3-�GW�����e�����C�Hv;?�j��>5!�]�A�]!ӛ:��
?+*�gSծ>�~�~�,�����IV�Lv>n[>��#��QƧ�Up������
D^�a��z?����)��?[����1@=���^���"���S�'�g$Ֆf�MR��v%s�ճ�h�9�URh�U��X��F���4��G���.�������j[�$��{��h��!���׋������~����mv_�U�2ҷ�?:�#���p��f�%z�V��a�ʾ���zӘ)�ZR&�/C���CɅ'�Q4�mh�Tr�f�z�{2�e���9AE~�p�	�&�<�BԠ�h��Bd�ş��п�u(�jl`{�	��/1���u�|�̊���W˯�n`�$4����^JΈc�ӖrI�e5l�g:J�+\��tgɷ����>t����"�B�L��Ӫg��\��4|�p�:w�/��,��_#�{�Dn��nAσ�%��\��ӑ����6�E���Ia�t�p!`��̨��[�^͜ �V8���X�o\!�A�7e�W��Ч�ko�W%*��fJ��g>d[��������U��0�sʆ�$�ܐ�\�}ܸ�ؽ���I��B{$���i6x}c^���k�y�LO|
����>��V�{��fJ%��h���߬����.C�F����"��Ge�	{0mĶ׍�c�qމL3�����ï1e�G�-��P���r�e�B.��7���z$}�,O�����"H*ژ��Jfz_�0J�pQei�n$B�>�N3z�ظi�)�b��~��ƻu ,��'<䜄��ӮWUL�9�FuR�r�H� �c�Q����ާ{�����y�@NIܛF}̞.��sQ�0u�XÛ�Y��
�jY�I���q�B����v8�����|�h��(2P���+�?�-���o:12������³����5��T��=u<�u�N�)4\�}E~%u^d%��J+���R�'.�x{~������Zw}W�����r6���H/:�k0����d�Vp�;������y�͆�K�E�4G��^���g�~
��q
�W�������P����G_R�l��x��@}�5z�|�.���+/^zX�%�,�W���~�	GR]������뛊	n��N��Ur���_�>3<F�Uh��y����|��ʈGG�������-��ӇD�_�IHB��p#p@,���䈖
\
n@@:��Z�Zhw����̤�k�y�{��_��9�n �[Y�{��Au��Ym�|DϺ��>���U���9_���q=Q���%���~1 ��>uM�(���R�uts>��S�o�h���LU}9�ԡ[�.;��t�����p��\5��1�w����<�J�p:,��p1���*�C�ݰ�TH�:�������LJ�8�W�����5x���LeKȴǜ�x�-?9��v#g�Wz�Z;�c���M�մӧ6�<;�Tj�cU�݋���?��3g�]G�L��`_��8u������V�q#���g$=u\n�˕�Dx5�@<� �4A�j{�/�� ��g�b�E贮��W�	����.�7;!���/$� HM�Oa%��F��ⓤ//JEw��m����s6�`a���b
cd&�'�3H�E����[%M�;n-S��1(	qs�q��;�8��N��{*�4 ��_��.e&�\��Jo2�8i�:�	@iB��P)��7�����7#��F=(�x�By����0�L��L�^d�N����r^��BW\���Z-���WBc<��*�B�\�~���=#v�o�
<���k�:�c0�΅H�e]p���	X�D�<)F�$��.y�i�r�q�|k�bh��@gvq��������A�?�.��Kh%�q���GvA��?+���}h��1������|O��w-�0�ꇐXp��`����t�υ4����G���N��[��@���
9:B���A^C��6Ȫy�+��%��:��zO�y'ܠ�f�W3�W�FB��K���&-�o.������|���<�w�֪��!)�������CT��U�!{�� �#�J�D�4l9�{���to�C4]�uCY�8$�|\����{M���0|&0Du�Wr�� ��i@�.��Ψ�'��ޝNO'�5Do����dq�K$Q��x��P)��9h�hi��� ON��H�W�m&��:�0 qʺ|X��+�T��86�6�<#�'h�F�6��7{��f�	�y�Ѿx�"�6��C�L�NL�Veً�]'�tz3{ei�Ws�!B��2J=gk��MY��O��nGbݗY�ڡПx3���xw龜3q&QP{���q��A\b�\����.�eS/�Ѩp��vt�NS�!�c�.1圕��S�q���3�~�������bh��G��ɡi�y�u���#�����dL��O9�����;��	!C������x>Õ#�y���,���S~�_Col���k���H�~=��9b�<�����?���SS+�y�^����С�+�d�|U���X$E`Lݚ'�������Y�̲c6��j�_v��Gt?O:N)P%"��Ε�i���L	�G�"��r�z��P���V���H���[�HJX��gH�c�|}�+�FԳt�L`D�?�	�H��%��x���8�ᔂ��-���[�]M�V4�8
���n��R�Q���('B )/8�f�+F��?r���*����@�z3؍�o�6�eNU�w]�O8Qm�0M��/:!�AH���|Tݩ��@Ѣ���(\*�$����/;��*��p9}��,�dQ��*�Лξ#$d<
"lM���-b���1U?����V��
�3�Mb�!�e���u���m��N/��%էA'}�-��TђzD����
 ��x�5d�:� �nw���}�n��<0�����l��CB��4-���_������@��z�&��XT���E��Z<||����=��aP������yK :�p�� �6ʰL�Ue��=�UD��T��N���:Z_�&j.N���y�W7��̅���/�0���yc4��-�#Ax�?��� ���,נŮ�e��!xķ�7yY�Nш4�(��� E(��5Iz��o�0�se�sG[(�u��Fה8���^Y:����K���]0�)��8��l��6\��B� ���%�<fO��(��4�SЇ=CϼumC����9�����9Ê�0#n]�'�(��l!��d-����3"��G�0#%MA��t���i�7�7$j��M�0҉��e��	�r��;m���᥂O������]�\8�b�~)���V��T�D����TЈ�MMӭc�JõJ���'1�m6��?'��7��S*d?�%5�Q˜�������/fj��w�Y(��t�~a*ә؆:�r��)=�4��܁�X��K��ax�pܱa��^�D����n���G�xXQ(m�?v":>Z����'��{�l�����2���W6ڈ�����@?�(n5��Tǟ��6� Of"�.�x\�d���A��Y�}��YwA���Aӌ�./^Z\n�B�����i+J/�P�B�ņ��d9Re�!;4.�A�3�Bt�mU���չ
y���M��wz �$
�8��9�S�CE�ov���=��],~Jr�	^�^ȣ�EJ��<��e9��`���D�a,	|��a����tn���B1Lq �ٱ7��G+�|���7N	�i��9~�
n+�q?@�0}I�k��D��=��L-��v���vQ�
&�?�ЁH��6�4_�3zx./ʗ�i�>����ٿ;uh���d�G>�MN@R��Z<|'Pp[��*"ްr��h%���=���t֡��ռ;��ڪ���zC1Rz#����t6�̈́y�ó�1�quP��@&�ص�ʄ[|����3h����a��}щ�*��|md�����k���I�on�,�F�2�A��#h������CO.�t�=�hqd .9�R�������tm��ĥ�#4(���I]�c���i��gep�����a@�ͩ�O�v�a� '���/AO?,��t��|��	<~ѽ�k�/�kwB��؍T�?��\�c�?�O��ۖ��U?�L�Q�z c�ݙn$��D0Ɵ�ً���E�D�'B�2��Ȗw��X{6]+1�Ī�,�Հ�ng̐0�#�Ӵ��,�u�JiAF�3��'gm<}�������0'X�c3P����u+���Cn1d�ֳ�?/u��zޠ����_Wh�Wk4��EN��
	2N��\��U�-��B+R�1r��Y٤���=�]�/�z��ơ앥�!D%<7��w��Φ���ɋ�J�y�M���a�K���m�}�����) ��ٽ�Ve5�HSG�5"/`�����6�dcGH�jP���^}���[/p��c4J�;M�K1��a��u���'	Z]���8� ߼Y	�������\G.��yfs�8��kH��ŋ
/����)�I:�A�W]h��B�E1)9.ډ��7�|OP��e�{�H.�7��cn$@��7�=�R?p��W��O  V�D���-b��K��Լ2�j#��x�h�,��kI���qQp�%ȲU�8�Gg�?�z�v��iZyP�W��~�B?�õVʼ�1F���RQ��OT}&;z�j���₈`�����e���\>�r�"w��ǂ�;�����YT]������k߁=U�~h��6����1È�9�%���� �8��^����DW����OA%���r���\l������-v��O$������n�5k��fv�j�y(����v�~N��[��n#ٺ>^��8wY��h�·��̆q��0���Ш��D[�+	�����N��5����)O[��O����}V�L{���X��ы��I�=�+ ��m��N�E+t����4-��d����隗��[T�0n����,�G������������肑�PЋi�m���v���������]��#�T.^J�8�]J-R"�q�Оf�O�����x��^bkwŃA�����"7�&�>!�C���O�� 8��I��;Ơ���u-�r��y(��l�+g�G
8�����:Ft-I�j;2�6o
"F$�6��VN<[wܙ}V��3��Ap���gq�nˢA�HK�<
n^���������E�O3"
<�uc��J�h�/p���c�L(��+ǣ&h��xtn���Ҋ�#�*���W�R�ex,b�/�-?�n������'�~���;��^zb�(��<(��=ݸ�-�"�|yֈ�E�G�9�00�U�[�A��!��֙���EQ�:9A�~�f������`����r�*<&�U�W��8������p>4���_��� ������ke6���+�mG|���2�\��y��3���mx�ް����y�N$m�ۭ�ť�����z����j���7�ޓޟ%��e�I]����|�9@�݂��b��w�溺4�B����������Y�}���Ѳ�j�)c��\k��/%i��i��+��V��O��7�{<W�D��T���$�!���ot�[��_��`X	�A��nNGz��<SX���C��+_�W����	�!��IS���Gx�'�&���'�PF����\efyX�A}�Fn��(�s�}!8~8"��x�9���*vB/ђ�J��*�^Vpa)4�pE�v�8�<�� �"p>A��{26!Ma���6̻�0B!PA"P&V���PѤ�h�RX�^�^��M�w�)��@ٳ�����e���g�0�z9����� ��_�C�㬺N]�I�֨�?�L�5m���Y^T%�|+�Y	� ����?�	t�=H�B�E�7:$Yġ��$�����.e��n0WϏ�`�*�?�t�ޓ����%�F��֯��y��́�dg�\��ՙCluWw���8��Ipnә3�su��`�1��ݠ���R�,P �_��~�i�z�2�&;>���:�*��^�:��?���%E9ɉ����Ӱ�Z���:�����>ٻ�sg6}�ǟ��o������!m�`��2>�<3F���D��&�_U{��`*0��9	�����]]���Z����B�ӚU����MkyXi([�ׁ��ƍ[,k�b��'���A��c��A��A*�>��Mc��8W����.��Ԥ�J�F�[x����j��$ 7���G=��.��.�_|a�^��֞������2�Xu\��tG_����Ҋ�LzŶ�������߄<��h�9�s�jOX)�Nn�a���cb�F�Q�6f��@�U~�%��2��-�㪠s�����y$ ő,l��YW�!)��=�Ѱȉ�w}��X2r�)f11>ķ5�G�̥V" ���쾢.L��X�\~�0�ܪ��ai�)'=�T�z�2^����A'[�t�'A[�(���w�-�-R�Ό��.~�'1�ӻ���ޮ
d�B���я�o�wn}'���v�~�:XwR�vLJ�w-�C:��$?�m{?��y��	H;�h�Z�Q�ѵ1���B�^�qP~3(�&�K��x�.d�ױ z��>�ޣ�m�Ԡ<O�j^?K�ǖ�N$$8;V�D��/7��� ����i�T�D���r�@f��u�+pg�8��[��ډ��w�,dm
�����|�_3���bؖ�ȵf@#��gć��/̅�-�8��'?N��l93X��.�^l�g��\��l9�q���M��cAMPx��k�9aL�H�3qy�1�L�0�fB�@
j��$
r#Z�ſXۊ"��)�߫���,ß!\��T5�b�]��L�JW6�A�b��%=��:o�����4Ϗ����5�s�ĩ�� ��N�d�̘�P�G����(1	>[�"G_�:��n�g �����Ⰹ���KV:{�iŭa!��䠽��w��n�������oX��⌝]�{W�1���d��*�-2���-���+v[۽�����#����F��gX��
��sca;�������x>���/��^oH �+þ��Zc�?���z�σ�s���WW��-�o��c28Cɠ~'NWs5P��-��΄VB�҄��D��]�U%˭_E������{�c�rA�Δ�
�nQj
Ts���Y�"k���#��~za� ����c��&	�t�G�i�<��~�/e�?#��B��k{ZB��A�|��p;a��L����g��6��|a�����r���+��/����T=���q�~a�b���zV�COIjS��x)9�$�P�0��}Z��A*�}����k^.X����%��D�D5�b�#ތ��ft�z�>1s�j�� �v����oih=?t�l�0v�D
����h	+�CYl��/M��c�����J<��T���K<���sЖ�~b�����Y~)߲�}G�?�^����=)
�:�غ�6,�UO19��ͻ�n�P��Pe���pK��A�^�K�[��
���������r0������[Ֆ�.f�ˁ�����c?��H�q!��?F������|9;���S�`ް��9ֲ�8X����8>�\^���'�i󝑪?۾������m�J|�����L�J6���������31���H����+��?ck@�]-~�^���m����x�PA�s����QQ�T]U@Tm����CR�C���������AI��!�i������������O����~��w�fs�г�����b�{:C��c�-OU��edB�4O���˟�}��&r_�����u�x�r���s�|�X�ƪ��aN:FP��:��	�5�1�F�<i_�q�F���@�ր�j
Y=\ȵ&;p߅�5�S��������D]$ @�x�K�j�Tm��#hKOgX�V�Đ\z����������B��?2f�7�B:<Ȭ����Z1��Ey�9Wq��R%~�5D�z����%��y>������V���u5�����2Q/�0_���8�����]�;��+䢏�T�nTt:D��s�R��+1g$�D�g@��������_�T�}��J��{s"�:�Q�b�_�%�ۻ6�����ȼh(K�+�F�v�������O GaY�Q����]+۽+ϖ�|���>�H|n���@�T#�4a�Tb�~q����4��,�sXN��T-���I���1N>D);��he+}(t�����&���Hф/fäC����e�R��UT�;+�+ �no
���4D��Ӎ��^Ž�E���PJ���{7)0~��َ}����K�޵2��K߮���c������O%���D�~��s#xme���v���ݦ@ğ'�X��`��~ι��r��I�={����9���r,()b��=�O��'��s�\D��wn_',r��\�|��2D-*�,{z��R􍋅���������l�����Z2�q��ψ��y�>�J��K�^Au:J46ӵ��ƅ�����~W�"��̓�Y�4~����\��%��7f��ě���W�p1�	�f���I,:�߹&�&8{lс]���LV�F�%�Ł�64ck�����"�{I�DN�����쾉��S�z�|7g)������P
�H.)Y~�$���[	p�*�B�~�]�b��,���<��of&�O''e���Q9��X�o��nX���I��N�ag3�Av��ڂ�HGֆB��K�I+��_t�ٍhqXK�MS���Ԕڨ��R�\J����VKue<��u��~��X��]����Hk��|6 ����O=��l�@a�h���,rjS�������̏�+J�'���+s��>�'p5Y�Ԡ���!O2���`-fo�A�����i����$z��5s=�uC��l��_�菔���r��
����@T����.�){��kw��}~�b沗�Cz01P��Vh�;�姕Iw��"�����~���/�7k�r�ڶ���!=�M|�,��ԍN�չ� �zj�:�K�� 6Ώ��&Pý�4������c{i�z̏���-�ڟc	��J�UF�ABPx�Z��蠠��J�����]@�x�Ͽ��k�SO�E���]�9P�����E����қ�R����N�/Lx���Я���T��@���XީH�UH��w�o�F͊v���
<��'�����a�7�0���$���|-J`9`�r�h��nܽNŹ���[ޗ�n�F���������i&n�����dG���B6]���G���ۭ�����zfШ�L�|~��+�3�=������|���X~�9���9�*w��ߋZ�O��H�W�4�&
z�z�E%W�Z_������m��/��"�+Ut|�p�(���9,i�������s�6cF���� �I����{7��~Q�~�.���dyZ����dw~�U��!t����`
N�������7O9΅����ᖟ�C*
_=e�=6|&*��4���]i��Ɇ��(2�n���;|�I_�3�|���kƊNQ������"j0�h��>�K�
�ta
� kb��xJ��������tr�Љ��;#L��[���a��G#��S�bH?aF�����d�![&��槡r�}���]t9D1(3ΩmZ4�1D�'�?b��&D��9���E�v�z��T	&�7�\�����PI��j�Պ��8�����٫�<u�v�����@H>|�~��r��닲0�9g�����:�Z��"jO��d<���L�F�d��g�%����,Z�[-����IK���,P��d�gn~E�0��W��6��D1f"wDRؗ���I�Qv�K����7����\�\�?a���X�Z�'E�����h��74ߗ����#�v�w�L�M �*������#��b�&�T���m- �� x�C�ۥ��2�I�Ȑ/Ә�������t݀��|������?+\�A���X�S�x�.7=q�B��)"]��:��B�oNB��e���]��q���o������ ��@w���nA�3ԏ¤����O��g�ww��Ƿ�B�w��ύk���&*-�P~J�d�$:�7ܳo��Ϟ��f���=�<Yܴ�a�r�Ğ��"@��z��w^�S�� �1{��?gy�1T����#'�p����r��	����P�zB�ʫ��N�����s&����kqqb$t�ͪOh)�:1��=5��?�����8]*�*ꐔ2����6�ϓ(���՘�l9�':�#���-eS}C����i9��gM> �K����k��<�1�3�(|����L�ǟ��?�Lj�l�~/x��e��D�$k�i�ڗ�S��\z^����%E����RE�E"��Z�ح�Y����]�P�����X얥��g&rW�G(|�.���2xBZ8�<���5�%��$ʊk���&����Q�u���"&ۉ���	������YMbJ��,��G�x+�P+k���S��G�ۯ��8���3�3(}/�bwؤϮl��h
���}�#�{%��M&JzV�li@�!P�$j���*�Sf�K��2���Y��t�L8�2�f8*�>��Y��`�t�`��5����b�cGO���mݩ$(ГهuۺI;�A��^ж@�����0F���Ѷ�!�=E&�T����m���K��xpr��)C@Ԕk0ַ6������*^�}j��z:|?�5{ޝ��-�M}�{R+s�ܶS� �o��/"�{�I])�,}��;�����ȻӼ b~=CR��m���a��zZ)�q��)6\�>k#�G/ܮ���]�aHƧo��ⓚk8n�H�s�������k�����y��4T�qr"� �r��9��6t�x��F�t��Dv���5Ȱ10b�q9�G�Ώ��&jZC]����6������iK��/6�ŋ�Ȯy9���H��-�]��.^��ԓ�A�;��H��Ē��yiD䔖��\��U�1f�C���:��,Ҽ�|�w�)"�?�����2D��P��tC�Q�&;ȿ�ͩdZd�M��f����1����`��n�]�i�	9C���D�בYm���6�(8�
��E�֓�B�n�dB�D����}v?L�	7̶x����L�>Q�>(���ļ4;ͷ���D�g���^زBx�]�7U\����X]A����%�&��~�Q���ԇ&�|˧�B��5���G�y�h�ؿkXNh�1�'�S���n��՝�����G
n4p����4E��l�]��gG5��ۮ*�PD�����6w��*��h���f��=+'gF�Cm�ͪx���+�P�/FZ�9  ����[g��Z�a?��OibpV,�_?�r ��*]�S��>�]2�|9���Dͧv1��g�����:]�m��� ��#�|F�L�n��:��b"�'Xp��~��n�q�(Z`+���K,wU�+���K!�4zL�Y�\����(��,�pp�;��PCV#|y��qd߼��4�	��7b�֍Y��=-�+�R��r��h#R����$~Q�)8})c��]���4�::8�Z���1%Y����qP�㟢u�d!x�J�0����$�ҵ���Z ����[�-=�`O+��s|�^��!w�c ��T�1�ݚ�汊Nb��Ԥ�5QK��h6������DD��}0$���YPkGIc�o���<9�����[����ҟk �f ��D�+�*/K5��.�Dx�-����u[���,,���J�i��kL)�'Rq��3X>�|n߃��*�}���D��h�%�<�*3���e�b��P�=Q}FG�fJ��<�a�NZuF�'Ӑhz�ֻ\ɱs!��Rw�oZ�S���j�H��05d~�����*�߈%�E�6��b~8����w3��0hM�/��^RzC�ť�k���v����2�f�4���@��g�6C%����>��f7����CL0�5{��+[�mOܭXݏ�X�^��;���őz��)�ԼIu,����ȍ���P�ؙ.M� 6�;���V���_��Vic�=�n��FvR���i��Y=�ЊB��+I���$���O�9B�X�<)�������j��_`�u¹�>)+�'����Dֈ9��'��Ab�Xwԣ�֐]����M��HAC��n�����x�GW<�6�)�8�����8��d"�K�v��&r�>��|��:F��B�5�G�#!���~��z�q��.e�[�6�t�����������-<II�u��tM������ԟ�4����hL>Ho<���db�'�T�_�6���IY�=��57�n�x-��ݳ�mQ�v-ؔ���jة�+���-��Kذ�*��������3N�?�4�L� ��s�}T@(���#����)��T�R��|ILe��}�;�O%����� ��sNJ�~��w9����#=ւ��4��^X�pA}k���W{i�P�#k�*fQ��A��@٭]�����z��Bӳ�O�ѡ#09p������+������ՠQ��0��'#_tc��Ec~ܫ�8Ҩ���UHި����h����a��R�<��L-8��*!�)hO��(M}�J�b�Bї0
apƯ����W�ƚ�L���Ԕ8�o>�w¿sm+1�d��q�����|0�
�H���׬�	�����l�"���F���E�O�c��H�p���L@�sl&� @����P������f��5֖�!T�G�R��Z��Ƶ���^-C����T��Z�}U��^l�2��Hq��������z�۝�"&�r4�G"����n��^����f3��Ft�]���v����n۝��MC����9�*O\P�p��q������֭��H�\�-�Qҽ���
�H�n����6�j����B��\�G��
�\fsG:��}\'qc�	�4�z?��J'R�S�M��{3�Aﻣ��c���u1lD#�.e
R�dq�r��<_�[�ן0�9�d��D�2a~�19ی=d$�݄�dp6~��4ˣ�؋}G��"�b�y�SZ��!R�>���ek`� �Ë0O�Ǯ�!(��y�Q,��.��Q�N���q��3�g	2�rM������ 7S�`F̽k��5������ln��R��@��}/�W��;�G�v�qqO��&N�����P˷f�����E:i�GLM~���&=߃��-s�X�i�g��.@��9�� a5� ����L$���Vyy�w�e���S�՞f2~)�F�����(�S����x��9�vO�X���D@U�&�Sg�M����d���+ ��_�Θ�Yv�TY�Z�y���������^��wj{ �?�5���,�C��T|��`�r���{-.���Y�����:yq��N$_-�^(��n�o`ﯯ�Ӣ��6S�!��@��4���E�:�^$�t�J;�f�g�����g���)6j�d ���C� ������s��U�$�O��.--�!~�6l2��8fM*���淭ٮ+pD����v�$o��Z�7�A��7����d� ���O����u�����o�l��ku5��T����G�)*B�˦zM�~x���M̃�X���Y�H�f-�M�\��eq4}��nK�(2MJ��ή�WBC����r�J�P {o���u��j�Fk�l�z�����%�l�
5��.�w�;)u�/F w�ӛ�߂S�+r`�������;Zw4�~�ͳ��?�-~cv�SI��v�!?w��0�����K����z�+Ub���vg����@��ᶣ��/�Ҷ&���p��5;�z>{*ѹ��Rp��v��=���Y�(6FX���^�������%�3��FH$��@�}�!��D��ځ!�Z���0��ծ>tey��P��FόF�ͱ���I^���qQ���Ŏn{�l~�ܟ���s��[��S4�=�[�Kd֍�1u�+����àZa�t>L�h�Z =�𡬰���f���CsǑuF�%�Qb��REr\x�>--@ r�_$�B��Bx�I����5��j�h����j&3�F~�����m
wEI^��h�R�8���9���G�0Ǟ�z��B���I�CT�ك��Wh�p��1$��u�rBlYzX�����%��I��N�M�ҏ-�ޒ?�T�(��ph��+�{b�%�׾�}JY"�ӭ��Qȱɨ�b:�"Jy�`������y9�:��n-������%�P2�'�wiu#����e�?C�_}��b��-C��	�xc�0ߍG�{K"�r����c����fR�v�����d��7z��������o`$-��K-�a�+�{ȡ��Sw� �o*p��<4�vlS�蘶�|��EеP ��8�f�}�0{	��(`k�R�2�s_DSZa��U����D�}e�1��X81|���g_~r���U� ��G��������K?q��e�����Y����at��</�ޑ&X����G���2�5�?�ͦL�R �3�X�i�/���ȟ�kT��m�����iݣ������9�g��9�٫p�
������3�h�	�k�(��������>ksԙI D��NޕNy� �ԣl���Sڣ�iS��oO���^��I:���ť޳�nq���^97y�F�T�-Ǵ�����!�
.��m�7��$pHtW��<I0!Q,(mն���2����c����i��Yx���HEPȬ�J��OOت���'9�z��B��I[0�"�ަ:��F���ƍ`�A�b��R)3S����1�{S@'����-9o����1u���~Tߩ�?�+�۬������7>~2O1�G�m�R�hT
�ufS��e�5�� _o� dd*�nS&���_wM(Yi/\����0 U��r�R���և�ׅCDB�����.@x��B����w�T]��n��(d�ī�I�(��/����g<���S���C���w���l�o�T} ���e*R�Ғ.G�/�5R�o�2 ˸ȏ����]&k�)=���;@�Xb�e��-P������N����2tP�,���r8�(|���<\]�ޅ�e�C��V�?�ރd��M��ZKB�A�N���fp�.M��P�OAX���o�S�.���̏�2��iXtk��4�L�?��]ɤ歃��LK���|�~��b�AM߷��g�'�[�ȡ'��5�e�b4|���Bw�sD�L�б�vX�L>d�4)��O�����/�����yuI��v�b�q��R��'�=�"��\�;�%��j҉�L6k�����ϓ�N�|��DC�u���W�_фW6Sc3b��-BSp�>I��-u�=���3�����!2QB�����j� k	��HF�}:�l����1�\�&/�A��SA��ayҹ��0ᖢ�8O�ƞD�o����b:��	�2*!9'�)OȹKu�y�Z���-z�\�&��y���qȁu�Tg|�EY��W>d2�}�f�ʃ�����$פ�R��>YG��$�)��f�/�����^��/�.�7�~�0&::��7�����P����O�,�u�_����`8W������	���e�I����Ӌ(�}�,�u�y�6[�(jR/؁el⺲n2]`��.n(��[�rX���L1�#���l�QL���8� ��+�5ȣ���fT���@~7�j�RH���w����M��}�,CU�i���Qr#C��Ҹ�0�r�U�Y$�j��hoN��^���:ˍ��0l�lv��x�>�S�����m��>�f���V�t��7T�	a֞�M��U�X���y��r^X2����(vI��ޛ���������$�nA:�[��(��#���k=M��y3�o]�㜽&��`�@ H�	7j�& $#��G���ϥ�Q5T�3�*7<4ø�>�<[��\o����>ћ�N~����vR�����3�0����dD��Ɣ7�9���Y��`�ƈ��z�?���Z�a�y������p��;
yc�Cz�6mg��]ȃ�2�Z�>;�^c���{�o�6d���@^GA�=O����:S�EY�
�uj��*873��y��w��/��E�I:LGԻ�m
��f"dB��K�d.� ��1V�o�C0a�*�`�U�xZa����laNB$�Js$�=0�~bt��kG��͘���hQ6�����*ښպ���S%�����~��La�ՔO[E9�S��gi_$�۩������c�t�5����ԋ�(ږ-T/oA>�F��F�l��Vۊ�O��}�5�w�����^|��̤��W��TEly#���M�ze�(�Zz�|�#�+Fa����q��1v������m�:']&���E�=y>h���@�Y��.~�=�~Kf�͵���"}��֘��n�|Q���-�̈�6��?���[R%��3�'�a���\���4|~��܅zp�X���	<_���{��g�'�A�%�]9�:/5�?��!�k�Z'm�Y�. ,�oY�A�{��p�����a�a�f�S�hL������;1�a����&J����lc0'�`Q��X�j��b�Ʒ�V��H>�'.ϑ지������4���\����e���7U���̞� l ;�YbJ0-�Pp3!�þfJ� ��l���X$B�0�HHq40�}=*5��m�|$���o�;��߫
��KJ��&�q��/!+�\�ֳQ���84^l�i@��W�[�Fo_�z�6Z����$���o��&~���T,<�M�O?����o��zM�R��@WT����cOO"�{1�Q�=��O�۸��J������S���������ݬ:�Vf� �3�M[̷Ƙ��Cb�;��~]ޔ]��yM�3�fE��IT]|�뢨�C��c�����'<��}v�S+~&$� �g�)/����a�����������~�NbT%w��*kg0����7�pb�fx������x/�=� %��i��O�\^Ɉ�w]7ެ*+=a�(q�~Wy����w"O)�:Z��-Bc�s$�Ʌa�����+�+�b�Nq����e��zE�g��p����]+����c� �)QЏ�X��U�\!��_#��Jx����I�`/%����P��{2-�J�:������K>`[Ej4��=���{���_!���{J��kQ�o6�ys�o�¼}�lT�&<I'���^��=���IK�%�X���8�ҍ9��&R]��1��>�'[�&n�殆=W_�ݾ��S���h�넪��j_�	��~���Ѵ$���`	m�$��t��[��B�ۥŭ���ē�́����F'�DvW�bD	A+��� �U�5���*��T�������-�N��+�֥����6��;�H��<TΎ���{|�n+�$�g*��o\�J����?Mu�3!��8p��<�L��	BOM q��bM���.L���M�_/!�Ke�q��,��b ��xӶ� ��E֢�Sc�R�Qn��M4�Ey�_��d\g���h��Z�֚�;9�_��S��� ��C�8��P��F_(_ �/��֝�k=�z�R�Y
���>6q�)#v��nt��Kzyw9�󓓂�d��L��������$�_�ю� r�L�j��$9����t����[���Oԕ��q�"I�'��$��	^]�z�E��3�\����s뾃v� J���v�4���?
�Tv0��q;���͇��d��S�'���'�[lH~��Ɇ��H�zH�5�,�?�U����z��E�����ʐ����kwi�A �; �/��;ϔs%�ȥ�‧X���7�l�DD��j�3��Q:�<������R�r� ���{ި�p;�/P1pF��x�g.s`G�6=G]��<Ą���SP��d�p`~�J�8�)�c,�sj�	�~�!�k����n���(נ�&mz���f��n�N�Y����
@q�N	����T�۹���:'S��A�P?z
X$b	�ȑ��i�8������MU4��5ݨ'�g�dhpN�"��iPP-�Vrܢ'��8,
XΊ)�\,҈W$;�>�ql}�fB��8�l����<1���ڭ��a�p'@�鷣��'��a�(��Y�����y�z������"*�^�t��\˲Daw�B'ʀuaEYԃ<��f��	ȳ�?*�B9 9Cb���\B�RV��rЉ��d�3OD4�����Ɠ�I�$�:\���\h���'�)��?���Z-�7�b��M�ϓ}׌z�V����a���T!֓�P����ڤz�����oJ4R��%����N9�vN��8v�d�����v�U9^�v:�*�Ю�+Ժd�Ra���_�т��zmS� �D{�$����$���Ⅾg���Qj�������5��q ��o�0�������@U�E�#��C����q"=W#��[��Z�A�ژ��$&[dS rF�ͫv|��O*Q"����{.�
ު4�۟��Ɨ7���k?�;`��楣���BE+��GZ��0�^wd'��Y�N� >�.fr1;�����5/ߪu�|�,�e�|��WV�`��<�j(��q�!H����HVq�;
�V�oӱ�Y��>f�^38|���u����Te��]N�2@4r�9�m�]%�C�2^'v�H��X���
C�lev�����şn��є�����c���i���G䨦�"�7���~�6�7+sX��wԍ����\���`����2x��b����*��,�]�1_��s��6�f���f�7�,�$NF6L;�ۀ!S�
و������p~ 7����:v�ǊG������J�3�^!�MΛR��J�2J}���̎�tϝWAʂ�'#?TC�U����&1j`xK�݉	I��.�^�5�'��1�x�ƙٟ�xBj h��LO�&��
�p�O�鲂��tMM^�����d�X����ݧ�$�cN���8iF��}�lo��F�;�`_kM�%є��%u u�-�W�� ��Z��/YCT;3v4�Q2��.L�5S�ɵ����zV���
��ta�{��1�v���qy�N&��Ipke��Ymly�/8F��A�أ� ���h����o�t�K��",dʯC���w����P��)F��e"��R�2���֨�њ����o���g-��h~"z�\��/�w�����D �:��]w.��!��h�4������F�ԃ��I��,.�v<��|��C�[��7ܰ>,��[a��S�����a`XS��;hyb�/�~ 7��> �V����捱�<��぀����հ幝	�%����B1���t�K� �<<�z��oo;��ǅ�:a'k�i��z���$��d�s�Ї�����>��~����Eڡ^�]~��0N�;4q�����l���=������Ny�GSҍ�4^�S�NP�Ҥ6��d��ۭ,kW����;���1��S��"�V  ������\��8���*�c� �O�������~�����
�fz�2�-Q{d�Rm%�������y�������i�t}���	�!fG������c���o�!h�F�|*�`��+\���aܳ��K���:�㸷Clq"�u���`Mv�uo��/f�}�ܺ˓��+I��u�/Y*�(b��ȯ��mf�W�إ{G+ �����F?8���������τL��g�'Qoçݻ(���V���%Zo@�u�|�b��T�;8����j8z���J�bς(+g��G�V3;a?�ʛ���|R-�z-/}��p�8g�֛��*��ۑX��v}��-�7.OG�iJ��E�^�w�����w�䒂��ں������
r�kp�9*פr$hoK�~)fŷ����c)IAk�{m*�����2�1Y�'U�,qi��Ǵ�J�j_͹��~h�<f��3~���߼��-����ʢ�3z\�ڛ팷�|�=�����&�J���e�<�~5�x��%y��Z/Oǂ�ء���ƿ�i/�PJ.�P�uM��kSQ��[#5m�����V��$��'"���ǳ�T��c��ZWv��)U�e�.UW���Xao�Bg^�ba��J�I�����v��@��*��-���7���i
I��ҠDG�=�_��*����k0��R����/ˡ������ͥ�I���lnıI7��(����Z^�W��qϻ�g���XF���|�91��X2l�%�0�"�_��F"��pɎf/����E����X&�D�~�}�����_�RN��C�����h�� ��Hh�Pu�Kƫ�I*�Bu�����|��b����3�v�6�n5�ʛ��]z� ����&�n8�G�I�[:��5ng��(��/Ă�՚BÅrN�~��O��B��}y��d�B�R]��u��կ�|G�p a�$�>o��ᘣ_��q	�*���wk����jO�!�a9�u���\�������5D�E���
b#�u@��1,��� >������k�\9髾��Q�<��/�V�ɘn���%��6>�P�a&��wk�~��;�Z�X{�9q7�����w;a��D'�
�	h|C��*Z���ݼH�aSc/�;���x͝v�.�3������)x�u�So1.�a?��yG�鹪E��,;L����`!/3��n�ҋVd�XOk�?E�F�Jb��K��5��]J`8�����a���Z
L'�T���F]���q)�oj�q��}O��$5kf!�����vC�ю~���iB��c��jV3щ��HŞ������*��\m�P]�O��H=~|�p{
�ۙb\�Ĭ�?�q��b�F�8�� y<)-���m��� ;I���� ��g��{��}�xY�0��t���³�	^�}h,��`�Jd\�Й��d��h����/����>��	�W����bX��k��e�c7�͎����*x�8V2kz#�X��X#Y���掱�ʬg	q�%[��yQ��t�
Gm�s��MC�c6b�MІq�y|7�#�:��Ö$����wp%�~hW v��a���r�E�+�?�D�����(�Є��^�$�樼"�"�M�m�Lgע?�q��dw1!4l�q,��tp�dS��N�c?�������g��~��������Wِ-��M��d0�������]*NQ��9�[Mt')�O27����N�F�6b��/�e�� �3�D���!gH�Q�x^���r���@/��T~����Eq���I!�<IR1z���$4��|�7�Ri�&�X|E��Q?%����[$T���/a1�*B:��e0���;�����w��a�D�І�]Rޞ�3;�Q���K�O���c����R��1@yJn�c���_�tD�qfBno��G~v;�CM��m���h㴿!c�r�Bgo�$����$�WM'urx���bfsެ��;�EςOeE�:�F�Ra�֞a�gA�"RO'��Wo{*��[&m�F�p}�)�_	�y(^W��.� �H�Z�ԯc�)��QI�Ec)Q�,�2��k�TҎ�ym�T#�Aw�q�O����'��k��h�de~����������1W�%`'X~d��{Z2��zץ�Iv�Tdt��w��tc���c;D�'�2���D�����1�8!r�=�
Bհ9����2w�CD=;���+�@��?�&'�Z^�ꍍ 4��-Si!��o��\�'����AH lVh���¦��LŰX�|�M�G�P�*�|�1�p�V�>�R6㉃��4�;#�P�u�p�P�Aco�f��m��n�]��6�2��ۋ��4_�����yg8T
���ho�^I�&���<�C��َ�$�-K˰���ݳڽ��^M�e:����A�-L��*x����E�N�<�ۉ���ՙ./|Cq^�l����7S�BKq-�B�^+���~��>7V�'�Lb���D[�0Ა��P��2�_��ڬ���?lE2��?�g�~���)i�\IqT%�]F�<��3���s�J z`���U�M��J�WD���Sp�e	MFЊ�om��c�G�����y�cϝ텨+��S��s�ݼ��(Y��R�we*�3�Їf��*q���yMOҜ��(] ����@��j�7y��v����]�[�ʇj6�q�)�/Lچ��֒	r���Ře�}C�#&�U���0����U�t�<sP�d�w�"}<�V�������lx7E�e�۩�$�l�g���ֱWD"Z�$��t��%DՓԊz�%�;h%K�M;d}�k��5�ݎ��:��E4XN��~�M�����B���#�g[�Ȼ��'�!ٿ��>+�ѕ~b���@���3'�x��w�q���Z_s����?&�~Ys�>#� �	���T�U�2�䆽���1Aq.[>[hI�q�W��O@�
f�
�(��\��K��QLf�P����0$#0�q�ur[��iZ@�jB%�P����%��e�ڟ'Q��va�Nt�4S��Z(,�q��w�}{L/��������ۆ��Gr��/�{u��'��P�.?V��ŭ�J4EDG\�g�NUU�1(��F{]���$���d�A�m당  FgUx���Uj&'-<��M!~ko~`�M��"%��ʹ��aQ�G����
�]�f�Z�����0f�x�Uq���ր��ں�q�=d�BʆF���r�e�1:F�;Z$s�AS7��?}�Z�\O�{ (�=��qkל��4��o2����ŵLiNgn~��1zr"H���(T��~�S��d!~�g��kC��^b[nd����C��e�k�v��v{��Ө`r�3Т��Vr�;�h��v�Nu�7ׅr����Ho�c�<�} ���.�M�M>�L�᭑=�<غ�){��wЏE��9^�����k�'�r/Z�����A�C��d���"-C�IX�	aG��-��DK�y5�!��.�#���$$[-i�~,�����6o��&%�;c 	����fn$�iy�;�>�5x�k�Ya��	bh���ɦ��&�\k窾�$BQĿҨ�p��B �tho-P���>,v4�z�w�����g�>G�S��r0���uK� ���q���L���t����g6�0���:q Ӡ��k��*�B>"�I|��[GK*�6�
�T�Z��u\��Kf�Twi�7�d��O�F���>ɌŝW�Xbۧvd�����٨�����Z-$n�2
�
-h�3s���{�8	-޽�~�ԙ�D2nz@���iP�eglS����erf�����߷HID釪MR�u�ʙąj�Ue�0���Е�Q8A��ᯧĩ��8j�̏�/�{Q8�&[���(N�� ����J�i�������0�͛�	��?}���Yn�fn��}�x���&�/D�M��.$��|(�e��*6���d3@�E���m&U��(^���y{"�-��'}����fJ��T���U��H*l�kc�gʸtE��u���)��l#I��`M�_��m�!�^����1j,#Sˌyhϕz����r��cq2�SgY����S�+�}�y�P,�Ư�.�r+����k !=`�<k�r�W�-�M�O��[�ڐ�Z:���*�*bV6z	�F��~zo��Bg��N���#�4���0�q-�Lx���G�UV�'>�t�R"�up�&3�r���q�����y��o����f�t�z�	w�;
rs�t��|?ݙ7��*n�i�Q����G*=�0��e��d�=�z����s�Z�7+�|�W%��ۢ+%������I���������� ��)ZD�Ԕ0X �C�	���j6�S4~#�wn���j�������#�BJ,!V� Uܧ�5��|U.�â�-G!�K��W�F�єTC�f���
�͐?����Re��J˓:R���/��=�_��J���v���b�Y���ktaա��q��xd�+#7�tm�K"��1c�����h�����7��@+���o��,���C�R{�|^�lo��=��]_3�Z�����1��������T˞�<x7�(���Ёێ��u�dfWk(q�Tk�Y�	�w�ʴ���
����q�1�1t�\�L�"z�<�{n��6J��'�8�1�n�ǝk�`ŅÔ6>�I7�Wz^���XƯi�WnP�Ns�G��F3�1X`��k�9_�l
V�L2%.�������K���6-B�p��/l���@���c�fJ�Dn|;7N!=���Q��R�Xp$��2fͅ>�� lbg$��33��nx������q�8��Y!���P��aqF;�0�Zlp+V�]
EZ�;C����Cwww��������GO�y�~�3�M�W�V������}��3-���������R��k�@/d�N�DLwE�͈H�sx�����·�l̚�t�L򥋷�4��Q�<��I�g>_w!I����BE[���|ڦ���c Ї��rA�́�����I\����Ϛ�PH��֮]����Ӂ&��`n3�w���E!1H���1� ���#�\ ��`7�S��+E��c��Q�h����.�E�M�����fs�=�-r'B���s3>˼$ȓ�BB!����ܻ��Y�j/o?�Ԉ���ëٷ:	h��+�<���2Yr�5��Y?�n3>���p2A��}z�>K!Pv����&��Z�sH&h�@3��+WV���'�؅�rC�W4ƻ�<�.��j��A)��a�#њ�~�u-R���/�Vt-��9u�\�kk#�?�/m͕�Np�-F v>i�o&�`X�	����c�@�d�yrԱ������Z�����d�-�:�k�w��j^��	��c����'�����f�\�ȿ���h?����{�d��~�k+���G�'��� ��\Hl?wW��r J�#=�K��4�iH"[���~���؝q�fOe��
�����ŗ��b�)um���ڗt[�`{�oڱ�$!��'K����Oa��a�{�d���#������.,�*+��q�1���(�~���(�t�E\�T��S}A,K��ނ�JR���;�PC��;�z�uR�n���]�!�N߮�-��	C������J�c��Y�[k��	�	�����%/}2�Ivde�'o�ߠ����/Y�>�)4޲�~�9�bNt� �K�v�#���<WK�F�z�o��C���z$}��|�R�FͿ����_sq�y���].d�}[�]�נ�@�ƣ�/���pO��F�-Vr~
#�j�/��c����2pSз�����*��5��mI��j�(�j+$���
�'1����U9�?Y��	9�����r�u_�<�~
���� �u<�ѻb�?�pޣ�/@`�qB��s��f:m��q|4�t��EF���?���CL�j���lBn� ��煉��+ټEL��F���ű���2lA��G��$t��j����o`�eSӠ��a�N AW6�ݘ$Q�U�a�S~~�&X@I3���=F��ǩ���]��$���ֶb��������[>����~ֳķ�pxN7=�ꟙ�]�;�j�
7���Q�����P��|�I�gH��Z&��x��u�� �,�1��z��U,��;��(R�à��_�M{J��s��?�/�̣u�,Ϥ���l�7��窌LA��q�S��55�_��3B��y�.( B�DMBk�B�-YC}Q�D�>��e�V6 �uI�0�i����9���Tm0iY�	FO��������t�W|�VW2:����@�F�3�B�ˎ�r|\\��[{�����=l�;J���@�=����zM�v�;�+��-�w< >�����n�fW�(aS�����N��2�C�_�i�� �;�"۵���tz�9�(�PX8�)m��E1��݃1ǆ)��,!��F/D�s-���tE��6���'g���O�$�����X?��=}��/-S��#��E�����o'�:��N�ƣ�k��"�ɟ�6A(_#��_��0�.ӘŁ���39��@oƩ���;��]}x�D�Ӽ\�'����Tp��M��F���n!��uO,���}Q%k�2UQ9�P��%���0��;nRp����ًQYg�5�& �ϣή`�p��,񴲁����'�0�S}��B)ť���t-�� �> *!cqF�k@Z��IU�+ec���X�fї�@���`��]�k��[��Ef
���!��a��ܒ��x����4b�b��N����[\I�~��\�����g>�ցd��� �"k���>9�Q�$X�oK��HM��nD.�3��_@�߳� ���x�ĳq�bo�"!�rjXƌY�GC$��*}��2Fً���\b(/&��F�7 `0F'�A�l���}L>:d7h�Z(@�4S)Q���0r�kz �PM|���a��}�T0�J2~"�Q����95v���t���]�J����i���7�A�|�so��d���|fIg�)�|�0S����.�ۙi��We�si=$	\��.�]B� Psq��4�Up�u	ZO�7�I��5�C{�{��1NK�v�+�m����2OR:�
���:cÝ�K�;A �:a�/�Z6�Eip��Iu�C��r&�+��.�Z�O*��Fܘ�v�o�,l��N�oO�F>�̀Y�v�*�����Zk�&��!^._�����P�����ۜ�3O7 ��w�ڡ�}{s�_�;�������Q��I���Y�IHŬ$X�l"V����RϺ�k%:�?�x+8־[93������H�Ӕ�?
��ۮ��e7���d��gv������d��?��jD�dI���rs��2���� � _��h��i|bn����ߞԽ�J}A�W0?�ۣ0f��i�.��@ӥ4P _��X��r)�)��$�%ej�w�}��%��l�1���R��S}��T;�s��-�i���1Z�Jf�� |�����#Z;JC�Ь[����Ӎ[��`���y��p�<뗻2�����M�<9Q3mW13�,§��*fN�'���T����� [6l��$��o\�әdJ�$���h�L�j"�)����c��J��_��V����C�	�Q6RX�?�<��
^1PS��3��}�˕+<e�w��^G�@��i�Ћؙ��G�����΂P��-�O��dd����_�	���=��qI�CU��㾵0z��ǒ�Qx#��u$䐷`6���&��/�UW�/�mE��:�^��	����F��$W93i0�0{txND����DOL�%		�q�������1�Q���Q�M=4�������#�11�p�y�!A1�T�ݶ��]�b�.��+���ƍ]�J�o�P��bC��l����]-!B$�{�_��~WWpٞ��
�vG4~-�<��C��Gy��.�sk��P�IP�IL�!��U��	:}��3�=�'h��t��6�lj� ��u<KE��4X5��c5�[ǆ#�u_��Fz��c"��,�u�h9֭4�M~#J�f�<�@ғh���iij´K�)ژ@�'���:ͬ�j"���]�ԋ ��*׹��-��f�ȯ	)��q��w�t���_P�:߯�=�?���ܚ��4-��I"�e�%�������u蚤�֟��݃o��N�ͶC�#8��}�J�x����A%.�Bt��Eױ�xy$g���;Ջ�%a���h�`A���$�i¨
���>�=�;��{m>$w���D�^p�,��͚��z��*�/w��w]�\��r�Ӿ�Z\�s1��Kw�x�q~nQ�#�<��uc#'���A=Cj�{?�0p����@1�aʰ�3a[؜���?R[�r��)�w2�8�n̕��D@�j2����BA�6+����f���/WY�����)��T�G�4�$X�叄b��
	�[����J`��H]�~*���` �|^�-����II�)r�h����a�����*&j���p�k���� J�&��í��n�P�Ŋ^�
7�����WʰW����#�4�${�Q�� ��������-s��*�]V�.YO�!}�H 4"�<˵I�/�_�k������O��O�뢥�/:&�QI�1��(���Y'�E_���"SL����3���7��/�b@xF�C���H��!ˋ3-O<�����g��!��+b���)l3o1g�rv�Isqn-� 
����T����:v�F�okɟ��J�ӶS�3�q�@��Du\���:��AN�r��5����L�~#Q�΂r���}3�вc�����Y/�V�Iq���j�؊2YH��o��tUo��=	�3�=��������@'T�����M���I�شB��Db��µ{�$b�<�(̾�?Z��[��\}��X��鞓/�qMQ#YJ7o/ ��Y�n �8��M���ei?t	'�цT�������n1{c,o-n	W��ف�����5�a�Xkc}���"/��;���$lF˓����H����Cͯ'c�Z��7v�$�a�'"\58����{e��9H��jm�ܢ3���p�+2=��RG'�f��-�/��JQO��}*��c�m��嗪So�ۿ�������ly����2�%L>���g.���Y6��x��*�!��_� �̫����y3��)�=|�
L�imR��/�$B�v�Wò�;_����0��޸A�p�w]�]'�}��O(����{?�Ȋ'�y�e4��W��((໣'�GB+t�'�\�e���U��՞��0\���2O6��!���?��-����w���~yr\[ՆUH��~�k^Zf��S���6[]�2QH�@�ҟ�{\жf�i�z�� C�{��[�1�̡m�d�C1�j�y-�u]���Ϊ���ʪ# �G�	������@��Ś���}� ?�J!��<I����6iղ�BB;�~�Ӣ*�B0�U� �L�����o�){,4�ϳj�S�QB���9��F�@Yz[c��	�R����¢�O��!|��7O�^;�����qa�����z��{d)_�x����tg�,'�z�|����QO!�/��e��D���EjX��y*`m`�R�nZ+�ￇ��k�6v'�È}���FW"H�P:p���B�~��&�{Ҡ�4S��߉���6�h�m��I�ı�5�=��,o�m�%����b�Ҹ.��\��ƿq�C4$�T��#���w1{B��.�	�a��hQ-/���9���1�/Xn�L��%m֭mmTU@�|�z�w-|_���� ���'>�ې�1r��ل���mj<Sn���t,})zL��$�G��
RӄT�]r��wq�+�	��.����p���CN���;q��������~�eC�i�|O��L������u��О���������߆1��T�)�;��7ZB�V�.|vh��XG��n \����M�aS���_&D�����"t���IBV<�F��7ֵr��7B���e{}��|0v�7�|�;&ɯIt���6��ѣ���ۏ�b���	�%��������#C��7w�QqX鏯��fa~�ӗS������*��R��=�m^L�vt�;���G���� o��.�_E��ql`��^��ߎ2ԛb�w�2{JY�6��+4ѹ��p0��9�h�o���gx��BE؁��v}�hJ�5��������b'�pt�U�[ �J��lx��A�Q��]5[�"\�!�ϩ<"������q���6v;Tk�5���
+�Ʋ6��-��﹃��:���m�ut��v�u����+���^�$w���_^�#���p_^�Vg�/^$�m��i.6K����"�}��<���ϱH��D�����@g�~�湾���Z�y���@N�J�ˢ���4�n��f�;T�t�E�W���3�g��o��d4w#.O�!���R(���n'(5��B+x)H�� � �i	^}�J;�J�;7�����gUbSk�y�`�8�?��K@�VHE�y�0,|��h���9mP{�7�6��ZT�� !">j<	���a�Qɡm��a�����^�}c�/�ۢ�����%���~5���Wvlo���ǟo�L>l�<=���H�\%����!�!zn2�(�����{�BB�[i&�z޷�c=����ч4*�r��o�Nv��$����Hd�X�V:�T�e����6����i�k��z�g<����@�Վ
ы� ��t�bz��!-��֐���x��������H�W4��>ߎ�'�iϠ$����
�x����ϾL9��l�o|D/s�d�&vF��ItP!<�4�˽���/f���hʛ#��1	���pKeJ��z��R�lv�Ʈ��~���u�[�3eY�lv*���ʟ��U6;�^G�`��bvnE4=l�XB/ҁ���b
������$��[����1`�����˖�`�g�?A<�����q~q��0�wG�x׼Z}?S�\�0W91i^\��Gu��D�ٝ�+yO�MXb�衐M��V���i~�!�;5�a/!�|�c��֪���V����a�&���C���;J:���U�����O!�;��<�0qv;s!�J<�ٖ�t�����1������'��=�P:�q����_��B.����Õ��q�i�yw��]H�,�4��KA��?N�BkzLl2���9D�	w��cx���GK��~P�%
WL5�s�����A8�aDI#��>��?�x��=τ�c�;-����!R��N�S)u6�Oց�y�$��f�wS��g�s��n@׷��a��H^CΰhUW�<��(O�{]�f���~1�����$^�##������y8x�����_�'�HX�� >*ĳ�`�fE#��^��fm&��U���s�	��^.B�`ذWmI;��J�:I��JW������<'�mm����@}�`n�7^3���Z������H�ۉW���kX����;I'EhKq5���c���g>En4�p=�3��U�R�<9���tI�/]O�~�E{烩�(�ػ�x]�n��������T<=�[��z�����(�����[y� X���L�l2��/��H�E��i^,�w�9FHTu���f��)7� � LT��|*ڹ�	�!X�ra�H�� �Xj�Gx�)��.�5YG�a�,�)`��9��wq�b-N����9pc�3(�j����n!F�V�w/� {Sp����i�ߜ���ea��v�W�6Y�~��*�ľ��{�F�2�yY��`ʜ��gC�\��������]4Z̪;��b�"�D�g����}��7���H���h�T���&*�[���S�@u+K+�]�I7b����Vh%�&��=����EƟ��Mw
k,��z��.U�v�2�^7���ĨO'��h���-���e�)�8zX2�t0g�1��疼@P/�h�(�>|�w��:���t��gL��h�R���q�'���V���0���4�t[Amϫ^�D��I��a�HME,���Cg��<�׃�����}0�������7xi�Y1�F4&�68�G�A�3n��P��W�wo���}T�w̄*�@�o�����F�qQ{r
��� P'��e[��m�q�S���� i�هZ_Pg�9SN���?�j�e����WԈ��3fߵ�ki�&�i������8lI,��m��!�S��ߝຬ��;ν+ɩ%��pr2�o\�*$\j~�ǠBΊ0��6^�q��'�2�C���Q�,�%A5uv�3�eyԝT��Ҫ!���{�q�^��������@1[$ؓZH�x�&b�z���.�zi�sg����P���В�����~��oh�e�Y".���gB&�\���N���㠦�Im�����B��Y�Z:�1��s�X�|?��-ݡ�������}L�D���\��#|�����%�Ҿ�I��CQ:�FC�Rm�= +��"ȝge�9qh<���>i�F{�h&V����؈3k!V�����.��uqDh�_��$M���d���9₃;0_��1�E�t�7x�*r'�z������,(�N���(�8�b1�?V���Ɣ���Bv��s �o��C��*K%��X��=�a�Gfdr�ئ��w�LD������h���ͽ�MmH�
��;���h�>�}��1��iF�U���u��3�,+y�yN����>Um�v����k�~��**C�쫞�uk˟��>�+�
#���^{x��֌�?�? �v����З�YV:�N�e<�Q�=�3|����	a(�sofNb�R>�k[�T6+}���39�1ţ���i��pB�[�ëo{@7);�͍/!f.�BI�Ġm=��Q;Ξg �>�ub�;������N�<A��!W��PkS1 ��D�[<6k,i-")KT���`XΆ�[�� o���A�ҹ�5���zy�tJ����#^���b�
B������&?��^;q5��z�0~����AD�u���p|�D��C���,K� ��ɒp�����柏8ܺ�uR�݂֬��"�Ncf��Q�TF �h���,��[�'�v@�YY6��N���G���ZM�^�^GF�6�DZ�';K��Fw��,�K�����7j��Rݬ�dk�=�ݰ�6ȯ���Ή�I��-��9{|��Az��@��}$=�)��).��ziv4���o�x\��4�;N�)TОu;ʝl��$'����3�A[n��k��?�,�uܵ�^?��\��+���W���өҐ������?a����!���$-�LdfiV�����Z	q$�d�s��!M��bX5����}�"W���N\��=O���ʐ��oM�D5�Zg�8�<���pyv�u�q��d�}��:����a��Np(�ԍ�=��ܞY��&D�} ��D�8JO;:���/�p���n�����8&^��%B���A?��|���G|7nLC@u�OR�������� �|`�a�}D��a��|]MOo����EWw��z�������x�����X��;l��7x+��g-���Ζ�ۮMZ�7.L]�u�5ސ�+w�Jr��$�:/���zBʽ��ug���*$���o"aԷ�Ѧ�r�3�N2�6�x�}D����=������\�`�Kex��NF��LG�o�����L�lT(�i��������Vd��w5h�����������[Is
V��A󕩩�����'��*X�O�n�����������⤞�ōxD��[��z�YNXx��\#�G�����	�}�Ybٽ���[�M��̐��c�W���fMt�:	]��q����\�D�iB �-MAa��rR�ܧ�`U9���k>7WKU~f{�q����7�f���J�M�l�/d^,��jQ2�z�<ӛ �� �k��Ç� ���x�췪2�W��ҍ?n����xm!]̺9Y|ms�T�<A��$����?��u�[�U��-�fϊ�Q����]Y�������b����:Q|S
����%�����)^p�?J���O�Z�Y��vfh�*����Y/�:��Yi��Q����<�rrA�RN�tI%'՜9��ѹG���~�&5��+����)�E. �'�$�u#Z��U�'{Uw�?[�±"�9�00�f������H�6��^b�+���Yϭ��T1��d����2�)�Nˎ�o6+vbN�'�|�Cz(�F ط�lz��s|i�̰�8��r�����7��keK�Ѫ��b��+�+sW��-;�UK�n)P���S!�\8ɡܢa�R�X�\8y�8*AȜ����Rf��4/_��"��ۧD�d='?7k��|y�Y�I���<h������qs��������3k�����u�Y�R���<)e���x s86& S���`��}�~r�ˏ��9����V�M)i4���/_e! �Q:+3^������r*��>}�����yy2�2��9�T@y: �h��sS��㶡U��/5g�,.�4�2�m��_�.6��kZ�<�x����ts뿧��RL#஼�/m!�N]
"���w����b�)�_�Ұ573��^���.i�o�^��ܪR�CGU���@���>WOڵޜ5��z:p<����)40�4R[yW�I�d�$-2q��gu7�3=.� ͸�� ��8��-��Ί*��gQ�V�3��0t���q:'���s�Jn�E=Meјpu�$v�����b����k����˘��W.ٶ��hv�u�?e���9E;%k�0J�ѹ�	���z���"�_�$-?��a��dZi@��x_>�=��o\���Wq���ހ��}�~��\<�����m���HM�t��'$KG���⾔>..v,-n�<w�+�I3�||�D=%����'�vŲY��� a&�<�:l�-,$��~�ؚxm�v��"�?�	N!L�/[Tj|w8	nq+Q��ɭ�JK���ķbS��-�}bv��@��Bզ�G�]�ֹ���ڟ��T�[*�"ʾ|p*��)ek�*pX�:��g�w��u�T8+|U��<��W�DU^Z�x�W�T��B�	������=����L*��w��<��{�f�|c�N�_h33>�K��  'A+V��-ˀ��p���_y���9b�/4g�H@����^V�#��F�푲�dG��s@&'�Ҋ��`n#���%�c��yw�哟��2D��dܵ�$S�B�;r�j�|=�Sf��������k�s5p!ǭ�m�딹s���_V����C�����:d'��-������A����8=��mD&TC#�j(�ݒ�-�[K����7�հ�a���0x�_rޫl��b��g����#�ٍ��q���=^v�l ��\��xlff��v]��3�`�����3E6O _S~-U����p�� \�
F�����5�~�c$h[d���#�vn:y��aʴhW�|�*���!4� 	���K��������i�`����;�_�b�����g� F�GT{��+���V����k�V�W�e�<��a�Mt���RU��˛nj���^@Ҟ:b� ���;�POs���b~�/�)�:���.|�9w;hN1�J���$���\z/�rsR�zq�v��>y�j%�7�?<wG��9�p
���L���GJ���л�6�t9!�I�-R/�������_J��}�����Qչ^�Mq�Z>cc��Tz�2X,X�r?���� x�����!�
�ٜ� @�{��,נ;Ѩ0S�`��3R�ǟ <i.�[����>���hV�M��&��8�7����k���
q�6T����K?���h)K�q���$�:-n+, ��M�Bre��S��Y��M���d>�B	�
��ѵ�.�����,P���ǧ%�=OR�g��������->������o��-ll+�䏳��W8��7,f�c^�0�#_L;ef=��mP�l">T�wi#Ɣ�0+�G���؀�QZ�%U.6�z�T�6%@�w<�)>c*���n�}��_�'��,2����������K^uXQ&Y�zO=�_�A`=9�}v��_�xǵ��P>d���㪇+V��)|Ӹ�Ċ'�)OE���ֺRB���4�Ψ�����n<��I��UIBob����3����B��YvW�)�h�真���0#2\H_^&%yl���PH�����齣�t�M>����k�I�}���}=c���e!����i�ĝ���Ȅ�+sa��YKx��o8�O���Ĵg��.�Z�~x��[-p'%e�-��(�5	$���>��%�-Y̺�����r����Ǹ~�/5ʳ�*���-˞Փ����Y��1�Qڝp����/	�� r��7��xX>wz��/<ohl_�=mL4p׺=���{�>;���T]�P�
�"�	��t��~~'<`�x< �3��Jh�,-��y��O�y9@s�h=O�yB k��_�'����ʹw�hʏ�]��f.�4�7�Wn`�WY5�Ih��M|�͕(�+�zF:kud��@��ï"��R�3��\�0<�'Fm����LR�2�����e�tx�~��6.���Nh�tS�*���֫l�J+�����ʊR���I;�`� ��~�XM��ܦ��׹&��1�:���a�|I
&q�u�ʯ���˔��*��2��I�/;*�据4Q�K�oׄ߰9�D�bb�.)�Y�am\��W�]�*1� ��,��#k�nt��PQJrSѕ�,DTB��F�5n�8~\bc4�K���\�|_����.�1�^SՕ
{�V覕7l��B Ip��k�{O\����9������D��A�%I��tp�S��~�c!W�.C�����8
�k}c�������ʄ�GCmc�r��a�W;�T�<*����ɇڑ3��{���4��$@2�G^}�/�o�rC���\����w��������̨������ifH��n��c���!�����c�؁n�+/���d�j�;I����W׭~l�1�Yr8~�xBtY{�03χ�\��Q�m�2���:�؟3��H,�J����Wæ7�rl�3,�1#��w���du��=1w��^���B��;��
�/���|�7�6tЕFL�\�?n�X'�/��ar��Ú�B�_�ᅢ���7+c�����YS������%���ͦ=���VJ�D:�G1�����w쓬6�* ����S��q ]�M�$��&d<�R?��Ǹ}��h>�6B!����Z������s[;H4p�I��������}VF"�λ,l���0t�-���Ď(8�����>�buO/����H���v��iE��KKW�1C.>�X��}�Ґ|g�99 �����-�8���� V�����sl�?��n�Wn��Q��vd`�l�$�<���ۍ�g�R�EU�$T�a}+�ۦ?�U�veH��ΞF$��V=i��$��y�2C]5��)У�f�%��A�,���y��0Z�b�
'�r���0� ��U͸��׶��Ԕ�#�� �WP>�k����1�<{�T
��޽E�����(���8I��#��uD7+���%z����Y(V��[��ę�1 5��l�%ǅ�1ۜ	�cگx��ŕ������]�PFȷ�&o^�e�]F�=��md�K�\	�vÇˎ!њ1��  ���	ή/%�	{�:ө���o[٢Sٴ"}�1A�T���cب�Q��[����]Am�+关h�"_�4$;�=�܅�H��+��}����=a��h��k����ܣ�:�H��<��3�,8�k?6?F��9rו*zA�˔���������7w
r��\Q�]g,YK��'w��߭��<Β���,4������&��)8�B�=>��˷�ܜ"��n��2��I02��~tq�g�{��i6�.C�*��f�x�d��w���F��J��r���VC�r�[[�n�`AKc;�����dw�
�c�1t�jU��'<cQ�mm[�8�G��  g���M;L����|�O��c�Bݣ�����|���Gx�#�?���G�&�������#�"��~ 8+v���붌��̐�+>*���|ܬ��`��׍�w����x�A��j*������n̲+�B�s�?���k�߾6D{��hd�0Y���5Jbz�A+��k4b7��IĊA&�5(~��i�R���2P{��N\ݝ�t�Oh�0	kr��$�	Z�ΒOt�
V���d�Ub,I�������Zʖ����Ax����X�E��ญ�@7}ƀ�x�W!�&�^|���Rp�\�������A�#���e߹���u��I�@_�H.��d�x�asJ�OQ�	�=x�*%~Uo�O�kN@�>J�E� �����,��6����R��ܰ����%�c� ���6�x:��"d�L�h�⤈��W<�J��1�-9cL���⻇m)�&�9�D���t�޲�ac�ဲ���H$��4
$wU�w��;]�����6ڹ��-�%�c�01�6Խ�9bҊ%l���>�4#��S:���� �!�;���-��$@Q��-)�g���DUgF_�C����,ߍ���q�FF��C��[Y�rݨ9½�d�ްn�g�M��ݧ~/;�K�i�m��~�%&_�_|�����1�>��V����o�|Gp��E�`�E�����wgkH\�/�`]mb���Ԥ((G�[n�淞�.B R��,�?�ܟ����'/1�_����(���D$����1�TEꉩ�V�m|�۝��"J���km��~�#EhwM�?�9�N��*a���(|�J]H����U����n�/G� ��O�S�Q*͊_�%�[Ъ��yp�[Z���ؖ?�jd<������_Uޤ�����/���E���R��\P	Vo�;�CK�| M�Re�Q��ϓ�b�Ds�����V#)��w|΍L�s�� ��ܑ҇���+�"��h�_�n+����~��J"O�����j�W�x�Bnc�YE -��]��En���١x0A~�S�{x����& � V�����Q�}�{5A=Iv�o��__�J1z�x�h�Gc.Ða�|yL�7��ɽLbMk4o�]���#O=n|���}�� �W����{���D��  ��s�� �\&�P
�-��v2�ˇS���>��ؿ���:��S��X�F/
e��3�9J������.���J�����4,>0?��g��$�o�5<�������*55Á�&��3<!i���ٷ�3���؇ :�"B3��L5�Y� ����9ۈ95)t.�c��_G�KA�9����R�́jU��;�lG-j[��*m�n�X� d�>:H��rv7P붋���h���,E��͂['��D����$l�t1���+>�L�u��qG���렺mc���
ҿ��� [���|(V"{�i$y"?O��P�-}�oMTW�� ��<�?'	L�#.��t֟�0ju�e�]�2�p���n�I�A&�;%>���Jw�<�N��\����糢7�3����Fܳl��B�΍T��c�w
Lշ��7�Y߀H$6L��1W/#>Mu���O��k^���B�͚�e��Y&�7W�i�-[#�y=�F��%gO��� ~FbY9��nH�U��o���q_p��H��/p�T��Q�\���A�P	H�a����?�&����ԩx�kֿ١�*����?��G:�6�P��~�.@@����E᳠��������8�t.͟2�g���y#��|9ŋ��7��Î�Q�Qޗ���8���d1��=
�J�
/ ��`<ʱ祾��������1k"��ɧ�;"�gWFk�Z�7~��_r����l}�m��.b�0��d��i��3x���'k�	�|}K�1�V�������uG�n	�<4�]AB����*�b@I�̩':ܽ+��KP�C<�~��x�W��_��Ā���?��|T��WY���Et�ʊE�W�ʙ}��r�������<����]�!�|�3����ğ�����
�
۩���b��5��!s��	q
���-�H��@�H<�l����{���2�>}�m�� f<~��|M�7m �8��;�����=���Q�� ������;c�����F�����*5b��,���M�q	!
�OԅgE��Wa�O�;��W�B��T]X��z~M�#t�.�O����返��">&�۟��k)��i	~�6����S[Z2~��DJʚ�_j��Y��Ym�P��T��J�c�}��B�<�~-.n�6n����n�g�?V�<��m��s�)'z��}��uV�Z�_ѧ��4�wr򷟨�:|xG��Q|O��6��y�'s�_��. ��� �
��۞1�~�5n��W���e�hyTI��&A�����8�q���Qֺ�XZs=j:��+����̹h���ː�ڠF+�n�ef��^�=2!~��b���v�g+��JUId����E���0��O~[��l�A��'�;����QM���&�v��^�2͚}���h�������?a���LRV|�L�"�B۹׳�~A;{E�0��g�x}ăy4����n�=��|P��G���4�Z�H�j�E���ã��?Lsm�Ӱ�o�β��!*�k)���LCİ�]s_���ۯNjX/�`qG(���Bv��Z�uOuQ�F��7��+�I/��.b�^[����z�?q�\��e����S�E�7�߸���MZ��s��&����BU�	TC���qጝ/� ���[�x�m��$��k��)%�D�B�=���v{px�N�� ���v�#F��"QaU|����r�q9�1�NHl�r=5�Ζ��=��8ЃV/�[���U�Ǥ�#��6�þ&<S�������^��/n ���_�=6�n�_eыo_��;\�j2pn�)/�T����r���p쐰8���;���Kl�An�/�]wtW?>���J� �Na�9�ɏj�ioQI�C�L��e��͹�s�q�c	^�~�RNY@�����!TT3�4T��� R=������Pb5?�����W��}A��zz��#k��t3�!Q�����x�E=߈��-�G���n�fr`��Ԕ7��(��Dĺ�mp

�oB�7�5@�Y7o7�ã֒����Wģ�\����|��Z��<���ֺԴ,[}X�$-4q�4T�}GW%(��ŁBaW�I����T���G�$����o���.YD$<������S^��_��V�����d!�v^�7F������.�yi1��{���������} lOᇀ�c�7Υ�L	�q\����FϪ�yB-�2��\���"�kቨe1xwM)�	��zYU#�F~���n%lG��N ��:��ˌ���Cd.i'�S1Z��V�c�
=X�dc����W𑻨k���7k�?���v�=*��1��#�-��j����n�J�/�^J�Rܡ��Z�+����wV<h��h�s��|�f20L���Z���N|�6s�$B���z7x��k0"�t�<\E<��yn�O��X��0�ٙ�D�� �0y;�#��U��V�ŹmD�,6����U�k��*���k��9�mH�y!Q7�P5G��Яu��\g��
s�V�դ~M�N���*䀓�7I��Q4�B�"�"ٲu���䚥qG6���:���m��&E��j��1]�if\�}���XD�J��r�@H�o�B�Eұ���U���Qi%5r��e�}h�כg�H�Ω����=X���E�9gH�=F�Ld�v�p�9�T�o��ҽ���5�iwGP�b{�^�5_ XR�;};�a��F��CZB��z|Z�_f��x��6���Rfn-��~�'�)۰��k(p�c�G�5��%�s).��mN�Dq�ٖ��L���~�:�$$���w�#�N�^��ǇM��k7���q<�O<�vB:��p�A�&���Kz���s���>C�����\ӗ��{���*�����o(�.��23�gY��Į(�ѹH}J���s����{��"���ǯbG��M���Rmغ<�BFV1/7��ٍ�bߏ�h����b�T�d�R]8� kA2��v��=�Eh�~���ƴ(+i=v�5;diൕG�D�C��#�y��N��=��;�[?��u�G�����e����{#�G�v�(�ohߢ�>X�,;D2\W�~���3�o��4J��ƒ�(zgb�Wvx%�u��s�@F�*�Le�"���ˈjcQ_�c@�WtXX��=k���lо�Ř>��]S�*{w�Yx�w��Q˧�9� �����b����VeQӴu��zM�(5���̶�y-�ٯ������ov����o��%��7������`8LY_/����뛑̙�.uu�S���WN���a{�6{'N�t]�M�\5�c21_�����A����Y^9sn^��6ӝ4�B�]�nd��"���\��cr�P���c�����%�v�c��-j�5�^��v'�/��i��:�Q�P.�q�zݼX7�Z?o]cy�׈h�B ����Y%���l���a�WK1�N�=`&J��S^�J�9����R�i'͗�1�%�BA�wu T.�{���w�/�ǌ:�c���Wa�Y�5��"[�!������Z(�9���2oF����  I�!�b�ڄ�w�{jҖ�Y�J�k4�;_��g���"�_�[���0}��t���$]䥜�gvx��!���BJB�lNp��b��]��3v`��_��@BWe�3*BFK;��u)�V"4G�`���%-�hu��N�y�3+�~_靨Ο"������,K_п��(kc�}B��K��?�PE%Y�� l���A�V_o���־[�,
�y�TIհ Ēݿ|���/����$�:y"{����Roz�E��� e�BmG�-׿<��w��妹��D��W�*��M�T����'"��Ԛ��/~_��p��������20A�>`l�U�{��͜=�錮o�y��G�U����ߘz�4Ɛ�ʼ��}�ѿ?
3��=�:6���ё�䲧��$�y~��(;�^S��Zs5�+V� ʕ���L�w��+��eG6�Y�5�E���A���� �F���>l嫐�ipL��N���Ӎ塍d��:ְ�ϝ
����ˎ�%rD��H,;U��M�j���j�C��!���j"d�<Ӗ���m� 3��A��z�WC�J2��ߨW�V�<���P隩���g��0����ٶM��n�G�u��sif����S��.����_Q��)_S�#V�4�8ar	��_�z���3�R�躑�fj)��E�Υ��Glr�m�n�ɥ;�rb��q�2s����F�`;:��ش�8�wQ�N��i󮔄LX�%�:��&vx�jS�Y%Z�?p�������� ƚmMVS��jK�e!�4�zW������
 �����P1�)%�3K]�"��,ጱi�ֿ^|����$��V?`��@v$� Q����klD��J����gl��O0x%[�l��m�ш|3�fU{c1�O�qy�)�|�X��=�OH�p?����$���%�b�.���&c��C#ꕙБ��(@��od��;�����,5+�fQ�q$5���[�Du	��Z�2��b��p�;�}�)�bj4?y ��Z�k����&�K�� { �Ë���JQ
c	)�0���9/(��(���̑�:��[��U�c�eyV.9��ꦇ�,[���[�i$����/�x�n)���W5�
I��3�����=��X�c��L%�,PF��C���-���*`�<��eq��R�MW�qv9����df,�8ǽ����ƶ�!�KF��qާ�,�������%I���y}���չ��1��L�$^H!s>"f��w7���%�(c��ٍs~v?0�&UCc�3��b��Ss(�f�>	<�n��>��0�rOV�C����{�O�yB	?���u1����x��{:)~��(ͨ�z~@;ݖhC�~4�`=$ý���ea�捎Ss�Dw�\b,�V��i����J��S�(0��ܖ#Y��uX�tz�j��`g�,�?����H���H
 ���)��-�*8�B-r�*��3��e�E�P5��E�P�j16�[]�p��b`@�>0�\jt�Ӝn</I5yȅi(>�§�ԈG�},�S���� U�#�w>�N����eg1g�lŨ�j�> z.��ԶȰ��k�+��a6K]\Ji����/n��s�����)��5]S�Ε�=���j��
��	���\�2� 3붞L�>\e���tul�Y��1\b�\W4�h��6[���;E:%�����{���Vh'g�=�6Mn9`��)XY�H���Q��E��D/`�M���s��ا�&��X(�rH���Ǿ�C�%�@�Ӹ��H��x�k/R����v,�`e`����~ "��T�1�L��N�����.���B��߯��/q�g0Lξw�kh�<���|"*F_/)	h(��6Di�iȣ��L�#��~(EI�M�Zv)>�g�KZ�]9����p�u��1<//�y1��R��k?5��M^�g(ދ׈
�c/TYj�t֖$�	��v�v�}=�����=��r�O�FYY@E9E*U���?(��&�ڮ{֓v�H�Û��z����]��eaX�($;�^e������{��	|�WЦ~J�L�B墯�{ƯÕ4���q���_��|ҋ�H��H����RG.Lj���"��@�{,�āC���]�S�0@�3�,dh��+�I5�Q������������� �d�蚺��E���ޒ�o�z[���;��Ϧ�&"���_�A������l�m���X�sf���w�T�������۾i<�˴��
�����Zw6t-��\�7E�����L9°����O,aTJ7M�}a��t7����Ŏ��3�NϢ�Z�]�j�:)�׭}~������R6�]֜��Fʝ�{Oy�rw�TI����ļ��ݶ���R���V�y�!�N�MS��=�>6k��ǄYe ���Z�'��5�N�g������y�_����	n���Xo'pJ�vO#�w�Eԋr�ٸN����C5�{������293^�� �oԁ^Y~� @h�7�k1�O�/�w�(�h��ǬQP~����]z�tp��=�-��Ƹ7`��԰n�瀞�����T
͟cu�F�)��*t��` <?��K�<:��r@��c�g�๺�y=	������{wF#�Z�xw�i�t`(�#�O����$dΦ�e�x��i�xm�PpzR���.l+s��g��O+�E�o��{C�hu�v���z�ޑ~"�f�#����U�V�ֲK�n`$uw���-�@�D���r��@-�0��Kl%t��;��N�U��ӆ��;����Io��!2��+��{e���\�`G!j����O� �M*�_��OB����{f���D�2"!e��E��� �7�����R�="fl������{V߂�ɲ�]� yU�S��Y��WhZ0����P^j��7�
��=;.��O0�����jT�;;��/��m+��T�^�o4�	T"�y�6�#j�=!4���4�M>rq-\.�%ӻ�����u�š�����p���J>U_��2�sw])�/0
'�'.�[�U[�1�k�U8�����N[��Clmw��S�	���AJα�ۉ�3�o�\�Pc*�i���-���ɟh'������^�[~ȴ�d��zO�B"|A��S���6�^�g$�M�vp�+ޚ�_,���8�La*T�0�= S�KU��7#�{ԑ7�sIN��`�q��ޜ�?��L�����G¼��wkɯ�Ki�6gF}����/�\7Z�9,�;�3I�������)kتARb&�d���������-�43�x�g�����~>��x�s�8�孰)��ο����lNd:5�V�^~�<�l�����|3Mrl��F��``�#ո�N�u�Vj�2�	�OX#���=ш��lC �`LP5!�W��8 �:RkF��3ч�Y�/��ci-�b��� d:�!���Ֆ��ce����0P������Dԉ�˙
ε��x9S�C<GU?!��u2�s`�Q�?*J�����(Z�5@1�����7d����n k�?�H�Ϣ *+96C���a���!�(�����zd��6��[��B��K���V�9�sG�9h�m��m�{������&�,�B7���k��Y�5��1�V=�Vz��c��_u�-�P���$ �Rg�I���8��#�-��?����B�/�Y�&�!d��J��!u�KR/-�e��oy���A��U+q8ZF�$�tI���D3-��Ԡ������-h���M�o[?������K�r���3��6�#����G�n[�/��bT�W����خ}����SH!������!��9[��|̲U�b�~��4k��W�ҠGD�Y���`C���|��k�7{C�ћ��������Ј�(�:��=��&V�Õ��Ƚ���߃:�4?q����%Kr8�f��4�(e9���Q=o;ʻ6gO�ϑ��Z��Yҵ����dY�<������K�Ak��fZ�g㙢A�ji�Th��kOF��~�).W���w�g;FޣL�H0�?֕�@�J���j�ϑ+����xǸ�MZ�(d��8�(�8��r��N7�+mĒ(��Ww���H$���w&��:l=�~qQ>��\7�<�~!�j+��B�D��%�@\d� a�i-�JSL#������؊ƔEM��"�ES�m\�8�y�N������_�CT~*vZ��g/@wv,UD���N۰b �7��J�󱉦�lR۹���{������X@�9��w�#c�1&�/�3 �X���w�ua�����r)ҵ�������8�1�XB#�gi��]:G����]*d>�����:��d�<��o�N�dU�f���]�Ds���Q������Y\6�h�a��܏x7UT��w�T[+���6�ݒ�������$H�a�ĉ	le!�w���:*l�������`�q֡���&�9ۄ�P�l���?���B�t��I�8xA��Ry)���-�4�|K`e�r��e����_8j,�B��zŀH�y�����2�0ڝ�ާT�E�H�A��`�+7�N�Xi�N&��˔�zL><u�C���JN*u~y��5���3f����.����2�����2Գ�9P�n�
�vU��b8_���(����=�2����0�+�ۧ�%�O��'�=lJ���o�1��H�:_�(��qӺ��t��8�j��,1�z�q�~}�����sd|b��[Y �D��A�o�L����	Hx�p�Ma���k�Cp�^ �b ��A��?�j�e*��i�z��yY�G���4��p1�-��CU��Ly^$=
�������W)�x�$o��,��w�6�,c�H��P������f�~��hD_���)PXE��������P8`��Y�R�0��Ju��������e!a|��߯��Y�%ފ��H��.�Qس�����VcА͜�r䉽�1��2}!�Td*}��.�CV,26Δ��_����"�����9g�q��z��Sa��?`{��8C��P��������QV)k�={�t�� �b�%����V�����a8������=��s�};i�������Qdr�lr����y`�Nc���d&�gd�
�?IOg���ߟ-w�n)r�ٵ��,K�²�MI�B���4rE��e.����;Wn>�A��ȨM�7_R�sk��[���c���X��wm�e������j�.�#Igl�G!��\�^c�WN�x�[�����P�o4�}H	��L�ԁd9�$*������*~����w��ZF��Y��A��I�E�zQ\`V��Hc�E�N��[N؊<|�ON,T���Y�rQ���$����M�9|���U��+�������tIvpkT��'��09��C�&A}bQ�ã��"?��N��������!�}��� h:�:�k��'7 �t�:���u�]�n��N�e�@�+h��W�Q��T��02��%%5��c[�2�Oj�؈z�(Y��Xl�2�Ym�<�-����Ìȸ5��ς��<=n���?G!\񌷿� �C^��rhPJ��.�j�ç��6X0ebE�X�R�ٺ}�A����i����+��{�m�
������r��U,�9ᣠ�Z���o�?]���X)�&+|��B-����6�(��zsc�y�[.���5f�9����Y�^��~�6�D��M��鴶J��mS�y2�ZԢ���=��o�kӬ,q�����a���g͒�qc��3�;Dl}�Ugp泶�L*��H*�R�ER�Lu��H��>��a�%!k���%#-��Q�(�u���a����G�JdDw{�դ2�M/Ǧ��*����G{`���;�5������oӭ�y��\�33���JС�dM?�+Udҁ3c�[5a��
z�8����:mK��Kȿ��@�������l�(�Q����"&RO����Ϯrg(��J�B��4�R��P]�̈���	�m�|��@w��5#���t�fqљ��IߡU��gjRٺ�F����5�5ǥ����9������;����J�_m�6Ow.�Ķ�mijS+�O%;0�����m��Ƹo�·[�Q�+����uL{�Vd�)[j�eA�ɹA�kc�\�v�g��
�2���N=AT�E�A�|zS���8xz����P)���������3(z(��c�)n�ºs��8\.W`������h��7�'x디���b�t���M(/��p.U�}-m��ZT�|��5���.TЬ ��(Ioysጅϋs���Gh:?~H�=��9����x�3��!n�3�o�����Ex�ضc�P�-��@�F�������(���C�fї��Ϡ�< 3�xa��7�u�0Of�8-�xP�ۀ�f����kHۦ.����cM��Ђ0�����������;c�D��*�i��6��9�ka��+)�g��;^#U��J}C$�r�nJ�����x9E�1ݵ�ƥ��d��9&DXgK[h�Z׭�T��03/��X����~��zYb8M�8!N��کHE�F��Sϋ�I(�U����y�a&#h��pUcBY9K���j ݙNm\Q�����?����l����;���E�� �pi��h�z�A��/��f����qpL~�\��x�y�n�LM%���'�\�~т��7�A4嚇�F�v�� |ՠ�k���̌�wHm�um%�""Uj���ӓ>�T��5Y��;MM
G���yq�G�����*b�{�|ګ�|�<#�
͟K=�fiOHb^�;~�Q�G��he�z-�^i��{�N����om�����2,A'�����k�����k�"�
5<�ź��lG��JV� �/����M�1�<����1������xڷ��0I��~�>#|�a���O�TMm��M�{�i-� �hׇ�*�,9l��C)�>��q3xy�@������J[��Y��>�������K�q)��
�?e�ky.s�QQ�6�Vo�iQ�OE5l���nt;ܴ��N�r��I������ƣa��`���ڻw�J8&�I坈��7���{�\F�"�Yʉ0C{�v�.�ׂ_�5�*�* L"�L���鴍E@�}Q�e������!�UL���H��G��2Y�L ��ż=Y���!�w�Ʌ������7l%3]�����\Y����_�K�y�A�PpK��%֐���79��AL_�|���gQ���KJ�F�
�uW\���k�=�R(�GGn��Z,�W4�s�n��6���A�g�a��	#f���i�]�� |�>p{{�W`pl@��XL��vE?п��d6eP�%1N��	�Y��G\��j졓��̱mL�Y�ZO��y���s=׃�+M����p�^o-�Kw#��l�䄳�_9��[ʸ�5J��!��/��Q��%4�r�B��/k����7�B��I�lߚ�ҷ��'լ��t���6����*&ݽ���.���@09�k�d��"8/mdy�p7���U���I!�rO�f�5�"��jX�"<�i���3���#��į>#,�H��AY,�n�����4f8��J�ع4C�{����~�z�� �TԬnVtw��Q�<�m�Q�K^�~ N��lz��疺���>�Y��������8d�k�	��?f��77Jҍ5A�a������C��G��9d3P��?�7�N˿��[j0�BiЬ��$/�f	��M�H�
)=>ن�>�g�r�ѽ4��!	m�$����~��~���X�Khr|��(Ks�
L����_~�HrV*��0��I�`����(>J;B>��7o�El]~^V4�q��Q��4���uЏ�΍]g�6�U�x�Wk+p|ܺ�t��7]@�5�`^rԈ���{�mj�������=Ϥ=������bs����H�
6t&���EUU�Ġ-�E1�} �s��8�G�P�H݋�l�h�^稬H���W'�´	Oy�ձo��!��%��z��<x͝~��JL!����5X*BxaI�X���&_�o�������G��%�6Kt��q�g�f�շ#��K�`�}g:0}�'�A��Ys��b�o���Z$�#�A���ֱ�*����L���ѫR�)�㹑�1��ދ�+�u-��_��liQ�1=�ɳ�C���MD/�A��Ԝ@d��K���Q1��r��4����'��f��������7��Ʊ���ݭ�A&�����e�<�NB@'f�i{PWZX�~��� m;e�>���u���9.	�%�3���!�9�%�d�I��*`�fj��v<6~�vFT:�&|wrTpb%���JY��m���$63dU�����$q��k��#��q(�S,�k��}qbCݾ����t����5��b�}XՑ�BY]�,T,r�O�J��Q�~Hx%��KҶ2��UryTx��#Z\8�8:X�bd���>*��%n�x����E��gk��S�����RDX\W�g�R�(�NG��n-��y�t�&�G,A\!f�5��'�T�3b��<Ӽt��CE���{����kb��4+�ٍg��s�)�{Խ�2��	��������,) V �Ԁ�8
��䏃2<�1
Ι!���Ȇ�'�ۅ*��T*Z��|��b�KJ���M�#]sdq�91�#�:��v=��T��S���ǭ�]R����7�F
�����ȹ�ø�X���v5�F����<�������ˡ��?�]We���2�Z��c��WЍJү2��x��t�o�KĐG�,3g��;k =��C���
$��x�rY�A�L��}OG�.Z���;��.K�A�H�	=��uu���EPL9.p�d���-�}�št'h��fuMn��V:��CV�C��p��$�i��>QY�dj�G�s)<_���Svn���7��k�W3(ԙ$u�y�L�aa��at��m���L/";(���|�kxD��Q-%`�~I��������x�L�����Jǳ�U�����[�SZ�������@�%�F�m�б���\��v<��Z����hSZ遞��.j� ]��]R͸� Y�X`J�`����F�}ĳ�=�_i�v���[=F��.~M\���ϲ���}�ӗ���U_����g��1��U'��3�	e�J��j"�(��fӱE� �n"�ज़�!��r���@]����)>��㏰���~���`۩�Pv��%�X�i���$�@�� �<����[�!k���O.��%��ڑ~
utl+����Y��P�si�-�`һe�dz���U&�ǿ���C}��~�5�-�ѱ}p���_��^y�ё��5�}5��9yC��	�G��� �~ɘH]��t��]���T�U�8I�7v�4#Ҿf<x&`|�}E��Û(�뚇ѦPb!�hJ�1�'^���v�2�ڤ��w��25�8�/��V� �n>�����Τ�A�����X�I�1b�Ն�D<�����f"Q�s����Oq5�P��, �{�{p:¸(�aOM�r �ǈkN`)
���xV�������0<�[�ٙ��\����WlBQ��"��d����Xb4�r�2�����ƕ�ڞ����[�,��#޹{ѵ{q�WC��y�b��?�tȤm`�#�2��'n�m�b?L�K��U��},���R_�J�bu�~'��@�������ⳇ���|�G�#��%S폣�����w�6���Bt�U���H5p���*�߼)�<��U⥯c(�7�!.0<P�M��r�*�JB;yW���o��-F�VM��gh5훴|�ɀ(+�����U�i3bx��K�A�17s�(i���d���b�KO��r�-^�#��b����3��� U�Ҭ��z<?1�  ����ơ�-��Aɳ0�����e�ө�4h��sq�����q�jҊ�O����B�iG�B+���C��/?~[�[|�bi��k=Ra���(o �Z��_����ZR�+*p��I��!�}������y^�jRH=X\�:�3	����
P�v�G��	�˒� ����ls�(ˇ���4��j����:�n���	6��U�UJҸ��H	9�3��>��|M�s�a��IZ�����WͰ,�+;�,D�����x�-כs`�� ={��+.޵�GO�П�:��<z9��S�,��d������|�\ 9BUQ��ħ�6��m�Ӝ�}0;�4��L�ŃF7NM���� -�
 ���W)^�Z*�w�� .�g^Wo9D�F8_�{bl?�:�R��-Tu�f
.�&PH�Kg}��:"M�!�{�2���2�Eh��3��6d([���q�4�vɥ �=����=�٥��.�?�ʆE��e���O��b�|ۜ�lSD�:�,e�K��Gè�_[oC=���J�J���>2$��׉X��;1e�$��#�5�$����mǡ�FL=�["c�Q��:���^d�`���8������tVA�c�=��e8[s.N�̣�y���b��� e
j
L�X|�E�O����;]���u�B{�K'�<�.���<!�{#�͑��:��SS�!��C=?�_+�6�d^�6����z<��z��ɿ�޿�Σ,� �+�ӕP��%���@�~�N��Y!!���[ڬ5/?�mĹ�v_f2������݁�Lﰝ���I��&�5������Brz!>�#n$ic>e��k�|��%��R�T2/������
ß����W��~P�� ��UU{�
�.z)�JG�*5ݾ����X}(��J���P�����D��"1��l(-�G�q����E��~px� ޙ���<F��>HC��z��L Žc���rBH��|qrώ+.�IE���������w��s���:�O[�U�N5Fͧ�Ugفϻ�۩��!��)����3��㴇���t�1�kz�����09*zf<j]��t�82&��yh��Ů-M��1E�yy����s��\Zw�u��?��ۼ� �u�0�(��` s�d�56]�d�����P\m��w��\Ɨ�J�ƴA��Wg7��j*��-����I�{n���p���G)F&��@�D�.����P�~f#SK��:c�HeJn�7��y��ty�y	�\���J��Ш��sQ ������ �	^�yn���wc�0%w2մ�j��Usa[�@KJJp� e�w��ib����f9912x��yA���k4��|K��D��nZV���I�=���Yjn�"O\�?5�@x���DI���kM�5���YͼI�B�ՖF�h&��H�*�6�F�ZqY�޾Ui�>�R����.�-�Iz��.~S[�x��+�yr-�������!��u|x&M�g��a�~ܴC�
��%��l��#J�02i��/� /�ٿ��o���ѷ���.��^�ds��ǔTN�+O�L��F�����ei��mˑ�D������|�u&(D�.��u�{c)<���Bq`4�Л�޷�(%ǁ���N�z>[)L4�/,��rg��Rv�>R! ���n��`��L~�<�U���Fm���:�DJZ5y֔+�t����c��-yև�ԸTv�f�4Y����ik���P�؋ek�7�<��U��%��آ5�,.���|䊼���z��D��v���A�?4M�M#�X�w ~�����y�q7(������l3 �nW���5b׸���\P�?�L�]����լ������w�h����4N��`,�T�ᒯ�L(�ۗ�P�V�X�p�8���|�u&�K��0�g��X&`c��}#�Yd�ժ�zá���+2 �+��h�L\X8[i+�֛���`q�o�D�8���67�_���0���p�=>>�)��C�&g6,�x���������(5�����=���zSR 4hl&F��|���Z:���xlV�#U����!�1�J��.MdJ�oꅳP�K ��q�TI�.ك���+����}frV��
����p��O��#���_%>��Rv+Rx��LG�g/@~�nK��I������Ax�
�&���1�������W��`����G�I4	ʤ@v����hGyz '�MJ��)ґJv(��H7Âc#������c77�sXSy���4S��Y� i�{Q���]���9>�x��� 5�6��ŠC���rS�<��o)�k��S������ѥ[��x̿���e�۹D�%u��C]9ݫ�����P��9�:����=X��G��)���hŢwr<gH	��}h��Ӝa�����7��Mϡ����s�׀��׀<l�!��ЗF�#��d�>jѠ���$}ŕ��j�I�يڝ�j+�"���Y�m�08�k�ݎ�r�?�ro�}m2�5�6�q`�5����?�������L�T�M��J@%MDv̸�+MT�~��3:�ؖ5�J���;K�a�\|_! cW܌+�ގ�W^P����f�p�;.���	^]�����^�
g`��0�}��{]���_^x9�{����~�`�o�UÞI?P%�>���	����(G���#���X� �Md�"����	�����E k��V��Ez-���ܫܯ��<Ǆ�o�gwm��e���N�V��g\+�'��^�8AH �^|@=M<IO;��Wl�Bg�M_�F}3!N�w[E�y=trͱ�h��(<�`B2�����������MS�V��;�Đ������+a-�p������
W��ůL����2��=��C�)�ROT�U�%Nz�r���nEM�l�<�M3���KЉ?ʍ\��P���4�k��s.�"bԵAH�av�?Y�!p�q��@������0
����Xfmb5Pvg��?yHƼ����ܽ�=KF?z�$o�5�Ӕχr~�1y�JrO�<%O+�d�=f0�8;���2҂6��Q�~�����j�xվ�E�h��nfA;���P�w���R����A��z&�S���Ä�~�[FT%�KO|}8��۽���n	�ޤ�޵���������G�
m���NT�mmǣqa����������(���CB?C���Kfq���_݋r���sx�mR�$�Gk��59�0��t��-��S�������y�x����,c��x\%���}�M;�%z���u�����f�1��j��B��݂�9�Æ9���8��7�V;/��c�N]�U4�h��41)�"jn�?�F �is<<�Ap3~,6��������a;�<�ND�y0���i�����ǝ��k�E<�s���p�d�\^�<t�Q��Ծq��kԕC#C)����m��я�L�F��n�����O���v3������=�ݨ��v�8�1}��υ.f�����W�NY� ?��йƏsޜ�i�r�F���� _�� �cA.�=�d�qå�M�+�9��$���I%g$²O������3�יp��o�P��O��?s2�I�n<;�-��7C�^��P�Ớl�!܇�֦� �r����>�b�Y���^	6����؎nn����W�<�<�˱���	N�/��)��\��L^'�&^BA���lAGÝ��CE������Yr�A�-�L,Q���FR��703��Gۍ�!�OG�dB����Ե�>y8�:���g��T�dC�L���c<���b9s2I��5oyٌ1�� ���)[�T�_��bɺGbw�A�pu�8L�O�4XU/��&�!#Y�X��sZ���G;=�%�����K��Ŝp��r��E���#H����2�5����-Ƕ���$<�sat��V�n�?a��J�k�-�g} ^���i�+6B��>�b��/�`'���_˧{���{�h��=��^ذ��/)�=VQq.������>�s��W�Rޭ��5�AQ��a�d����_h>.#y)�#"���t�咯9\0�|!���/5'�!�pa�����5Dgbp��$��ɿ��*�gK{ 0�B����nw��-��"ޢ?�b%�Ah2T�����$n���H�Ǌ�3m���n�����ޥ���w�Dd֣��\}���O���*t'� ?E�"�z�A����ߡM�I��K������gl�'��� �.X�A��r\?����%��Abi�~G֟А%�jK�|G,���%����N/���0QG�9ڣ4�t`b���z'�|K��Jm29�(��.�l�I��ӒZ�#��t�uǭZa�vr�y��۠���Thk�0�� e��Bӆk&��$,gj��d4r�߬�h�Qz����\��-�88gB���n1v�b���B�����8��ٯ?	K��鵠�4��V�'�@Ŧ������=)ҁ���M��\��4.�"�XRl���C`*���Sڅ�1��F��{�U��1FH��I)m��]t�)��c�'=Te���[���&]*�\��2$������&Ǽ�Q��[�Nr@\QbWT}��C�s��I�N�J�!��Yx��������<Y�,z�b^�d���Boߨ�?g�/�O�j=���
�P�S��F��7�MSy3	.���6�I������6��B���U��փ�e�髅>�E�� `���7�`���Il���a���?o@�G�L)���~5dF�q۞Ek3�E$���Z�����F�wS���xxL��Aè<���B�F�x_a0��v����p�yjP��8w �$�۶좴�tW,����Nl�d�l������p�}[��=��m#���a�!W�Ĳ�چ��uN��� ��}�'��e�|:��=Ћ�����;v+9c�g�V�BCS��/�U�`�/��Y{���F��P��Bڂ-��R+��l�^,m�[��&����Ta(pJ�~��2�������
�B���$��{��~hBjCc�Kw�q��$ъ�n��Ze#D�S�[��펦�Z�^k��z#N C�C����&���˔��#j�Xkm�d)|m�y�>
ݽ��P�P�]�0^l�q���]1�?$!%h��8$�#�N�O{J��ף��!��*�;�zM{Ea{��q`�Y3�ɱ�jUU߿�2y^&n��~�� �ȁ�e��h���#��@l�l�Ih_���jmXe��Kp���1���޴��5&�_�Ցw9J��b&R�A�r(�בh�vǻ� t����'O�6���5�z��mxq�%SȂ����H�5��z6�4GZ-;�o�������=<��2	[i���0�)����<�������#�A�u>m�^��u{r*�͚��x�<t?�|4��k ���N�/o��H����L��rY=�~(����G�=wTz����8{�3�e���]�s���5�<��d���f ���dj�O1'�H��#�ڕr�	6]o���Q�95ׂ\���G\4���]3�*������ϳ����gy����!L=����Mh�!�4�4Q�j��s�Ai�>{zR.���T��P�Y^䂦�o���?Wl%{u!
£k�H3Z�*�r�ar1���Yp�g�S`�H<g��$_E�Nt�a�<H/�H1��#Xl�8���\�uT[��?#��58�R��)�wkqww�H)RB���;��C�`��_����g=g�������̼df�$�-���������+q��da��=&�cq��]ꭳ�J�f$�!��>�0t�i�an��צ�eǹ����M���a�mw�{H�KQ�Ɩ�9�" B�g���u���y�[��Z}�N�ͧ�F|*�O3�ܶG1 �W��1]>�xƕ����WV$P��*��-}bJa��q��Y�ap��жy�&��G�Y���}1�z^w��'�Jt�����|����"�f�D�l�W���؀:��Q�WÓ�NW�
�֧ۀ!��G�x�;��UD_)?&�21�+���h]zD?.,G�Z�=�}����p/���P��mOK���b b�q2�_�����7�m�7h���9v?jݭ�0b�@�1@��݊�\��݉|�d�1�aF,27��T�֠��c�'W!mcY�A�fK�-���n{}ޅc��t�*{x��Go�铽��q*~����)�
���o>�p ��=}�oO|�"<�ڤ�nE���;�z�k��"��l�����u;������ ?�����1W��Ѝ,���Z��.�P�q�-B���D[���X��Zс�EW�yMB:��+�'�2�A�_�^�������>04��7�[Sا�D}wN����li��ȾV*��ֆ*1���������k�D$q�� ��AW�י�Ư��E�=��������L*ū�G5��#.��*ڹ��v D囎UC�����" ���ain���5x����8�"�{���N˭��4q_�L��̃�0'A���d)�����������Sv��˩��E�缾>�FG}�=�c5���߽�>y�ڐ�������
�o�]giC_��vO��/��
�|���0�ޮ��߾~�$�����p��e���Rqj��y��SHKPwe�r4�S�0o�ɿ'(��<�0Uuaww���=z�o^�����w2P�Ū�q|ܬ�գ�`����k_��nߠ�X�'�A:g���*Y�1�D��G�/_�g�#sMiV�����!츀�C�W�9Oa�����yHV�7}>�更��������Q)U��n�Ύ�b:b�\?�Ǎ��&�K��¹	d�FMh]/ʍ�qF}z$1���(��č���V�۵��-&u�R+b�l�C���X�Ya�uf�Q�c~��G�&�i�YV���p�� 00+5U6sH�[�&�Q�.���=F�_���!���ރG5)t1�/��G�t�н�������P5�y��<P$�V}B����f#��;�+�d]f'e�,f��a:=�L�����wSxJ�H0_���-�0�zi<l��n�7,��>�\�ͳ�C��e۳��,d{�>�B�h�X������+�9�3�v�w,��Ƈ�d����]_�S�Xz�m��*����n�^���*��_&d]��|�>�Sn�/TЉ��`#�o�����p����{�����qdz���!��b|���E�<��+BM�#U�L8QCC+qyu	���g���+7EQO�Dg��l��A�g����!��A���*L��t�P5dnaE�HY�x|U�����>'��Oh 	�r�n���+��7��G���@�:m^QPF�v�J�3nA��%RC��փ���h�)��ҽ�l���j��Ѽ��(�M4�_�Jڔ7`h?��T�m��z�@!�Zbն1x�F���l"���^k4�l=��	|``9=�b�����������M�dȏЋf����"�ơ��W8��f;�E����߁>�vĳ�=
��l��'O�ހZ{�������m�!���>&&�����aG��ה.iih,�jB3��KJ�W�5I��ip��$n6Cc�s,;w�bwZ���Ă$�(z�3,=��s�ܷ�+��5�~[�:h��\0��9m��ݪ5������?��7&i^8���g��ʎMˡ\�u[�@&��y���N	C2KX�Kj�TS����o�'X�O|��΀����4<D��!����)A��L���S����Kz� ��{�N�K���A�<6�?S��iJ��o���YZ� ��>���c�����>V��&�v����\���ɜ!���\;����C�,cr��������FL�ਜ਼sO(c�Z$�Ez����S�ז������k2��}�y~���^(6��˿�<�R��_��;H�8��4.5�)V������i���1�p�K���O|�^����_/��MFx��^���h�SnR��qY���/,5�*Ƭ��vwԓMV�Ah���޼BLF�� M5�J���L�oW��g�X7������ل�� �yYO�1��B.�썕guHn�s��έ�u��^Ȏ�_�g�7��6����T.�QN`��~��V,��1;��>__c�����W���CW�r"0<�<0�-���\n����D-P����)����U�����QFEz��R�1�$�GJFQW�(�M���E�6�ע[�1�G��j���-��&��ʳ���z,;]��v�y8�f.�cX�w�λ�;K����2�5�y{���5Y������7�/[?����gjT/��&�Ķo�}�E����a����r hRF���c���7��/+�q�����
P��GoZ�t?Z�W�{+��X/��W,�eX-5=���,n�����|3�U�d-K2���K����٭�V����������5Ѻ����Y.�~goOJ��.5��[�JL�R4��{�ҡuQ��]$��%�3lRL�OM,Zsy�ʓ,�9�-���y�_�$PE�Ф���M�,�E�C�7��F����H�I�&��"'�7�߶�������J�H0�%/~�Ý#Sf�n���o���?��7�{i�^��'���wxR��&�}��a�ap�!��B�zYYV��-�Ƣ�݋��<�3���N��0��N�Ӿ���0��kƝ5��b?��F�)ն��g@]��g^���bM��p.JJ'ǅ���1����/����K5��v�q?�k���ꨐڶ���?>Os�|���9��I�Snh��Q;s�}X��%{~`��p(�y�ɇ�g�K�d�X��zӹ~/��ԟ�����|#�͑��U�k[�B>��D�f#� :r��!��r��%��|K�]k&�p�+N�R v���o� ���YAzPQ�l ������_�g¬c��RN4a�c�>f.~�<&z�x���K/肚�3ݥ����8;;�^V��<F��,�4ιcG���c��/�V�	7Rz�:��2��W�ӂ����=.ї��EF������z!X��u'��j�'��3ž��B� 0�i�� �;�9�Ю+9�U����[�g���i;�I�Ε�Ra[�$��_���p~wx�I�2!��PS�Vq��@��B�f_�JwW�)��WfX!��4=��T�8���_���N��OjX_��W,��0Ѥ�g�~�����11�����d�$3���Q��N�Pe&gZt��٤�F:]Ϙ4��) �|��m��Xo��b�xS��&oy����~�{����D���AS���x8|$�7�L�܆�R��2ێ��@d)�Ca��/	�<����Sm��N#��s�W�2!�{޿������z���<�F���q�����f]�="�fERA��O�[,����F]��V�zo�r�٠/�3�a���マ|��s޳|N��8����i��-��������v̎�J�k��O�������c}��Dvc�/Hav���ܹ��oY���\ͤ�=�������ә�}�y���9�F�Ak6r�'9��$�!��˛�2/8��$�z��)�G��6n���M�um �'Vg�����^�P����Є&����oܭ� jX��蜦�c�n!f�S��B��dpX�ܶ-��ǟ�5�������,:ED޳*�?�Y��x��j�i7,"#3���#�%���a5���l����AW�4�mTL�V�%*X�7G�����F�~��_ �ܷS��"�����X�:-hXH�%���.u���d:g}��Mpf�Lʶ��~����h�������〥�e_��J?p�m�&M(�S��F����� R��yi7j4�b�T�;��I�(֎ɱzC���S�� 
�@)�lȎ����{H�1j7���ݯ��}��������4��R��b Xł&�F�l�u��{�"�����x���|}��1���pi�p��)�"�<���ˉ�Hc	kǳ5�QON9��]i���K�G�����E%�J���6��;��nr,� ̊V���q)`?Mh�rxR\�В�7���l�kU���90����#@�~��eD6�yH
6
ss��U�W����Q�f�i��"UW�71T�?��b���5�s�T�FP���q7,V����vpͺ�E�'g9�FF@O7R���M�����ͱ��o��D��QE\5̽ܵ6Dd44�Yv:����Sȗ�o`����0�?&�	,�/e�老f'�)�Z��Co�Ak:k)�D�wOJf�S\)�+�:��~�'ګ�Yql]{Q�;d�d�hc�w�#�4�ωt�<�!�#8*�H���:�Ȩ�G���*���WY[�X��v����jA��Hɹ]���].��n�_d7���i�;�X��3�;����o����Y��mTO������Ro�����|P�XB�K�l���]�d=ӎ� ��/��!��_��Y��!~�-���c���:)��\����Xl�����y'�X`��'����o�=ǆ�ҩQ�m n>f��s"h�}FG�>@s@��Z�ED�W��%��%��~,4n�|�4󳑞E�tWY�_eB������#�Ri�Gg&:�`���� >+u�te}&����[ql�X?�t�m-���9���~)G��n=K���@�F��6\�|G9���_�7���=>�JΏ�w�G�ѱ0`	J���8<?�� �������+�iUr���,�3c��
/�sW�n+�ܗx��ߞ܎�%�e�
XI�d��{݀�A�ϣ�j��� l?�I^��f!����,�d���|��d�e�G�<�VFaC�:~pT�L�L?��-��6�Eh~�2����a�o������J��?'�D�����Xy��Ih<�����B0	��<ڕ��h�"�,L�@��P���/+��s����Ud���N/�u��M�ض+Ke8K��uŰ���)?"�$��,���>����6��ḅYj
�K�6(-��\�6���|��[L	SQ��+2|������Y,ٯf$�A��?����y.����(�N�wdpB�zɐ���ZY���+u��9����Ѩ�����.=�!gy	�}��MP��&���'��g[_�n%�ұlp<)�f���`���n���.�>;-�P R�g�db,=�)f�aq��n�#����<8��gt��rZ�����zV\צ�����c*���B�>5���_���bF �S�1⍇=���������Ck��0}u=`�y�"��s��zldk��XU�����(�~	��@/�ry)ߛC�[ds�s��"��ވ��%�������EKmnB��]��7��R,E+$n+|fB100����Z��5x���³���tP]@]��*u���>Y�X9JR�B���i���p�����&O"��g�$qw�1AcL�_�ܓ�ZƖ��ǯ�hi��Y�Oou ��օ�>�ۤ�j1�nTDi3���'?ͻ���>Q����;�aϋ�+�118�L�MySQ�B���kF�d)�V���֛E&_�<.��_��W0����$G�Q�i�=�8�t�C�X�0�cV�'ap<X�Y�;�,�B�������:�������E�0;Q{FwX]����"p6`���=�1�%޳��ֳI2=.w�����곖%ơ��vFx��{��J�����:��c�G�[(�)L[�I�7A��-�/J�32��|����K�|�c�hL1��^]	m��C�5�u�!�3Iyq�n3�LF%#�8"1Y��z�]V�/����hр���ݛ�sscY��ɝ���4
��V�#�J�����C���x�o��p'�p�jU^�����P��%�H�٣j�/Pg�G�O�m6D�U�5JCkzpv�0>���� i#\fc6���=�n��~��f1��������b��6�efp�m�O�縠Q���&�&Tň��v+��bZ�+�n�	���k���	���_���p���{��}M��A{N�
k�?k��.�D�F�]J,S[���2a�^��+��֘��h����+O���os�{�6og�I�l� lVI�hu#
Շ���_|}>������}��7��;�Jo�'�P��9��x����dO�ІY@q�JX�^d�f���# �.�QNG���p��b�՞SkGv-�ӑ�Ekg8��VN��f������0���������R��1�G֕�u2�6��z��˜Ht~�h^צ���~Yp�zN7sN�;5�hh���Z|�.!����� �L�S�x��l�ܼ��A1D�y�y#d�	r�y6���%���X�tlqO5�J�a�~��e�vz���.(cZЧvP���̚�l��m���� �Ֆ\ �0��(Q\8_���oeaIY�D,ʋ�D��sܪcr*Ҫ��}�%��Nl@{���.�5C<�!��hʴp��@�V�GA�[�*���(��c�?u=�*�)i�!�S��8N����,� ҭ�G��4�B��bj)��F��3Rr�T,q����E�F��䦳?{��u¾x�����k��tS/Ǝn�D7��c�Sit\����tϧTK>�����b&٨�i	�N�[�k1
��SdBC>��.-����9��8Ñ�O��p�8TQC������ 5�T{UVYz�:�J��q|��MmR�|�#8�ыExns���27G ��qX	�]{����� �l��~YÍX�E?��ک�sx�9�=��/q�Zp[��+t�;KF�`�Rz���}+�	)�4��F(	�TrQ7��v�ݓ�'m+8����y4T�CH���8���氄��vq:�2��,$q�J
��7I󂏆6����.�ь�?��5�Z��=��]q2��݄���	�O'f�~������.'�'��I`�&�a)+�^�\��|Y�±���Y�aǶ⬥3��?H:�IV�r�U$v��Ĝp��M����ɶ���B�r� �q���,�;,�H� b����;�>b>�fJ{E��5O���&� �	Dְ��厊��s^S���&YPr��Z�j��'}5�"ċ�0c�{����t�*iZ 44���vl���bwvL�`�	���H���l��<����ck����.����ę����a"j���(�2<����:	���Lᯁ��!A��/�����&��zO*;#(��Ҿ����So.I�|��g�cp侹J�>/��*s�N-G/Y���~)���ϻ}� �>l�N�8��i;��l���Zt���Y0�{Lfh	G�`C�����"2��e�WiIKW��cHsH�ҾNHJ�*�D�:���H2�"A��
����4�#�H}9� F$�����)���5u�^�R��X�R��2���hN�?�(Bu�����ǵm�Q�|c�e,�[	i|�����ٱ��&\z�F3Ae7zL�oe<
S� �}R��?�1�}�:�
 ��MG���\_�s��D�#�KL�okx��ajĮ����e�2A�w� A�t����d�F�6ʪ�Q	����3�z�O���w��d뎉v�������P4T�y����W����-o��0'In��s�s�pE�H���C�����k)t���*����#�{��DQ����t�I�?��d��vw^Pi��O��~�ҡ����T�o[�KW2:<��A��:G��1�i[�ߟ�������a؋��AV��0�F�K͋��8�ǡޞ\�`c)?q�L&�`Yy��i�ws%�\�#1CD��s�զ?��Ӛ�}1��<�pX��UIt���v�g���y+%�S������:a��6��-A+�}\� ��:���%�H�0)�?���f��`�����]�50+9hCY�m����edh32�4�������	�I���v��E���C8g&�S�f�c�ջ���.��v�`�`ջ�,���\��ñ!Kհ��byu�AڭDN��!��d����*�NOk8�a�}^S�{#n��w{:3;�}�ti�a:�X�7G���ߥ����l�&k��g��+�[�į���΋J�E�.X.���w(����Vej�(�v��tf��y�,ZQ���K��R�ד�;�A1#�g��Y���X�9�Pb�d�Ŀ���%`���EͦBnӂ����WE��8����(����8@A����q��ݞ��zqj/!��]�zS�Z:�&`��\��8zp�vV�@�����f��wc�Rv+0ϼ�?4�}]���gzr�^���8��R\��h�����?��g&�fThQ�7�.�>	.�\da�c�8L}�"�YQd\�~d'�ۤG(s��?�t��A����Wn���O��݁}���fп��\��T�y	�K\�3W��L��K}����9�C���p.���܁*����?yP�}G�����C��M���/֫-
z��������k�0w�N/�H���0*�k�O�����%�oJ�S�<24s�œ�&t�)x�C�O���L2���gQÔlv�Ԝ���[�dj��x��:�n�Cctl�Cq���+�����}E�'�q7����:��;������S��K�J�)�Ч/�GH=��d}L� !�%�I��w&(�!D��Iqݔ�nI���"+n����������c�Zf݉(w��V5=#"���?>��,��	��<2yu����G?oj��n�R�E�p'�	�1(ɑ5��Q��'{ߤ6�T�S����		z��5�*yz`}>��z��jVv�f���a���肑�Ԋ[���_*�N;�(�J�r��?Ъ��ސ�:e��np	#�����Em�룸_�8��� qï�L�����w��v/���ē�2�ډ>�����j����\�.1���J,��?`y��ֲId<�{�	S�Ìl�5U|��`,���F1�����A�j���Y�P9 ����v�U�!VJ�i7�-Ir���8�f�B�O5['M�[��ĺ ��@U���X?�m��&&ZN�B8��F ����+_���e^Q���Ʒ;� >NJ6m7���8rP'�RLVuY�V��#z�=wG��^�����C���8O�ZxNUu��}ZԇI�0T+��ܹb��/6�h�4R����4�#f*�Ո��%hC̱R��s�.�kj�_�b���x|�@RM���)�����$����fP�K�ĚS��s=Z?�[���J���'-��[q��q�1?��i�j�|��t��6F	���ic����돫�<��N�B�r��/�&י����^G��<�R_(a�&RǷ��خ7{ȣ���{�}��}.?s�ƅ���vR�H}��L�$5�t�*�����!_yӽk�����f#hTv�Bl�,,�:�n�3�bU�GE/ǅ�]X\���ӗ�2��#��o���ݗi8$�l����b�z�A��8���,X��0�����b�k��z�<u�I��]�?�+O��k�FHjѹ��9~��o`�\�V�x��A7�;A'�VcjRw��Ku#���i�3�*tEY�'���o���7��
1=Ǭ�$��Ɯ5��M10d�܏Ż�|g�Ot��j����������c(|w���s �h��L_ %��b��Xݸ�7��g�f�;�^�~�t�?��u�n����ʘ1��=W5y�xl�>�/��0�+�y��U���gAa+<�
��al��ؕЉ���� ��:P��+�ħzs��{��_��������v��}k�[�A�3��2�((Ց���6�����Yn�sB:2������wzo��
��%yVw��\���$O�/��.w<��O.�]��I^��mL�&�}�m�`ڳ�QE�<.8z�M���OH*�ߊ�&�Y��D���=�Qd����O��d�:�>�W��
{�ZF��{Ē� 
V#�w�
Dߴ�	���D��Y��UT�
����0)"BN���V�聑�^|����d��O�B��k��U�WpH�<Aӆʝ����2�V
\r0r�/�udʐmT�tG��T�[k
��F�%ªnc�m=��3ǹ���*��Ց�vEl�{�#K��B�n��J�K�UVR�����F����sW�1���/X vzT������a�it�-r�Hy���R�tS	?N��d�'��ټR�g��m�z>Ũ��~��ӀlB�\��S�a ��fp��|h�)>LJ3['³����k;���X6'߈��)�q~o���
����/���
�k&�-�n6�[��y��,�VW���ҮF6��g��B�A@E�⏗hք�En1���f������ Pww��e�f=���jsݍ�췇JL���J���=΍e����ю��X�	Wy�q|�.�����]�{񪮺ݶ�
�
S8./�0�Zw�g6���x��&v����m�1���Y_�6��j">n��p*W�H SA"���^M(H�=>�[��:�"h�1�!�Y�>}믤lA\���W�Bn�L�H�nhlWSL<���<-�޻_��}���y�����!�[�?蔐�c�i���qa2h�~��ϯ_� �g}�+O��J�b�Cզ�K��'633Nd|s`���&�
��$S�E����V�Ƶ�U��t�(���n��4y6􌘳���[�nt���r�p�2A̖	�-��so<�Q�e�g��w5�����2������Ck�%��*D<�[�:��Z��v��=����F,u{���N�f,  �� ��9g�ءG��<ß��^���yo�G���� Ɓ�
��P�mw�MO�eN�CaKǠ�9���p;��	�0�H2s�������ܺ-*�A���>��߄�R )REz��bX�T��׆��2"5���*��N��EA�Q��$;��t�<�T��d�x�M�n��f��)�s�Nd���6���/k��c��j��I1����z�W���!ŏF����.�Z{ԇ�����!�v��9ie������}:��..NL�:;T69�t|�ۼjgeh�xaB�ӄ�Ζ>U��;�s���'@��;�����Ve���ꇘ�rN����#�HF9�kB�̬֡<h5�A��D@R����/���Q�l�`�⁢�4n��bt�#3�%t�&h��B��s�2y�ܐBL��U��U��[���2�陿;��
��b#�PYsL�[�^�iË�����P��v4@:��9	?9��T��9(,���f�AN�oPB�j~��z+a������o��9��M���Ge�̛�|��<D�h��"K�����I�A��� �gKH�4�ړ�N���/e��0�F��4��m��47��Z�"�@ ��.M���@���{NlVN�r���9��Z�O�W\<3ȢCe/e��B�}K�?8�ƌ�[�
��o-O)m~8ǁxc$8���67+���U���v�YLr�R���Y��J��s��ab�����r�@�&�)"}4�)�Y
�#U��tg��d���h���5�g?�_Yܧ�#�l�i�h��3X��0�6��'�mR9�z��;�XH�s<ks.0XNf,t�	�H�흃���R{��R���g���:�������w~�_c�^��bI{'u���g�~?8~�Jv��6��)ԡP�����)�W��X*I3���i�oA�5�/�����x�6cýI{_Lg������.ş��y���Gw[~E����#2x�yn���s�D[�/>�%�k�i="�E����E�m\�����%i;�r�Z#� �،�X�S�J~&ǳ7{Fp�Z:1�k1Y�d��-`ݿ�nV��� �!��ʼ61Z!z�9�(|����Ī���O*�H-$��HIɓ�������4���8"Wg�i��j-5�k�����c�<H��P^���z[6w��x9��\�5�m�sJ��"�R��m�yS����N�kJ �FI)+w}��������=Ep��FP��Foe'|�l��.嬳X~T��c[����e����XܣV���IUN��؝�H81F�e�؛�g�a+����k�[ǫ+���h���CCs��%���p��_%�Ѩ�����Ĕ�щ4.h�s'��a�,�����Ceq`���k���nC)��D�&B�n'o������pa{c�nw�����M��5
��͔�07��c��*d'�����ϳ̢��<���a�@՝\�C���Í2G+BQ4V�ߎ�?�?WQ�a�O��*�^�;�P\j:��q�T�	~��s��
�[D��k�~��գ��'թ��̮%�9�[Nd�j\Ȏ	X"QuW�l��5��9��yk+��Va�}�D�\����*�J) ?��oOG����lhջ��m�0l]?��
R��XEG$����x�gޗ2�k���<1ӧ筪F|J���δ8�Jb�.$������ѳ��2l�?2�\�k��6�����`�	��qEG����9�X%�7����V
�-qu29TМ��˃�;��>n�RMI3q����'�]�q�(����i�� g-��%,@v��) ��- ����cUs� ^�gj�#�3�nw����[<IR�b��w�֊�m�@���T��g-���3�忖cEW����Jh��z4R,s�\䴐�������6m��V�/u����6�R���_�0D=���U�y�;*E�xz�9Az�j�k�_Vk�P��l]C
J&�1Z
�V5���>�<��Ǆ�����UmM�ӏ5j�	����$���D�:>�=S]������B	|��8�G�1��v\�ߒ�/f���m\x�տ�M��¦w9T���~��8'F�b^Y��W�(h�Gqbg{���@����2�f79�K*H�w�}����w��,�������~Q_�UJA<���3�d]-)��fs���t���i	Z�*�E_s�K�^��`�z��&�F,ܫ��X�#>����#�-��,Q�b��3�io���|!�[��JDD�j���@�	p�ߋnP�9zo�B&��ƗV������{ϿۊE%(��è�Hl,��Y������>�_��Y��8��c᳂�ѝjm��pݥfb�����ԡ����WF�Զy=S��E�M�5�D���h�|Q��ԯ�v?�U���D��RO2!R-�m�%V�~ֶ�����<׍��K���7;Ҟ�LUX�JJ�2q`��ӊ6r�U|j9ӧJ�^e#=t�`a�;7�y�|��m�=�d�5ڔ��JjiXF�>�z?!��G�S�'HG֠�H$-p�+�V_l7:=�Su4r�E�w-s ��Pc��gzn^C�Zw9��=����gE�H����8�:��m@�g�֪�6Ɏ�>֛z��(V_��e�|�N��jvc�[Ǡ�ϼ��W)� ��ؓ�����M?R(�$�>�rT?9��Gh�兩F�QҲ�J0�x�"�l�o��l�w�M��h�	�|��)��/��縥@J�rDyi���؍���T0ך���c�g�[���OƏ�,�t(�k����P� s͖���c��Ղ�9T��Ol����%�;dh��R� ����l���M��4%�7J�w����b�]�� ��UMpx"��r�@��e�g��V�x�,��[f`}�Dp�	��L�"�jX�vV�EQ�$�1����}C
�[�_�G ���/�eѕ/W���_Ds6�7;��V��9�2���{">`�4k�2uj�a�~4�0�v�Ҩ5uYf.S`��B�� �|�]��u��ў�G����@�w8���s�>
HAs�Ʊ�|bhe���A��\���񑈘2�Z������B�7�N��bV
0Q�J��:�;�m0^�����&�[��{q+Z;;�!FMJB�%q-oZJ$������E�Yu��f
��Evm�V�ܣ@�N�z�2��*y�.3e̺��I��m�qV�>���@��Z�]98p]ؑ��a�v�k�h>��'H��̈���;mq����tF'8u�嘎e,���b�_֑�ҩE��i#�Q�o��f�v+Q�[d��8�o <�u�%͈�1��v�,�U���Si Ю�0�"�	X7�Y�Mb�����J\Z�Ap����a��p�R�2�]�ݍ-�!݈�Z��M�������v?���Nr8`>V_'��P&60#HvX��l:������>3u��e�)E�"�^�R�6�8�%?�.>�?�B�j�$~|:�a�*U0�#2�o5�z1jԿ�fQ�����喱:buu�B��0-L��+�U�P�s����R?��==�T�z1Y�u�B���4�p�"�
2VQ�`o4��0����x�gkeeA.��M��S�Qq�Y\�n��1~��W&e����Z*xr�.�(�F��p&8 zFg�����$��9�k�{��J�ZyRA���:@ޚ�����\o��m�\L?y͋�(0|�H�NvX7�?�����듀V<֣��ʷ��(!�ʃI��Abny޽m\��"�����۠E6��Ȉ�����b�*�5WЌl����v �����S����5>����l�?�<T�{GK���������VA�B�L$S�9��z���2����E�Y �bR�4�(����#�
A�er[�ЬW�h&���Wl���< 9t���W�i�3^���W=9�o�Qa�@k��Y[���ZHa��@�i��*V*�KӒ��Fk����da^��ݲ���a���꽘���ا�͵V���TC^�iv�{F�e7#�CkF�ΔG��S�$k3�a�s�W�ū�b����o^`.��m��*N|*Fo���^n!L�A�����S:{���6�0�+�����՝DXCn�W���H4CD��˟&�q�X#�3�L ��ѻL�����]5+���@�K���V$/���Z��9��=�<�	�D0��U%����f��������ą�:.p>�]2�u5�����Ub�#�1r�yE�e��V@��.���?Ct�֋�a�W&�ȏ?>�z{I g��s�
���+�*S�~�2�]i4���s
co&E6�Lr+�ξ~��bن[��m۞�[�q�ʥ���W���Cu��F�gZ>-�% �&�I��g:��lS ���H)���ؽ��^�����p��}Zx���o�����;mu\�����j[����q��H��.j��&�z��SЋ.��U����v,Dk�!�p�WYs�3�G��<Sj�֜5\_h�H3]C,���Q�Um�kћX�1w���?�K�-y7i��Y?�%�"����eLe���K�
�{өe��E�A�8�[(O�&�G��p�d~]����Ia*ӱ���Xm���t8�E��44T��=�t���y���Hq�2��fJG5�(cJvZm���<g��5CU22=���O^�<���8,�3�N%�f���_�n�b�͍�Ҝ�3W*i��-��I�Duc�V�PB����'�C��ځ0�h=��Cf��D�^Y���2({��ć��荕*�A��+�YJ�C������ԨR��m��[� ���� �1�L���y��=��[G���5l�{�v�r��f�x�	�������V,��m-�Q�G��ƍ��!�+zNR��i�#�1Xﻕ�b)8��4d1�UԨ�4nWp���K�rg{!�i��qǱӈhb|�޴qW������L��'P��h���$��+��~�?�cU��:��h)��������86"a���_�@��z���tM�d�8{��&W���h������.1�9*�*�-�	�{)H^/�@&���N~eLM�m����*��&��F�����984�3!�	~�"H�/�*ge��dN(_㬢�t�[G���N�0��C�lD)���X �kS�V���+�ta�\H��Đ���*t4ϟ����_�m9��]�F=�B�o�jL8x)����
7���p��Y !w�@뵐kIS��
Lk���F�/�#]�6�`���{|�t'X��r$�\���g��G�:z�_����&�j|����(ր�朌��ĵ.x%�_5�Xvz�b+00P���?�ozkY��"���nv���"��R��������QC��~�ѩ[$^*I�F������6'֮�_�UZd��vg���>����3!SSfC�
��*��h�����uÑ�#�i�/���3����y�!�����=�����I�H�2��|�Ӝ�68iqd�J!�;UQ��Wq���z�MO�I	Ͼ����|���+;����z�ߝ<n����ܛ}�)�>��Ͻ����ǒI����L���<$�ɩ�gc�c�"ۤ%[R5y�kj�<��/)�H�уG���T���Y���������<�Q�"!��(�0Z<�Y�A�}�֚�����w%�2z�U� �"�cA��FK"uf����KYj��u��swI�6�P�;٣E��I�����i73
9X�7���zl�c?��ԝ��+5c	n���i=ޥ8�S��{�����f��.r��|�q�pb����V������j�k�Gq).��)^ܡ@���+ŭ��;Ŋ(R܃��Hp,8������?�X,��'sf��=3��Ü�tK��f��q�#Y��8^�^ƙ�!�g��	}xޛ�[���P�f烷ֽ�>�Kا�N�����#nOc_����ͣz�����! F�����U��;�ɵ�ͳ�%��)�Yi�<���A����O�q��x��ڎsKM���/NLG{��j�8g����x��~<.���q�I��!��Ǐ��q2��&�{����C�$7�H���.<���:�U�������$SK��H����z�<ml��:�0j)�g�̚&�����dԼݢJ��''�"в�g2s�$�������0uas.�ZNѩBM>�����-sD"��Ik��BLv�N���^j����wX<ƭ��R/����m1�����8X?�p���c���b�i ���>c��l��9����T�__��1z��@�0!x�3�?Yc�%����� ݜ����WO��iD5p�wtc�	H��tA��c�ػ��꘯� ��ף�f�.�h��k��]��?@%,��w�![{�v����jŚ��I+�yl�.k/gD��*�y��r�]a��&�ы�o��
�SZy��.��N��v�1���<��|��5�Ѝ���fszVz�{-5$����WT�2S�%>�MV*���ݯ�"޳QC�@Gx���<��;�tO��x![4z:<Q=@���4�N}z ���y���IZ#�%������(;"��ᮔ����!-��S�T!�I��iY�,8��*�&ꥦ{hY�{Ep/��i�P��hM{���.�S��W_�(
�"���r��V=��wc��w�E3�y�ڠ���{D�X1}Y(Yj;5�����<oҽ*�Zev�Q��c^�5ѱ�����]���,Y���� v�"��1�t�Z�e�~u��Ja'�k��ح���W¯h�q�6Gz�H���C"E�=�`��<�k�5��z#���hr�z�ln��Fp=����8��O �7m����-��EI����@�����~���@f��𸗭�+%�|����fXr�s�S���=(D�rcQw�Z�!S�h�uH��~`����|�߅`�b<������}ȫ��	|��2IyGӉC���~�0�#Q��U��1�P����=Z�)51���J󖞮����8i-�쥃��:��p��5�5S��=x#��h��}�/�:*���l����z<_���f�G ��/$+���_�~�,`��k����`<ǎr����T��~��mG��tš���S0zn��p(���#�w��� ��ɫ��J�Os�ǚ��e���0�&�����i��sz��Vs?��Mw����7X%�5m�D�,�u�2�^�b�ى���EB�LXǺ�:E&�.�-Ƥ�mW5!�sR� 5�M���5�%~��ƕ�����n,FwŠF5������u_��:	�<���S��^�@�<�`��NN����tXR�x�I�t���p�.�1��d_D�K'�`ǥ��/�����9�?MP.w��u��H%���4��,VF]�򦂹��NQ��$�}����{�f�~��I_k��r.��<����*����#�/���<�Cs]�����B���������4wF�g�P��P�l9�Px"*y;�+�d:r5�O��d�gn*}A���o����KB����;��4d|e�.*�|����=}L�vb� M�I��u �sp�����;P^WmϽt�&�KL&d��x��{�ZWk�5ʼ@��+	����qݶ%k�d���:<��F�>c�4������#��R4���֪|1��CMַA�T$l���p�z����5i����U��n�_.fk;s��W�.� ��6br�S��y*#B�9B��z�,�QV�����Ũ�l��/>�����a��?�}�Fy��O�j��Y�&K������˨B�4��zk�9�s��B8a�'?����f|����dZn���H�G];e�F��'�&Udp@�(ͣ�"��LP��v��a�_�~?��`������W�v��b��.�;���$���}�+ΣŵA�-Xĥ&!+��%B���%�68����\1����)�Ë��ɞr���~�%1z<�K���J:꾽�	���9�����q�Yl��cH$�\��%�݃5&8�rg�����H{�]�P�_�O��b����uQ��b��f5��3Xy%��"��"a'l�2�����ܗs�-n-T3#��C���ֆ'����J�Z.�B�ō��oB9�a�h���s�}X�a8v��Us86�"|�2��}n�����)�c�\?�75�|����/:��\J2�����=av��sϫ��_�UV�����̸��䤵����}oQK+&g�bV�պX�18�J:��W�C��`<��W0N:�����*��7�v�q���b��W��e��� =m����x��|;#��M�H��<�M����`�uɎ���*��[E��苤��YΊ�X�8i���T⏧�����-�1��P���ȷ�C���s�_?u���%<5�="�������p�Į��qa�1����G:g��:�s�s̬V��!&�o)��I 7�^�ɵ���c�c$�@E\F��Z ���-E���C�X��g��׭e�3|Ve6#�0%)�|��|�$Xk��鈟3b�)�ex?`p.|�����V�H��������.R�oV=<+���cϧ�=��ү�{���~F�gb�8�*��Q�����z�O˕�`��?/�Ŭ�Nb�o���m��6�p�(0������D�ڹ� �,g�F�Q2���D���T2�uÿ�U_�V�ĵ*O�Ì�8�Aϸ�.�Z��_�R�6���m����?}^�X|�uЇ��4�.�z�-�݈d�8���n�3=	�p��Mo��o-��U�V�!����'W[��a��a�=��P\�ז~z𹷞�z���ձU"�0�ܠ��b9Q[�c ��о_���9h�w�ˬ����h��O��*�����(Z��wj���>yG=>UR���s����?���tp�Q��̭�p� �[����YWR���๞nݿx���ܥ͓h?�3�`�$k#KCo��R�P����3�}Jy���eJy�u��ж��nѿ��.��_X�Z`�Lp�����L����9����r�V�/R�ͨe��QՂ����"�zMY�����F't�X���4�m�O,Z��=�T�	eB������G��`�����j������V��X^�z�9?�׽������{������hw+��s~���8��q����cܻ�aV���c�橨��Z���X��^y��#���R֭�q%w��$]�Sq��ʥUk�GiW��q�i�4N����o`�C�a|�1�Z��N����l�VJ���1^��<2�`�ͅg��)~�2���)��|�9G�,\7A���T+���˾�Nb��:��I�,ꐲW�F����>9Π�w��
��5�h���Ö�ߥ0���i�����7�9�@�B>y���$��K�f.��A�4��R�_<`q{�����w����
�Z�hg�F oD�L� ��}lw���q�Piګ��m� �@���w�j|CWNW.Ff�=?�J�n�L1̜C5�Qҕ�)�L���P�L���>�/!���`߂�/i-�r5���{	�_M-���UWn&tڪ�{N0�{^����A����$�&�|�mǌ&��;��cky��,B�h����������/� ����y�F"�g!ϣ�O�1�����w��\�)ˈL�A��K�z��-��`[*Q��o�~���L��#*�܅L���Hn��h�+��j|\��~J -�*��u�#Kk	CD���W7�o%��2�W${J���Rir��Ϗ�ρQ�V��?�:�}h�&m��E�R׮}��0l�w�k���������j�Ct��P�U3��-^
`\ǧ@�/�J}�-�`C���g�^s��a�=��锈�^L������x��j�m�GM�� 6���veU»��t�)�<�:�~� ދN���=E�?5��|�������g<H���o�}"���lsn?��2M'�,T�Lj�*�KZ(������Qk�_�4o��T���� ͭ��]��4݌��t�������߭����I��sC��d���s�+����D{2��h q�1��|���t��?���1��g ����_T{�+��&�%�>�T䳄����b#���}�¿�E��W�"�ʜ	`R���Y|� �%+\�&In"p5��`��_���E�i�&X�] ��(��l�5p�v2$2����1��B�zq��C�Bʨٽf�pE��l�,�}��z�qR�6��)v����VF�=q��?�k����k��$�S��:�D� �o!��n�{�Q�c���)[<�!�S>�_�h��)��kZ��~�Ńs�3HțȂi���?˼�DR���P�\D��0�Z�nj;���:���	}�>`�̽Đ�g&�|a�����A�[g��FSċ��z��|Z�;�A���җox�һY#ݤ�Q~!ufy�Sg�8��e����{�oV�#.ش��2�4�v��j5�p����U<`2jx�W���EsT��j���/�f����{��ת3��������M��Ċ��<g��� �B=L5C��4��+m8���~��7Gʖ��{��5QO� f.n��X�Nx<��	ѫ�I��� ��%��]'��,��]��J
f.m��5�}{��s~��h��[��V-7�/���G;� �;l�@����I��п�0�[w ��#tgw��&��U�k�s�A��6z�b*ujy����>�YQu}��s�:��ϻ���B���J��`:�α7�g���;g����Z4ϳI��k���,�󫬂�o������V�_�I_�[;n�O�g.&Ǉ-v��qJ�E�g��a�� ���t���ҫ�����h���?��K]�^�⯠z�ԏ"�[#.m�v�H�����$f}ȏ�N8��C�:M%h�31���*w�<o�s�)�����K��@G�2�g�fx?����~��Fo�Q���s�~���2�*��P�O��ُ=P4���x�c�P��0�݄Px��@Op15�>g*��!h#�L�t���`�gz��uڳ�2��/�ޯ�~'���|��$�ZAfd?�w�@�"�«!���^ua�\3C59~��p2�J�!h�I���8q	+�x%��\��������rd+s���A�_��3OĈWׇ�����dmW?��z(羋�#כ �T�H��\��E�&�+�K��Je,��81ĿԜ}5�u����~�i�z�I?`�߻��{�L`��T�6ܴ�Ξ��0�C jq\�B9!��D��/V��l¯&W�1��D�3��;8�tsN{n'�{��^��{�G��}��wr��}/D�����q��%[�J���Oz��fީǰ�eF��^l���)6D6�#!4<��:س��l�y~��~Q�����ON���ӿ9���V�WY�����B����
C�d��g)�P�r>�%���&$�N�zCH	&��BOpGe�sθN罎:�n��0��j3������x�XZ����G�~?���5b>Q��ӽ��;P����*@�n;*�Q��gϴ����8W�<�_ax.ɀ��3�m�a�������Z�v� ��r���&V���S�$�Z���Ӡ!�c�W$�'�t�ⴺ+��Z&����4���׍�Ar��W�J�z�X��L6��^1>�t����4��C���3esW ā��R
G��Ӷ�k3��nRq� ��P*�������WVr5���V�O�7)���yk�+�����sy>��iѿ�7��ĿK�
�6t���Kj5I���c^�F�U���zv+%�/�6���:�94�co�+�>ϊ�3��hZl�cB]IHnv��8-מ9˼�����1��T��eݛ8�y��eX~��>θMw�en�?͍�`�y9b�Xc��"|�`�����1'��1K������D���5H����ĀU1���\՞xj��g��'v=�>�;zȟx�~�>��8���Ƹm%j�j*�twI�~���enV4/(�_|h��Kz>�~����x�
8�8�j@l��=7���Q]�%ɣ~�5�����K>̫��B�֕�d���Սה�3>��9��FČ�Q>��-��o���{'�z���PM�\�˪� ���Q��U�e:�ڀm����^Wϵ��.o�מ�����'|�*e��]X�֟� �j�o��!��ˁC�Z/�J�Fe;9\�#jGy��7���=�#���GY�G�S�����Lԟ%h:/���R|�g��%i�ǩ�Q.w)�������!Q���#�%	��y���CN[���� S�ޝTS)Y��� �K�����b��&P� 3�<�����i}K��qjt�����PD�&G��	�VE��|�[�&� p/��H�J���GG�}�)��pe&o�.�������?n���<���b�K��I�ɛ1�zd\�������&��\���Ӻ��k�F	�	����{���9�c��g�:�-ǐ��#4�^�+q��z��,Q�[\+�л�M�C�M���XXpV4%��?�bTҼ�ఙ�0��Ⴀ��
�!� �J!\u�ٟԋ�K���j�u��Qw��e����2w��^�8{�¯�ƚ��@J3'}~�{g�@ݵu��2{��8-uu�3Ӱ�Ͱ���E�����'§;���F��$%:_d�w��8���sD�A�i���Ht.�Z����a^��2��q�7m��j�N�UΫ�Pc��ԓɥ��4���b��=��C4����'�\��8�C�Z�N���k샴��r�ң!k�����~@^���=�^+*�!�?f�c��f�8�u�[�(���$b;	��E<�U��ư�X��4��A������n�۲Zz�������qC�%d:v���D?B�lH�[1�����Ե�ǽ�6z ����#���O~�={�CԘ��F�b8J�z���}	��;V�lN���<���1�8]�OJ���i_*�xl��K���%�����P���ˀ�'�0����A[F�>�P�thl"_j�^�5��d�@��%kS��N���*3��s�˵�g�U���u�L�Zf&g���������W��ѢM p3p����4��=����W��`�ea	C.��og��<-��nV^�L�KA�
*Y��z��9��y���T</��㗜��R^j�~5HO�ѣc�����S&�}���+As$�QFk�8o�j[[�K�<��ǳz���#��^]߀W�!^�dC�m��"��}��o��=�m!��)��7]��.����b?�Ex���%ͫ]@ս�4OC�k����Q��#Ղaf�l��j�����i���r[f㻱4f��o\R�,C/�<���K�'�6��C,'G��Q5
�z�.D�r�1���H�QoS���bєP-�u�%�o���������iX����]c9gTB��~A�8����l�p�z��s:H����g��#]-��WP�Џ�0�L��u�~��'����!�*�4d��'���\̏�"��(���~��\��tuQ<�8�l@|���<ʖϼ�Ur�i�Z�zC:D�Ѩ��̰``����!>F5
���0zX����X��s����U�,��;bE2�ep�m
m.���BE	�*s��y�?��%R�	�uG;rK�!���7 ܵ���XQ��*5� ������Ab���SY�';k�2l۽��m�/����\��7�`p@*%[�X��
�i�zQ��E�6��Ùe.&$����#�W������"�y�h=�����c	�E7.,�r��0�WU�Du�� 9��x4��Ll/���=_�u�<�P"Z'�7��z�ľ�SdW�uA�J8�|��G���u{�r~L��N�0�ю7$,z0ٷy�G@�[)�,I-�y�%����s�����$��ˆ���	��t줢l�Ƃ�S����LHGn��`�7;�?�jN���X+��:�����0O��B�;9�3�� �-�ubA��Dĕ=0�y�aD��m��q�.��1$(1�����;�aU ��-Fm�Lo^E,�9d����u�4U>3���e,m�i�W����Bȴ9������tH35���s82ѫ�w�IгY0��Ƌ�b׸���y���{�R�!�]hY��?�c���j%x��ɢ�X��qd�~�}2$Y��~�Ve
��I��̙
���1>���?��_���p�h�N�Э�lV1�$P}>��u��j�A����<�P5 g0�yKsb���{��ΥB�0�g�G�Ф�f��d�% )��#�{��+�e��w�:���(�J�M��[�µ@�tY����ĕ��ٵ�ֲcpT���F�{D4@�s�� ��˔>�P���	��.$�@.�P���6*�
��amS]��5Ϲ+���|��� -�:�p�`C�F���Ke��,���w�|
�9��`�r��;��5�j�j�v�:�n���9Ȉ;</`��ޯ���������=�7��;����U���~e�!E�Q�*.�N��H�Cn��@�D��_>���7���N�~/+�t��.�Jg��Op�Y�U��d�$Ҫ�]��{m]�	{/zߚ���~C��]u����-�E�wX�C@NH�#���xPz�H�OW"5tW	:]?4�B�/�#V)��6D�l�������k���A5F|�3O�Y��w$t#����۷�n�&�cz���xk�4�X.�GR�%O�>|�%��qt1��m8Z�����غl2}}Ard��+\P��y�8Rg��仇��9H���� �TB"&�q��?��E�����I�������d�>�r����ۘ�8�7X��:~s�R#���8 �m�B��Ï㸛D�ш%��^�������b&리&[����o]P�锜Q���X���Y���jZ��# ��=��E�/�Hu��3�N�%�e��}q�V������r GY���Z�GV��_� �pS�)I���Ed!�^�r3C����pX���t��G�A�rN �;����Y�"l�`#��KT{�!�� ����YEq��v0y�;��*�_F��7M.��	�{Ӫ��)�B$p���]n�\4>�_o��a��=�6~�ZY�`!���L�0h)��n�4�\8w5����:�mb�z\�ӆv�;�'cIYzt^P9[7�f�zѷ��͢?9d�o���Øqf��v�{\9O	+�{fb���T�����^��R���s��Lp����t֢s�����V���",`���ޏ��Q�'Y4T�5���N{`�,�����=@��~*�{JL������7\>�ye)9�M��%q��0RAI�.o؜�v�l���P+����bbK�X@eh��,0�6��,rr��Tvs���補��jA�:�V����"#qCy�?V7�a	�q\��Ez~�|P6�>Y�e� n��hx!�c8���S�+>i�=)�T����oof��W��W
:����}-��њ̪���w�0F�-�h�Wp�5����?�%I�0�R�?J���FW����	�}��ۡD��gR��dC���d�P=�Z�G�H�����'Ҏ3���H歎��&�5)���D����m�-������uqa��!�:���,���?8��E9O/$�A�hXgMݸ_�� ��{���OŽdퟫ�6]+����_��`�+ŇA�{w��j���⏡��x�sG����;��"�qCّ���(_#��DِG'���Z��*�t�ؚ
Mf�Q�3ڴO<�fw��x�"kBΔE���JQ ��Kk���FB/�L�>��&���#��e�o���uܼg��������,��ݢc(��x��pp���(���R?Kﱟ L���	������5�p��C�Wu��1��Yj+�'��)�ca�l�9�?��zne��C���ֱ��y���@��ue�)�����k��r�y�q~��ReE²� 8B�<����<������ܵ1��p/�\�	HY)=��.~�>��D���k뀈��Ӱ��t�q�٩���-�揼za��G��'�V����5������;����H�h3OVY��/>	�1!5ȅXńo\Z��Ё��KNI�Zƕ(�*.����#��r�� �J�t4��L�2��;����W��5h}�p��%����f���R��ʀd����I�&R���š��V�ɀ�5
e)����(M��W{�Z=�*�	7,�g�o�ĵ��yI��ʝ��i�p��-�B�bܶ&��ɰUw�2��']k�	I"�W�H+�f�v��Q(��E��'У!�%�Y��x�K��y�k�F%�EO>?&P�ٹ>�[�c�a�Jdp�ܓ,�zm������+�3��[h�p?��w�1�}ں��o�d����_Ы�"G?���N��D� #�ȸ
ʈ#D?L�R+�m�Z���o�K;�*9C��"m�ƻm)!E�V���mv:-}�ĘeT,rZFHeq׫Β�n)�b}Ǻ&zD�k>(����̫��x�c����d����370 �i����S�	ě9��!��~/8��x_�����Z���7=LC�r��1��%�<�c 6�*�3]�)��6~[9Uw+��`"�ZĬ�8������ɦ,+�JM�髚t�i˱�dC��m�_���o	��_o���p�h_Î�3�j�g�g�AX+S5�<^/�3�;0�2�(]�\��y��q�<��O�� ����o1,h:|EB���Q����o�] �8��ݐ�U�k���Mm������!����>f4m^��0E���.�����E�P��Iυ�q�Yq�Y{�?�9�lb�L�H~l!�f	c�e^;9L���rR$�K#N� ��'�+E�LT��$O�݅�S�ppH{�gw	��Q#nB4���!\�F6�F6y�Dp�M�`���Og���S�0���E��:�<1���۱Nx����g��(��GmK$��z�&Do�u�w(����%��EĈ^ܒ��J�����^s��G}�ZWU��,1�9�)��'rpG��g�)MH{E��t�Ʊ��j��{���
X�Q�Tx(�����?S�����=�{bt��BkS��?�M:�7���-���k�T��a:���|'��B���G_>���鏔�ob���u���)+��R�D�fꑅ���&��Y �Z8L	L�>b���<�y>�("v�@�W��ќ�Z>�0���@�.R�āc�C�	uW�k�p0d��=,��\�U��I��?�LR��CR�tŃ�υ�m>�zs<�X�`���^�\Kxq]�3�-TEG��L�q�a��y��k� 8�_�w��,���V҅::EIz��]rm��Eπ
�B���ӟ�.K�v{*������=�6�i���q.C_������ߠ#�2���"^csg������3�K'�sE:�vi��bO+��il���,J�n>����M#W�>'�U�y��P}U�y�N�m�B�Q�����2��K�{,s��Vd���ƴlC�w�-�8n>�3DSPN���?��
^Y2�og�xqz�d戲��]�if��f�o�!����N�+�.Nժ���H!�������<�ڟZR^g�A�D�?�[M>}�.��ș�17tF���u����"q9��Մ��k��5�ި�i�]�=�q:<g�\������	�j6���@���U����c�
`z����%�ݷ<�EΠH��~�%n�'���J�{�v�0�v�Wٻ�:"�Qh�e��̼'�]��=�M��������n��-ޏ\E/�V�����Q�I	2d������t}�8au�z"��.��,� (`x�y��5�ϰ�����Z_���r*-K������<����rq���>��|p���������Zj����ƥ����e|<�tG'�maH<��o��ۄh�"'��6�{O�����U�^'څ�W�����Ǻ;_ݻ��B� ��0	��Ow��O� Yl��ǳ�Ɍ��x�9d��l�`�\6
\�{��@���m�XR~�ӑ��{Y���U���ҿX�r��Ϗ���C�]m{������T��&*J+8�|Jn�͌@��ϸ;'����x'k�u'2};(pIᏼdl�M)�YE~1;�%��� [?�"����d�7���w_\��,oK+�m_I)�Ԍ]JFD.V��<�
I��u�E�!��p�?�{����Z׽A�VS?n{������e��43���*!��� 0`�RS��a���𣚻}�]�2A�=����w*\s�U��HfR2�y�K8��X~,�Iҩ�T#Z6��Y�k��S���U{4���Ɍ��ޤR��~J�M��NS�`��.����i����W#���� KsI��s�^}�ռ72����������xU�`�T��b�2c��78����2�bmy��2��2z����=����bs�i�ޱ��f�t~�k��޹�L�ӘJ��)%�|+�����,�ݥ�/a�.�G6
)�C}�޲|G�ز)�R����kf>&Ew:��}�<��O����m-\��y]��������i��z�l���H�/<���4߼�p��&���m=�`]���-�R��0T�~{���"1:���-)
A���3e{�1Gz� ��,2��u~�7f� ��gX����Q�,���{��4p�	��a�R�������-��Mt ���f�ĝ�r�h�[n�!*;�inn4
��R괸K>�
�|��v���R��U�x�?݁�����A�%��&�d&�(ğ��_+r���Z��)�G�@r���H�<T��B�h�{KhY8t�RcLҍj�-�G�HsLp��[
��ѺF�H8�n[��Խ[�٭��=	@�|_�9�����H�8#66
��]h�F8!�H�'R��ƺV��z�OT�UKT��23��W�P���-�����U;f�
=�k�:�M���$m�lAdP"u��u��ۍo���f��*i&5�sٳ,|����ǲ���������)=�ȕfw������'��pw-Z1�Fg	�}�M0�E�Y����0�I~l$1� &�#@8��;���Xy�wq��p�i��ta���Ӻ���V_�ݺ;��ꀤ{��+�ɢ��x�V+�`d!�d�G3Ꮍy�X��'���M��ϋ�ʂ��c��>�;�$j|� �|r���M������$�Z{��"��`G�I�S���Ώc�u�@������2��/i�v��T�w}�G�k<�!��F�����I^�chO^�ϥ���P������{C5+�7�3�e��0��bla��p5�Ϋ��ZR�����<~�`����h-�S:p;դt_p��RUf<1�blB�ďP�5\������*�����F7\�rh���~a�>jey�u#�zJl"�ڠ&����J.ɠ��.�=�Pg��3h�cU�����y��ZQn��[},��[Ӳ��1Ղ[��ZO=���(ahu���*��A���uҀ�k�I���BW�ǉ=���RaQ����!23���B�G���Uf^܌���F���5�	��"���U�������R�N(�=%�������f�EB�/k�^XU�%�L�+~dϏG����@=�3w�3�7�i^eK�k�s�@�$�YDdvѡ��5��g�lL���%���EVG#���O>.�s�i�,����:p(�r���[�}��y`�^ß�#ap�ǳ<�V�ysE���`�b�b��ħȶ���1T��B]��H��*j% ��鯨�(�so;�����'���*�M5 V�(0h(ϓ�P2�/�}�}[�7��B�!�[��+W�����t<����ֺ���nq�a�f��,�u�{�������zl8�Ǔ��eƴ�oȐ�����j�髆��c� >�E���uZX�1R ���C)˫���	�5�&\kQ΋
����������-?J[ P>�7�`�.�\O�"y������z�n16�&��U9���mH��������x7��q������j( Ӹ=�_MJu��,���nG+�)!��֙G��|=�w�-��R00����;�l�s���
X
�-�ǎ����`+T*��푷y��/?FM�A�F��Q�.�+����%�g�G��r6�닚#��{{��X#�Mt�,���k��AEƠб�Cx4}����B���C��s�.L�[6L�2Ӈ��k��6�k�k+(�i_��֟Į�(�G{]V|����`8W����"��+����e�Qp�YՅ��v����}32�Nܵ?�2����Q�>���Z.@�������f�+ׇ���R�6t�:e��EUA��,���I[����N��C�\����B�r�����r&\�2��o{�qz�I�Qi�b#�C��C��+e�u\����%Г�p��IbmI��$�V$���1�`j�i�_���ω����&<.{��(+}�8�잢���]��ڋ���VbwL'd�uv"C~�wrq2Hw���'��t4UJ�z-d��K\�Em�zm��[
�@�%R�xB��|+bq�q�Z����'�����K��Y��]���_��:�;��+��[�6����|�����_�I8�RZZ�O��5>�ӿ��m�ͺ�U�� �:툨�����ɒ-��j�(�'O{��d4-�gY�2��e����?.i��e	޵�(��mבQ��.˼��rH�dB>��>��sB:n
��[�2^��s�GA��*2���/"�6̀@D�N㵥j����r�������m��i��8@,����ǭ���k���fwK�o�?I��P{��KB:T���������ǻ�s:B�~~�Ε���L�}ۼjU�[x��:�
�J�O:��!�N�jm:�}�p���\���Q��CP�-�Y5T&�O��H^�n�88��I�Em�|�9n�AfD���Wi�7�P�w$#�Ѝ�t�I�Jb��u�4o>~�de[v���{a �
aƍ��� �B�sq�}�.�&$.x��@ÓȥgkU����<�@�����"��1Zn�1���9�48Q�@�@�ۉ�����S����;��#�Y{S�?�q��['GF��ɾ������7%��p3Q���͢�-�������!ެH���P��H�ͤ�o�+qz�߮�����6�c6ت���`�N��l��𠶦j�nH�Ns�	��^��e#��(i��BX��mx�E�2��-���T���U���&���E�>��٤�چ]��B��u%O�ˮ�(�:f����a�H������NDVڬ�N�Ͱ����;�Eת;E��O����X�w����-��Wc܊]-�q�%���7n��\r�Vp��\/�U��t}kd
����!�g�.�9������u>m��V��(���ߺ�c� �5w�jҟ���}�o%y�[��}*�SS��N�uG��H���,���,ƺ5����7����/z�js��sv��xQ��*�D2�ѿ~t�n�x��-�	\���Al]� v�4���p�s�D4�j��7}�zy<������^&Xp�e�s<(H�qH<�b���E~�8P��#�S�G�� �y;�#�^��{1L�~�z*x�s��Pz��CJ³�\�y�V����5��8�$���j*��m��cV�� �#�7�B(*򸿳R�D��(q.���K�'y�uZ�:F�!p��Ӡ�2��M6[���70@v�҅�&v;�14x�����I��۩�Yg�����Pw*'�<���~�n-	E]M��1�F!O�X�S����4���wt�����x'r?D��`�C�NEzX�6_�r��R;0�9����^A.�T[QOp| }D)�/w�u}\������.�"<1�% �g'M�=%�q�B�J�ut���E����Z�S4�1�����&��0lj�>�L}�Gw��
]���3�Bsiy��, �4~�	-�遅���U�h������[.DHC}N��\a3K�94ͺ���)$�M�_ݪ����@n�ޛv�c�YKi�+R��e�Eͳ!{'�~m��kf����=(�����s�:�j��*�$D;=��Z�4˰ȿ�V*m{�X�
}�'d}�Y7�~yn{���*q-`�V���
���[�����֢��q\�v�OW�5��Y�j}�?5��Y:O��
��y~��5�T�����L����� iÚ��L�����v�t��;�r��QF�_o��f�1��>�U&Z�0X�bB���ˈd�ʹ7�[�\a��5�� Шg.98.$���K��4���T��3�[,Kt��o��<K//�!�3����0�
!�a|��C���+� f���Qf�;kM�Lj)��ȫ��	��R{/3~�u��0[��� +��\Kî�֙�*._����6�1�=0��;���
�Pw��t$T��+��ؿ
�߮K�����
����mi������[��FZ�n��i�t�n�7��}�9￯�k�����~��1�<��b\�#$��|�Ja���h=vi�[!���N�SwMہc�4���P�F_���yK~P&�e�c%L��Ҵ)�ŋE�e�5Ɓ�_�Ĺ2B�'��f����g�^��G�Ao�d�y���"�oj9�4W��Y��YI����g�(2��:��L����o@�XD@�㗳�J<T�t!�u�Z��p:*/��z)�P�����~��zЍ�%��]���8�C��OD hB'z˧a��Ҿ~ִͺh�5+�3���nb��C�ÿ�\c�BR飼��Q,�_GۺE|��Kc���sv���ǮXk�_0�j��bD����q��q��]��~�F~Uݯ�K-\Ƨz�*�C�5nN}H�Ղ��Ɵ�磔���e
�ͳ$hi�2S���9^���gw�q	~�.�E��	n�v��'�z��$�.�a��ϓ�LL`��k�^Q����������H(�^ٔ�м�W�������E~�ɽ!�(:�"�����`�~��D��	�Ġ���{%�;b$+܉���µԦ8%�.IL�j�O�H���(J.ۯ%����?Me?�������h�u!�����s՞o8�9H�-dT5utЉ嗞D;��(���Jy6u�b����J8Lӑ����I�￯�r�쏺�IC��N3���׏�|�xc�Q��`�
�n�6�H��Eid�`|���*��	[6��)d�`����� ���+��{���F��|�><�B����6W���~�%y�ȱRn�n +����^?a�p�`� �f��q�&�D��ݥ3;�9?B�*z�Q��}m�k��H�������C�51!��=��v�g�xcj�{Xhy7�< �Zfg��ڗIk�\e�e���\Z�������=e^9r!#q�7d%��鷊��!k��
K��B���63�°��r{��r��+��g�������$y�ʱ[�^8�."�s��_�`!�ЇI�����,��Uô�=��dH�r��e�����M�3km^�h%gB�yAB7�ɰ��-�2tt:�U��ݬ�io��}u�+�����Nh��o073Q�R�I	P��ḃq�z�$��d���В��q�Ey`=�RHs/q�S՛W�K�dAƈ�K�uM�T��"��kJ8��� �:��9��_�>�K{�u"�fA���]S%�%|�Q٥���s���������u�ml�rݱ��Qo"Jy|�1BR��[�F�<�ݭ��cΚ��d<M���P�?~�
�����������u?uH3�RR�ѯH҂ϱ�Y�H{�JMI!Y#�����<sD�n�N���!Ѳs�� ��~{��ԖP��a~��q>k�������ts�� �^L�ZJ���'���Ĭ�;�[xIk�yP���"�U|�L_��o�Q�=b�Lm�D^�Er{���U,u۷BR���'�_�W��3�+$���
�b:����zirf���)��-�$�!:O��Z���yc��k��C�1g������W�Ԍ�����
7�
Igng��G���=~��O�#m�j��~f��o�8l#���B~}���� PE�~���J���c�tӴ_Od����
��VU���q���O���C�ܨ`�{��*H�E����:�^��淪 Ey����˩�4�Wh��s.
rx�4+x}�΢yq�E<r���;�9�Ec���{�
:	�e���ᚺ<|;(q�Ӽ������O%�[��gbbI ^�Rnn�"�H+�o�Ƌ�� �h�N�~�yN4vh
+	�[�l�jn�q�wP8֗��s�E:��A</�����lcZT=�F�g�/�<�KL��͟�1׸���W�qt���o��s�I����Icg��RY}ʝ5�ɉ�/�d\m�౉�~#��b��=��s�;��G��bwE��FZϝ�*��o�����Tq���~=Ͻ�Dd�/l�k�k1�u�c����<no���1�y��]��,��N�~PzJ<��$�A7k����S�W�c-�]9�B�:��=�K<!�^���*��C������ۋwZ/iˇ�갘e#J��3�(��Ny, ��u��NH��L�K��}��Ў��s'/�GS'�*�O�p��K��A/�S3(�Xé�5����M��4";��eƽ��E�8VD.Mɏʶ4k����2?}Ɐ���Ĵ��LR�M�*��z�f�b2��Jp��VI'2����q�gP2�������@`!��	W�k/{�4�0���,z�.��s�W�e�f7Y���ƭ��T�p�Z�i��^p�r-+�L���cC�8Bc��d����	�ͷ�	�.t��Tbp���C�{Ӹ�g��16���n���[ -\'����)O�� k�h�/��������Q"���?�9~�����+G�9�8�9��@��^`񤸆@9M��~G����-�x2ߝ��ը�����X�ё#���Y�ƾ|{�#������ҍ��LH�O
�'�aW7Ե嗆���،5�~s��<t�i���0���C���ֺ
:�y�,?�<�k��+��Lh�#s��,��o�m6%�2e�
rǵsmҩ?t���j]�Ax��e��;�s��Ʉ�$26y�1S�u�q>1ML���w`�n(l"T� ���<�W�7(������r�$^0l+ �`kD��JL��@63������]�{� �[���
}ު)T�6W7�=�J�E�D`OQ}u�K��7�������J6>�Zxd`IԋI�=ӊ\� ?����~���1�'��aϐE��r���O#\�ܰ�F_���|�F`z����|,Vx�u=I��[M�W%��ա��#�����-��Y���C��\$�$S��x;ڬ����o���u��Q���Ap	fI �~�5�����A:���n����o�7_��o;��3�Y�=����+� ��1�����U:�4�H����'+�N����C�Y܈R��:j�Gm,ҝӏ�Ƽ ��X���"db�G�V~�;���13�3]�F�����>k�G����R��H���Chb,_>�uȄ_�&W�83��2�1�T6A�c��N8���J��²��T���64�/�l1ٿ��G�ǉ<�<WH�!���J��L�ZI-����Q��ş]N}}{��+\�9��#�Q�/"����4ًgbʭ;(���.FV�M�X�O�>���9�۫�@�?����gr1U�^e B�w����:�(m��/�FH��ڍ0���\�*��m`����������+���j^m7'���Pf�lU['Űْ6�f�N���.p�u��f���f?��z�>�Kl^�O��9l�Ǘ{��Du��!i�_���%���!W[��tsL�dA��x�A�d!�Jl�����H=�h3\m�,�������K�X��ԓ|�e��.ˡ--P�8p&3T��s\�4�)H�,x��z�F4{8uo��k�I-\b�zY�n�D�{[(�d�p�MKf@6�,3<U�������"m�YՓ��#��ђCG��) 0��O�����`����*���F	�Cn�]�_x,�W!6��qcy�N֖���v�U���.��8Q��s-�o^�$1Z%XY}�]�5��vR�"��#`�iI�*B?=,�s/63y�΃�WC�L=�@�v�/�2kV]`���2 �c�NvU�����`ҟA�ͺ�?�!�g�R.~��]�B*]�_OVʙֈ�M<:��J���|�@ �h� 5�Gx~���Ek��5���Bf^���<N��+�����S{@�Gn�=��5f�2��K�?9	
(�2�ZH_X���4T'�Uu�V?)��F���,Tjۿ��$������7{���"��G)��M*cX��J�s~��N�e\�۶�����&˗����)<pF�[E��F��1�$4|	[����,S��+�@
#��j�b��[V[R+��껿zv���:��!�lV����73��7��:}}�됖���Lm�9���굂��[��|Z�e,�႞QT���f���$d���I4�ˏ$W���_{{��l)B/(+Q�>�X�B�A�n|}�d�"/
#�wN�է�v��B�qH�� <�
�׋X����^�&��f'8�b��nC�ػo%@h�X�
^��~Y���x�7�n�"I,7k�
�PH�{�?!ҕ�ףʾ=�W�@Ej�"��u�L�}�e�F�s�V���Ao4���8�~�W��#E����,�XJ=v�xE� �ԺYe��l�'t1A7L����>+bQ���h&�r��W�B�Z�mG��1,����y�P ����ځ{YV�7/�<F	��H�+?�9���ݺ�F�_	���p|v6��z�����P��U����xF���܎a�	1��r�fl�!�N��)�p����4�K��_3��,��� �"Z_�jT��iq��ɒX%� ��\9e�GD���f�ǭ�6���E�"���QV�$��wA��H�£�Sd	����}�Nz'�.��f�r���=�-�1R?�����Y'�r��Xmx��G�O�S��3��C��S}an��������y6��{�*k��B*����@�L����O��!%���m�pctVx�w��s'�a_/����Jc�!��-�������p��f��>���1�6Mm7��tHV�5�+�u$%w��u�{Wk4$&�88�?9;����C�4z{(�,�3�c��n�
�c�˄)��Y���`�n|+��\��ۂ�8"�X��~:�G���Of��-��K��ЧLR�!���'�|�⃕��7~0��ǀ�wv�dC�$Wb�)�h�}���/�!��+q�m�e}}$n{N��FRvz?(}{�9�!���G���F��I\3!G]&&Bʉo�!4�,�#�^��g�T���w>���W�:U^���j?��N<����/��gJ &pƞ�V<V]*eW� ����(���o-椛����n��>�T�
���/QW0e�f~��d�=��n��h���F��4�zq����p#��fOI�B����˅Z|��p�(����}�~Ƃ�v�����5��^7��A��|�N��_o���9�Y�J�H�����Q��$�A�@oD�~��w�鍧�-�ڭz&��I=6K"
����N�!$�~�t�g��ێ���l��f_��ݓ��?��z�}�E�I���o��YV2�&8���1g"���F���X�3�]�7���rb�2/�|!!d�;�i4
c�8@w<�u�z4*�ut�����.�ݑ�}���0���s�.�a]uP�mMw��\�\wgۣ|*c���V�D�O��v���/&�]����LXV�(q��$�z���`���L��FI�sv��?��{��]��G��!��+ꊥ��T�D$i��ł1�2����a��4ɉ�K$嗿sHw�<ǾH�@�А��	bD~q���C�y+�3}|b-1�;��ZOSLhZ/6��&�<�g$�y�^(�b�G� P*�W��R���8p��#�Zc�i81q	�����2����9U��aם�v�s��8!|���^$,ny�?�$"1F�q�A5#JI�OփM�PZ�9���А��gۮ���?��t�z#HD�Y{qh���H��Z���b�\�%'>x�Y�1B�X�����,8���0�j(=7�Y��s��X	M�m�g�
"zf����X�^�G5�C5}W���g���y��D�Y�2�x���q��D䆔�;ĕ��7��6�d�?�o��ۈ"�)�Y�� 2)�����d� aڃ%��~AN�+dEu ��	�|���Z�)p#=�OZ
���k�q�:�9��LSY��g]��7?e�h�[Gqj6g~^k�tTslӎ��p����y�����
��^�W��A3�$�%����cN����>�\��I9�D�w���־��p��Z��������Ю�=��g֌cOK��S��o��/\�	{�㥇#o'2@���+nz��,|�R@�,��Mf��49H`��!��g]�/���K���u�J`k���}�W���߽T0F2�]�*�\ٿ!����ّ�)*�M�G��;(���?j�fL�n�!:X��wqLo���.jz>�1�A©3�5Vއ����C��W�h�k�䭦�x�[:��������5n-�|D[�����<c�F�ouCO�bs��}c4� Z �0-��vF=lQ{��W>���le��s��}jYO<XƋ�R`�j��J��r�{�2��'�Q�w�1z;/<�?����Z�Ǐ��ھ��������QB��K[Ϸ��HJ ��2�/����ҝ��;���,/��]-j��u-P&� V��E@)����!b�M�P�aZT�uu\:VB���+�U�˻X:����
X�mM]��ǃ<XL�}MІ5�
�݉���*��<���A�$����&F����,�a��6�O����)��ۍL�.֏x�B�M%tC��c�D�a�<ﰕ����a`dl����n[�K�4�^�m��+}���5�8�<s]�؎iSu���Y+6�\;⯨�,�Em,Q�Y�����=Qst��#}A�=�)�����W��c�W��(Yj�(��ֵw��TB}�x�*����upI�Ah��]�є
�.(� �\��g��I6�?`I	UU�'0H�^�6Y����Q�#9"�Ff;�k552����kN-q�c"fĠ��@��$Z��O?�`�ݭ[�ZL�YU�b��.�juii�dz��ez��P�N�D�>E���.v�c"y�갾��E����T�� �K��k�%�����&{r�ۤ��r0��C�^�)���r�W�����BvYv;��5��+��B�}�Jj8���_8�.~QB	7;�qA��dv��r��&c`�U8���:�^�HS&�6�5m�|��;҆#'�f�9�'*"=AGm�3p�r��*Ӽ���CF����I�dO(ۮ�S��mu�$�H$M+���э��M��])_�qD��>Q%�n��
9\/���Q����<�쒡ZstH��=s=h�t�ʉ֑��>�#-c�݉�����-\!��W�],k�K OF������&��	�)�Rֹ���˿M	��$&���Ⱦ�䋠Y�X�cz����_Ә��Y��Fd�	��C��-�R�\E_�qT�h`����F���������⪖ b�P?�s���0o���^���SJ�1"?F��FVT��
?��R�|!��S��9����Ri���F+�R]��y��͢����*�_x��d����[��"EڽH�ۺ���Q7nc��ڳbt���e{5|{�V��b���*�[C�� �k���(
~��%V�y*��EIIs��#��4ǣ?��DY�Ծ�a�)�/�fN�ѻ�{�+�̛~8_��|s�vv�xی��#Y?�S��X���y���ƙ�)���4o��Cyy뙛��i�	{ka�ቇQ�w�JFY2�L?�^]��Y��6����Q��Չ*>g�ŷ0��I��6�������S~ϖ�띗n��ͯU��O/���	'�[=@E�^�6�F��y�������޼9�����/zk|�P�=��0-<9[�h}�Of ��>䍱ieGJ�Nhy)4��s�j���L�-ȝ�߽L:	���pr�����T(Y���g�HsfO�I���ń{�x"����^U.�h���R�p����+�Q��?	�8����8d5�5Oo�y���(�r��U@�����#����a�5
�n�:���cHJ�З!�/R�G!�k�� 6��q��o�B�^0�6?����ؗ�.��Η�ˠ��S?�+yv%y��܅�z�v����_���I-���?r����U�(���v�H)5�M/�.��8&p�	� ��!��կG@��M��o�+s}�kRaGZ$EK��!�T��v�z����_�Ğ4��#v<�6���V���uqT/"nӛ�Z�:�����Q��
���pe!���.�+ ��Ỉ����t03�#C���
�58Yp��vS~h�M;U	a$��"��1�R]��6���(�4��v<�%cWQ�m��Ó��2$��h����xI{l���O�|�;�e����^o>@<��f��ە��:�jJl�����~6y�T����ǳ�Z��k��̊��%�n	�+"�����e����D���;���gb�n��C~���it�y������>��h����('��T+�SY��SS��=[WL�����~&� H�6'��[yp>}�2�$�,��1J������e���p�fz��k�`�2W�;ەʩe��w��Y���5�����-m-�Z~���x���,��Ii���O��~�(OB�:����.�AgF�i+�S�k�@����E���ׄy���&�
UVa���7TiX��m�I-@e���y���6j�}U@�YE
$o���q�AN��^���=GD�٨�~���1��B&8rjK<��{���w|�A����G�B�ԧ�����~�ʳ�AK��Ǻ�c��S4|�q(:l�N�y(�Go�F�U�s�6k���W��'f��T��TogY0Y	�!�������z�<<��O|v�����q߰3§(ļ,Ȼ9��FG�BE��s��O���sC�ε�Ι�c����f�Ǭ���Ě�j�p��k�~Q������
j��[t>��T#���N=ǭh �vRx�Z�r�����A$,��n� ]��zE��e���~���ѯ��\��J6�Oq.����rZY��6�v[w|�����O\��>Ḱ�� �
z�������g��K2Mu0w9�[`��~㭯8Ҭ�� �3h�?y�\0�@=%Z�a<�dZWYܙ�>e�kI�q�W�M~m�hY!H١z槡������k0Ti���n͉՟��c��(�fG����������jO�v��g�B�5�<|��?D����g��ﳕ��P�\d���y_*؉LC_he�	9�HH=��K>�G�s�@!V&u >L4�}��.`����x��K��B�(J%r���c�7��m�R~	|�<l^k�e�l�a$��1�����h^O�zF3����d��e>AF� ��:ų�B��m����kx�+��mԊ�3��}��\�ο�� c[\H�mm��,E�]��e���/�Z�q�"�ѝ��Ol)���_���U��v1�6G�d����h�������8�������v��D�h��hF��R�v���y=8,�������O�6�L�"�Z�!6����l,�Q%7l��)ނ}E:���0��4l��g�r����*�'&�����C?~0�Q��y�y��}R���ӣ���e-�lg�z�6�[��\���OP%�Z*,w���e�1n�����ކ#�$(� �X2'F�LB[c�ݳF��b�~�5���O�9��m�x��_H2��v_l�H��5_��&���0"����ӝ�ņڠe`=~`��������@Y���?D] ��%� j�
�e��I�_o�X�ے_�\ҼD�-�?��}�0�U%8�E�b5ds`0~U�ӱ�I6[D����&���V�f�c?���!/ ���nx����6�U~߬���GV��o�%�ے,j<�Ӷ��o��Z��6���R�����Q���O;��T��nP��{\�!�Y?�a�O�gD	c�
��@G�rd�8��|2�\�����2�y�kh���cٖg��CnS+q{��tCB� �D��aץ���N���R��xA2?��㰽�(�ݫ�'�N����SA׻pO �t���Ip���C�9!�����W�����%�}��zoߘ�'x�8�w�Pf�#���o�=��+�goy	�/|o<$A�i�I�;r��&+EA ���Һ*hY�E��~GH|����,�!)-I���O�gc}c`Pa������D��5��0���ad�[���������'�u� ����:z�N��a(��<��򺄳� c�a�-g�ן|�U4��铓�z|87��m��_f��ﻏ`
.j����Q�� ����b�8R8������%䆇���/*�Ea�Jxȧd���NYOq.�
�?;n{���L^�8H�Q�Z��B��#�U=����@���A]a��z��)�������'aV�b,dP_�{bX����F���4xcUD)Ѵ�y�3y���僈����k�&��G]���M�K�#r4�-pN&8q�V�V���R!C�m&��4P���ҹ oƱ��+d�W�`;���������I��|)�)��1�O�u��JA��"���T�{@�qVؑ�[Z� y��%����F#�c�T���U_7��ŷ|�J�����N�J=��������Λ��Q�r�7g����F��h� (�:�ڃwd�1��0��>�ѽۼ���yc�$�"l��i��]rן������Bp�CQ�G��@��ߣ(?�m}Lu�+�?D�M���)��h_���	&+�T_�u���m7ժ&/����TROk8˟^(^�h9��h�߁D@^�/a`�a	��w5�خ�f��\�F�F�,�YR�le�x��y����d�gR�h���^6T�tt^=f^]|ɖ�|��x���]���HuP���\�}�`�i�"dz�����"h��짼g4mR�u���n���Y��Y�~��z-=0��.XXʐ�TJ)��s��J�r����z���.Z-g�\�h:�Ɣ����}9:k�<���p������C���W����?7?Mw���+�ڳk_j���9=���*D[��E,�j�����K6�`��BQ��%��*��E{j/�p����a��4L=,���,��I����5(�����1HYi B '~��~V�7�J�=��q��粘�	tL�u!4�4��}��}r�<,.�K
?��gvx� p����e8>�b�*=e��\?Iݾ�t���䫎���I
QP����d	)��Y�m��7���ٽ��>p�Ip�7���|�)ŷ89�w?:��� K���O��?,��5�+�	���Kb/`�Vx�x�M%�:n��i�)��Y�d�,e�i.��E�,'\��um���a������P0�L]�g�I���GY�M{�7/bGL�Zt��k��?��s�@t�
� !��l�īiZ���O�'���i0�)q?�My�O�Ra�P_zN��+3�����6R�H�ay�I �ꁿ�VV��{_Nk�6&^ϊ/N���٤dD�6҄B6�+k�c!�j���Nf;ƬlGjL}�-���O��Ӈ�%v<F����ԈMG�e���/y�%C���YH���먝�,�o�Yˉ��+@G�[�k>��N�����J?�κ�*8�|�m��I���jK��-�x��d�T��y��׽���Xǁ2�ę��8ѳ�Ӱ�<�M*Û�0��6Q!b��Z�/1ၻY�2���k�hA������M� ��Oo��Ih%�r��ܳD����Cc:��*g���2�+���U�
����A��L�3�:*Q6���o�2F�c���8%7�i��i��=yo�񪦶�S>�U����㓸����,�L��n7׳�뮊�$��o �p
��W��g�sT��7�D���$���;n\�9����Gx�q�6�G��հ�(I���&�:��!;iφ�a�Mz6{fS`k���_D��ۙ����F��6ͫ�-���7��Œ)7
S�����~N�vMk��N�7�8o��v���\;�d���m�^��K��,|��%�j[��X4H#W�����-1�UE �=�Z������w�E�N�jڶ�����ʇ����t�9}��;۟�xm�c�H�'-lm�8�;Ah�?Jr���1��n0GDcx�����2��6�rJR�02w����� �A���j�#= .sbY^��i2�Q�/���\���y5v��}�����\��W�YT]��[�󨐏�v���4��U��d3���5��g��B����b������>��2H�;�A6�����i���h�m�<NE�z	����Q���/���Y�!��Q��
����|��ob=�ͬZ�=W˺T,Px%"�%�rV@����'B.}3�O3]y��!��߸@s ���Tvנ���浛瓻64�����L���%:~��!ç}���l�esۖ��HP��m.�����Gnx*�y�Rq�h�7�v��D�����,EY�z��B����g��m��C��_άxS_*��Km� �4�����A��kxH-�i��~[�������S"�t�����dW���4���o�|F�ho�"�[W��v4J��y����?e:�5)`?�gz]��6lY�5{�-�甁9���h�m"pܽ����ثT��̹�^�z�N:;��I��5�FG�\}O��L/����eU�#>8��4�6�m�$p��eh�j-�-�^]��i���$c�m�(�i*
����M.}|y Ǔ�b���xoX�+���������� �w�5�|=?h��,���5N1ÒS���r�A�~}{���N�����E��o�K��d�^�&��ױz]�
���v���V|���q����T��ӇG���Z��xAO�rN�Z(�"T��ʲa��
:�o;�8��`Y�,H�EY�%W{!N�����N�^����ù��cu|L�k��B��MΪ]?@����*�l�X^��"��;�$�ׅH���	����;�E∦���ݹ�#ZD�d �>)&���d~G��E_�D�]d���~���>�|�����p �ku��i��
�N �b�E%>͸2��*�y�2%������2 �6����@Ȓ��\Ճ[�f�1��4�h��u�v�����202yU�����M�1��������D~Q�Yts/��`�~��&�κ�U���FyS�ֳ����J@}c���+|sU@���@�lq-�(�h�^�Lֵ�u�l3�c�d�h)a����59��2��jGk�{��:��Ml³aǷa�C��n`G���ƽ�҂����c�20�a�_�}��m[��ٲ;�5�+�x��/���xZ
*�p`�}<� �5�ɫp@!�j2_Ɔ��rl|E�<s��lP�S|��K��qv��&�̆*�@��G�Pp�R3�>��F�t����e!�cN�[T�f?&�����&�:�/�V%��Y���.ޞ |��c�q��z��c��7}D�E�� �x���������at��7��G��E��� VBt�����8<�K�)�+͈��ڼz�-�q��4���ϋ_W�>������"�n�'{:�ŵ?��C����K�	9��!J� 2��̍ft�b����tݖ\�XN�y��o.� �x�k��0�A���?��vst�|��W�\T��Fk�m���p}.K� )���%���?�yGW�8��A�W|� 2gTH��5N��'�ej��{��W	=����^w��	Y���R���m�5x��������I������RtW�<x�JP�h�9��J��_�82��ʀ5�+9��n���G\u	�z���P���=i;j���y�U	=	2���J�aғ���㪌;6^I�r��l��Ͱ����"Y�wk"��KΕ�����y����oL�&�9�W1�6iY�t���1���UL�C-�ZO�U8Wo? �����NjǏ%����w���=MRaQET�v��X~vp&*#����K��m<�|�,o�|曈�=�Gvs��/�e����NQn�uCN��6)�� ],�V=��JS ��_?*@}+����5��A��t�/��Ng���NҬU	BFM]a3���87�,N��@�Ձ��q���zvU�v88�2;w@k\R�䱻ɛʻ8�^u*����؞Qi��j�%��N�:Y6Ǻ�]�u
��*�~
�we��(�'*fM.Zj��?t���$BK��,��������`�F���NK�{Ւ�_bo�#�QqNҞ;	m����б� C�CxRd;ƽS��еK8iN��߄�D�R��3NX.��������El��}Ԇ_`F=I�>JX�������^&w%s�KiS��t�f��O�T���ѵ�zX���3���ե�I��g
�ſ~��ȏ��D/c�G��J�29�)H_����L�xP����!��H>PG�����<c�f��+��Ӷ|�*��H?���Tx*�	�~�C���v��p��N��,����.w<�t�O���м������MƠ�*��dz����ޣu�s�n�s�=d��%���.��F:zbV��%/e��$F�*�hZ\i{_Fv�����M8Gِ���*�~T�ZrW�L�n���R��Yʛ��}kW�n�̡�檴g�&�S��T�꽙�#��Z�����v�b�G<����|�}�j���u.Sis��=�^��8?O!�)�Y�6���H��U,��u�l�TK���#8']$e�������\���>��{��w��5��jB>%S#^��(B���.}2H�=TO�K@%b�����|]J�?V�	X�8�l����*�7s-�3��	&��(�) �|�_c�1qC�@�Z���wgU���U��+S�E紡*�h�8R��EG�5q�"'S/�'��h%.V�~ �v��.��J�	�7,@��~�=���3O��B��SY#�	����)Csf����!�Q|1V_|��cT��b�����2���■�e�c#�Y
����͕~��F[�	�,aM���Y3G��FD�D��{5�m:���yA�M����sn�|���$x� ٔ@U���d���M�vky�"�"�^AyFM���`���ث��%q�����c˥�r��G�:��r��L�����k/��͓��p��71�(�K�uB��wπ��ޫA����\/mʲ�Z�r���T���"�r��U6F����醲<R�>F���!�^�s�}��d?�l�d.ل��\"�x�mcn��%��	IH��F��JЅ�#��8��`���� �47����7g����j+ %լ{�=�m+B�;����8s�iK�H*fJ���Qw
��֗�'!���������AF4 g�����q@)�]����6?4t�
��m&��!re�d��=�q�
�ӹ����9ׂ�z���d6Bt�����*�	�~)|��Ř(,�l�m�uX��dJ�O�ӹ5 >�d@\�7b����e{� (���7?��.�'&{;i�����v��Ӕ��A�� 5n��KuY�'�M�	��}�z��9�:��$�I�`nv�?��T/��Ĭ:�v�i3�0��/��Q:_9�'����.���\�3����>���r>P4���������ƶ���n��ڎ��I�
�e�֟�A)�n2*��T�Ӥ�4�b�f�P���(�5A�%K��i�@��DS�6��yZ\�-,�V��"�T�9�&�ڃ%���v��i�?���fl��ш�0O�!�_łۉ��C�f�J��N��xVyrѸw�+�_KsA���7����y�4��2�\ꢾ"$d��k��2��+uZ�3D,���U�lB�ESJ��B��#)��U���#��Ŏ��O�
���4�p�ݡ}�_:�� ?pV�\�W:bڦ�4.	߆H��t��UJ�'G!��7��O��Oۇk�$��ϢO�8�d֬�<���"(������ы���s��I��Rsaݸ��0�r����o��M����MTڗ��zߠYնx|&襤o}$��m7ŕPRw�J<��E�98Lo������b��B�8��?@�?�5�3���lԽ>�*�� �>�W���g 0��Jć�"~lM��[�'��L���@�;D�<�������D���?�.��a!�g����u���5+h/zw)���_���ֳK�~�_�o���o�Y���ұ��9�:%u�`�ikuH=ӧ�Ŝ��#-��٠�A��������ŎZ�Z��Y�!��_htz��K�~�y��w^�*��LB��d�#���������o��J�c'T��^p-�g��ݰ��J��<����p�ǔk�x-������|4w���>��E��H|>s#[=;U�M���6s�=@������f���R׶T�|��Y/���.��Bw\��*ʁ��1�j����o��4ۛp�<c�t ��gx�{����"��eOU4g<,�`[�T��U*�:�pS��D�ڽ�y�yu��E��[�WWo����R�� #����k���t�_�?���P��X��LWX�����m/��c�l��h�>C���k��B �Z�X^N��N������]wP�!	}h��N��8{�����P����$Y	�U����+�J�D"~�U���Ի�v�\�z��6�ߺm�z"4c9��5��v%���`��~D;��@NX�3�d�:�t���!���V�^��y`x�=�f'Z����'wk�d�h���d�|����sY���zw�Žn�t>��)��FW��٥���ͽ�u�]�
&���f�S���{\z���8�qג�=&��ƶb�[���3���b/��6�|�i'V�լϝ)��p�NR.���Dį��S�._v�2W�u[����ʵ�(���8H<��	;]�����Z������C���!L���p�ᦕ�v�#>�����q�,�_���s:�Ux���2.ј��[����4t����̛��:��t��4�����������ۣw�����$ő�,�;�D�sOw]=�2ߴX�	�;��0��[-:����X��.���\g_ǩK�F���r�넣̪Z��t/�&>Swt+b��������y��T��ژ��zL��S���ΔM�+w;��+��]���>'h7�yN�0Ъ�#r���O������8]Z��zr������Mva�`��`ҡ" �R�%D@�A�k�6a��` S����" ���ݰ!�Q��>��>�|�O�s�s����9g"V
�LJ��O+��
��f���Tخ�PЎr��U�Z��E�#�0 Ʒ*�m���Q	^3�4��n�=�c����85����QM���)Q�lE6�6��B��Ş�˿%�lPx�b&��g��M�@���/j�Q��Ǒs�L=�{K[*�X;UU�'��"0�^���L}ܻ� ������Y H�!ӤL�o{���OşU�>���r�p����ֺ�P����{�В�w�x�{����
����b-7{���_434�#�U�s�1*32���.%h'�$E2�:��P�zn�Zm[Ps?����^�b��:+V���"���2a:(�����Ϣ+~o�J%�����6V�E;�詫�J�W�4�L�N�7G[yWi��*FW�F.}x%��\�LRG����O�ՙ�J��|���[C!�qS�Z&�q����`�K�j����>�0��/���t�KC#�H�=C��D�Y�A��L��ت����=��C_�w�2҄�F|������o?�9��#�@'LWwc���b3�c�����x�q�c�P�P�g�}��(���6���m�T�4?�ߚ��}���"g00���S�M�hR��%diЅs%)��x��%�)4��L~t��dy+��CIr);U�Q��Jp}B�绿�rKy�'��@(��i���}F�_�0H�m��TN)f̺	/�=AS U��X:c]u����0t�,;�p4�f�����m$͵�G��OmKJ;z,�R�/
��2f��A�>,q�-͟��a�5�s����x��cVw�xC}3�O:6 י�뚆c���0�����4�u��<|\?�G�1g��(/�0/3,S��KS�i
�z�P�&��5���Ĳnu^G9)�(ֲk�D���]���5�Xz��Z�zMn�p�uX��h_��$H�(�_��C���L�PliL<�!����Y�u���Ih�R��(e�f���#��NbF���큕�8���?���V���� ߳K��=2*6�96��!� �ʴ��|PV)ڤ�j�]���F%Pj��O����1hv�$�~̄�ë=�\���~���#a����G��KLz(l_��|��޸q�[Fe�����"vg��Lfc�=��\`��8��>��<�&��],�aN54��������t��H%�q]��B�B,��PY�@ �ni�F���0_�`���&Ŭ���b���0��R�iB��P�t��k`�<��Wc4&�ϧT,��Lhn��>�2�cϾi{�踣�����!S���ȴ�[���V��S��O�A���A�$�ZY�5�Y���I���~T��8�(�k��c��S�r�1��4����Ҥ$��Ӹ=z�8����ӪȓH��1��7t�Ŷ��5bt,�E�1ǒZ��W������o\��d�k�:������{�{!�|K�T���@Z*����(���>�v/�0�//����5Ja�rj.�M��	w>L~���q_��4p���E�>/E�[�e��v��&����L��=��bEϑMj���a��nt���>�H���L��?�B$XQ�r�霝����(Q�TK��f�C�ki/#�����J��~�w�_�b�*2�.ױ���(h�m����5��G/9�����)`/R<ϸ-���������k��h��f�Ŝ�<�،4���d��h7���α��]��02L
V�]��_����>��:'?���]&���Tw7\���$͙0���>:h�w[����lxl��S�Q��QT����@1��]����R�=P����T�j'o�Q��#�H�i#��l~�t��N�5az���ysBQŉ��v��{݉6�x2���|@��s�?�va��<o�e^\�'q��Pa��B���x^���Y�H˧��E�2���!�7���+z�iF՝���q�TS��`��j�4�P�N)�Г�q|����G�^1&��4o9 ŪD7	VI_ˎllQ�Dߝ|��,����o��M� ��u�EJ=�r��&V������<�: ��dy��<�tS��/5j*���we�덛��#�&��uHч>�N�_��X<�^�˕t��Hr	��F��f�5d.\S��;l����~����y��v�.Y;�t�]�g�Q֥\4�v��EF~�ޯB��:|�3\~�_�50s|�UWùW!]y7�T	�Y/���Z�(��jW)`y�J4%�Rh!���v���������ܸ��6pC�"�����ۛ��'g5P�Qy܋oإ�nvm�_�V�uU�d�TUn���(^t�6$_����f��V�Z�&,��9K+��Z��+��,WJ�i"v�e����w������(��>0�f�h���?{�G%�}�"�{�I��5�ܧ��~��U`�,��TU���FNA��S�����n�a6}�\�T�=�S�]h<�3ϡ��(m)�tV���K���( sVb��:˦[Qס�kv��'$�jq�籱X�6�V�r�Mk��I��� �3~���t�A6Hssg���ػ��� {2���咴��r��v��j�'�@��<>��4Y��y;����6��~��̠7-�1�M�xi��tz�.�iVw#ȼl���I�ZZ�̸ӱ�5���@p��i^��E�9E�ި�o�'��M;�_Pm��l��'~�����ʿ1Pu)f��ݾGӛE��;Z�U#�Q��E<]` B��V'��m�"^DR8
ܿB����rm1�$�^>z����k�^����#?�kW�����}SR{�UצoO>Mc���ʆ�K���Ҧ= ��`-�K���M�S� Ƣ¦�_P�Vg��o���Th���:�Ή"=6���pv�9�������]8Qq�`�>���P�_�	u��6�G<������b%��(���f�y%��s��JXE���� ��͠D40'���ѵ�c�M5'(�m����)h����:�c���}H�3I5�e�	!�X�{4�]t���/n/?�)�4g c���S�2���1 #KF��;=d���2s�[��2��&�a{�x |+MSH,�-��܂5��W݋=�&E�]�:�;���2|��t0��e�"~]�k,�A�o���!]�^ �=�2Y���͝=0v��d���x�'�l7�2k��B��*e�"��5����ڱg|��$��y����=��y1t� �ӧ������ű�ĩ}��nEr�*��.�yg�O�]������v�� �}�@�3}������yvmI�������۠F��p]�*��c7�D���<P�0M��������@a�����[�:�<��xX�U��y��+�Ҟ4����=��e7�S`�L��ݨH��1\��;WC�� g��e�n�[J�_q��;
�@WĶ�m�.1��V4�''ιV�P�<�����[(<�'�Q���$-��8�Vk�S���Y:	�5��9������J#�R��R�&͠6!�U���#�H���}b?ϊѦ��zNQ)� J�Bk?%���pr�����Hu�/F��������E#9��j�48�z5nikpg�.�ȴ��_5'/���1~��]���W��|���6�ͼ{<{���P�@n�����Sg��-ç�&�h�3���tN!�[fu~Л�yK����M�"O%�a��~���5�ľ/7�����'������V�'H�emtR�jA ��[�v)��E~>aџ=H�\�[����|p��1>�����u0�t�]5�
�N�z��jr����+b��:s���&�eK��}�&=����z���e�lJ���Fke���b�V��&���
"��6�@j��%�u=�U��X��(�9����?��O���rh�?���O��=��F7k��V|��eE��ˉ�E�	<i*�P'���;g�?2C��>�122&h��[��������`���>Ҳ�Q�
mg@�e��~w��E��Cw��"�����zh2<ג>��&1s���9��}��=Z�p���NցO�[X���+z�ߓ;�'@@�O =�(���ӎ>�/�t���5�J2�|5�L�Yꗨ�3h�-��<!^��0�숡�d�{�sv�z����GEV����+�̰�?��t����6,������/Ts��=}+9U�5��a��眆���	v�I����ِ<ǂ��yNNW/^<aL9hu�k{����=M���O�A6w7<�L��c#ffn����g�۠�?�dBG	���}��	}Hs)<��Chh�ϔ���ͬ���Y��������O{�\�����||��׍�y�����e2�m����D�߸���߸�>s�q�����q�Y�c��/&F��iZ���o�4M���B�2�<;��w׽,�Hi�8�M�z�r�r��j������W��@@5��^�wo	aQ�f�6�F-V��z\��$ׂ�4�_uS�9����oT0��7�5���֮Io[��#�v��_C;����L�!0�k��?��F�^�^�LY��ǡtS�+�j��JE\`�r�s�ȭ��	p�-tր�hq��6���8/��QDRt��]*_���*E������z��{[Jk��9u���y�k�O�%c[i��7P]Q��T���Ly����[�����T��Ȃ�AB�R��n���F.�4x��u�[�oU�ǟy�|&[������O6�~vk7�La�V���,�?G�!N(���s�-�	[w��'�L������Ꙅ���X���,~�f�I4D�%?()x<6����Q���>8���Bf��ho<��݌�U�u�O�����ؗVY�=O��_�9��ӀN���C��_�2)��̬S����u���%Y~������h�h*����M+�\��Kg�Q��͝�=������\������� �G�-R�c/��r\�6'�v��ð<�!Z�~��o�:?粳��U�YHa�aC7��gէ�Ƽ[�����M�1�����CF�O��W쬰uEw*{e�!&HI*���j��t�\����h��EY�����͒��Pr�uS�� E��uY��!�۶	��Y팣*��PD���;`U�1�� ���E����9�N���VA9\	لQU���6w�柩�%5�w��r�P�=�P��lX7W�p8G���F���J	���=�2G�F�O�_�/�n�]��Z5-�*�I�3R���r����Ć26���綍�n6�B3�v�t����؆����՗alBޫ\���u\���0uݴp�.6��a�왠�?jAd0�^��-|\�G�76����n:����� ��ڊKws jyJ�|�x/�9�s*��ԣ�Lq���I�$�ph�-O�H�Ņ�O�(7���K�Wؚ*�k�D�a�@��������K����ذa*V�,x��^1�i��hǖ���x������u�&
E\\?�u��z�-ly���K��B�[~����Ty�)	>쪞�v��sr���n�W"j.��R$��7B�Mɇ���I��+���Q��'�Z���+1�̵��'�r��Kͮ]��>ɂ,Qyf�>Ycc�7�:�9�=�������/T.j�E��>M�t��>o�#hs�М��A�����N��a;�x\�硺+��DG�-	d7��+Q���iA��ß�����}�&|�0RG-�ٮ�_������(���Irݏ�X��Nűq��kS��h\��],�e����?�ݚ9�O��Z�>����k<�}�o$�U�,r�g�Gu�w�w�,���Er�P�i���Be�p�2!�U?b_@�ӝg���E�g���6_���w��"�ȳ�a�4?��w�ij��9ff2�\�T :/��5�OJ�_�=;��i��HL��JUQ�Pj4�C�L�jc���a�h3���˟��IoyKX�'��VG.ض����E���Gkn_���1c,y�H0��ۻ��.sϑ�@q������v�'�-����&"�z�nZ[=��]��^h�]�������7e!.��א`���O���{
��o�5��#r��0*�r%�h!b�˓C�V�p��I�����G^�=����O�����<�yy|kF�g��I٣��q��&?�
��������k�<����}8��x��Q��y����Cz|��5o!�b,�^��#~��Ͳ��M��l��7��6�,��B���z�诮(.|��`���(�u]�"�2oXtY@g�vNQS�@�(|&tO[��.fp���4���YP�T�D���1�w��_��Ӡ�(��N
);/	��@q7-qw���f�ٔ@�� G�k��L���K_M��}3O3��W?�;&?J9 !�p��^�*�+bJ�kF
L$^b/���R*w@��C��q�َ�3�/��Y%�)mw.B	<���l�R|�}��T�SܷH��p`$e�V\C]�S&���;���W?��V9IgG!t�[%�ڗ�����L	`sA \��du5���U� ���f��Nꪠ��P0Ҡ���(d�VCCe��T6%��I2��p�ws2-Z�5�vt�KW!�F��P�oJ��1�ܓ�<n"Pjy�[�5PD�������?qg�Kr!���cOCV��Z#}7v�yy��%u{�uu��u�%���`>�y�fy��g>Z]���H���z�6�LCw�̶��ڇs�J^�W��~��kol��;�^4��.^T)#⼗�����V�͜�`�A־�J@��I��Q�N-�*H��M-�������˻����GV�Mj�!����+d*�Ɣ޻7YV&$��"�ԍ��f*��3��#�������O}�E2�P��;UL���+͠�2	��R��}Mͮ��C[\�t��_N���wg��ʂ��'E���]b��y۠ݻ=k.8�d)f��
v���=V�Q�団��
�{�VĿ�R�����j��l��҇�W�L�qhYfJ��j��[^TU-O���E�����i��>�?6zy�+�EjAB�F;cD�|���>�-t���E���U?+[*~?ĵJ�׉��Ď�{���	��'Q�2���𦠋Q�o��b�[�[ҕRRE����t�+Ԏ��_���tP;I����\/Cx���I��D�A�{RI[i���ZΩQ�#����C�_�y��{�𤸻<<b�q1I?Em�u�g�/G��6�-$ڹ�Ip̸6ڿ/���µA/�y�R%8^��	�~�_4U&
zzB�6��jK	�Y��ܼ���܌�%�]+�(ܠ����
�_׀).~��Xj������MeE^�X�a���k��R�&�2����	�E�^��ic0��]��ܐ�:�tԂ�a����l&Y�-��j�O��
�އW^r4�?���9x�C�F�41'���a���f���&1'�$A�A(p.}�c�|�{�'�b��!%߄�s2M����b�UK���
��1�<;�q�$����庼%����V����/d!Κ��+m:�݅�VG�`��it�+�'���I��2��>ZA\R̋���pSf"����Ŧ/�ݪ�`�8�C>�kfG'�|��De.��N Uf�~���Ϧ%��E���w���%��I���E��z����	��:8�f��7P<b1��_�\����G -������0K���!<[,^R��������x,������Vؑ�l����O�P��z�=���r�=��K
*����k�P�Yk��� ��D_8���Q��e�[�^}�"w��NyY����VY!�al��!>^��~�$֕*pSWy�a߷2^m���͆����_��]��������mY�
��2���y������f����{3Q��kDu��|��P�ŬW��pJb��(p�535f�W�N��F��
�huY(�E��j!�y>�P�a�m�P�����XC)럏�b�Ot1�����6)[��t�ߌ���#�`�YD+�lX˭ުm�KX�IB��2,ܩ<�X����ľ`Q�r�T���2�z��83;��CU>���x6�;�=�6�V^����v��,�� �A7�r�<���F#�.��o3���E�H�J�so׻Ū(C����^�3�;BƋOu���S�{L�Q���A!����
�Fl.��_��N���C��L|_UV[��\���̒]���{o/V��!`�9��{&;�i#����������,�p3y<H7�r�
+���m*sf�)$Z� 3Z�k|�g�dR��U$ݽ,P�\��8?��%\���N`+FV&/����S�3�=٤�{���:�q�n���W�nssa��f�{����̿����N�zog�3"C��d���9��n��g|�?���&�'�W�Vg���OΉ�&���raQGb�
2~�Z�Z��2Q�Y5
�,38X���D��c#8�mI�I;-�t&�jO��SU�}7C��}�W�_��J�;�����=+'�g���oLџ��ڟ��Ć��u��=����R�z���T!���o#�P�>�.�K�}@`Ek���~<�R۹����d�H���ޜ^;��=�;NF7;X��ooil�I &�
A�:���[��0�i7çqC�*\N;�I�l��F�۸�������4�xm�8}�=;n��tU�H��F���P��K��$���w]�זe����V�)�&q�,S���<�0g��v�k��#����#�[�ox	�̗��O��h�gc�L�n� =JT)3��`N�n`e�?�0�C�J���1<lG	����4A��L�3_� z�UCk|�mf��F�C��Adߗ�l�nK�Z{��b+�ϛ���W�b�kK����Jv�mR:��z��,0?��D6e��ec*ٖ�z*��4��������]������?W�q�H�c��I�(�S��<&ç��U�$tG��}m��țP׿������H�/�j��x��#��?�C<��OŖ=+k�Z��dm�ur0�w���袋-�4]��s ��V�1B@�Y���3%��+�6>ab�j�U&jm�������i=S�&!0��,Z^�8ڡ2?����Ć0���l���'~"m|��L��0�������vu�c!N���V~��aƚ�����;�'�=�6�X�"���n�U���ŇEݣ�zx��F_��4��^��];W���l�'�ZP4�KPK�;�ay�="���#�G&�M�]�QƩ���A���2EF�!��>���md;�][�w��{�38�s]Eή��`���`�g�� �.�6ɯf$��*À�2����F5b��0:x�u�N#ㆉ�:�nmҪ3\�BD�1uq�#������W�s�j��꠪[[���q�K}yQ���$��.��X���i����k\��TO*����,������0mm}՞�>�o���J�2�ފ~KaҪ0ߚ4����!�&��"Mж+#�6b}(0�VTr^��F�)ix��E�]��˺��-)*��8��8�˦�辽f��V����F���
ޟ5�	���#4innn�o�g�6���Bܫ5�64�]����?mG$������~�!D�cm�9��N�9)�G�D�l�8�>�\���Oe�wԢ4�^__OS���$aIE�4�>����W�[����D��k��'�Ũ��o͙�Gw�>TTth����񫽟�nRL)��%����o�A�O������ƱQ]�w��k�>���`ؖ2ò�O����Oi��=�On$��������cפ�w��N��{���w��ҐHI��B��Ox� ޹u$�W�16컙�ޚ�ܻ\���؛i�.?R��z7�/O����w�ɾ�˗[��#��4�6��nƛg���R�.W�Z9	"�.�oW�.)�.~�~����U��ӧ���dk�Dg��>�˞-v�&"�\�of��{�YW�a_Ae��4I]��	�H�L|��"⮷\��LK++��jϥ����Kɣ�ie�������v���ĠCU'_��Ș�������n.�9�莢 _�W~B�\�5�rw�2��{y��}����������حsGx�^W;9��R�b�D�r��A_]h���Q_����#Z6i�:Z�>��xh�s�r��Σ�a�
U��?{�L6/�P������:���g�M��E��g��D)�~��{]"V�NK��Z�Nk�7[�9���:�F1�cLݴ~�1`������ȚC�]����gP+��+�>S�c�(.��l��x�&��zƮ'a�����@� ���U�d�]VBf��Mˬ� ��F0�5%�P��?�X��f���I(�p���r�R���'k�%ؕ�!�I��W�@w�,"��ќ�����w%Q�w��[9	'TW��S���!�l -�M�k�[BАc73��ٟ/�Wҧ�w���~`����&j��Җ$��"�(l�}��<�MNNΜ��_l:� '�!K��#L
�۹f�a�5���|�;W��
<���6s��(�sV����̭	��RM���>�q�����E^iC�hc�X�BbK�y�ht��j����X�����Ə�<����R�a'�bY�9�*++�(�`���]�n�ЙE�:����Z�i�g�N8A������X1b�=�zF�YF2b�h��u9A�?�2'<��e�&�!��ܟ��	UZP���� .x0�@���o�4����2�2�߄�b��#��ll ��{���(E�$��'<>ޑ���2; Tȟ���CX��9�N&Z0�yoŠ���XH���|�Bs6f;�'2?��3B�}�S��3�z��ti�&Bܤ���:�WA3�C����	��SB�̾\��S)��l�ȋ_Ϭ�N�~P�6`곥SCd�}xd�0�F�p����וqC6_O�OSD�jj������Hx*�3v�	��/o*��:X�-���z ��}��č  X����5�iuA�2��Hn�Y�Yz Rm�G#k��U�5cSY����rV�98�s;��q����&W�lP��R��̪*L�@���T+l'?�����������,�Ħ+CKZl����!K�J�M�bU<S�^�$��V^�)���
�y�`;�0G����,v� (��ԏw�CB����M�}w�|v��OVJ?9�"V%{��ֶ3�V:�C1H�d�̟��lbG�|+��۵��ʾL��=mݽT�nRή�W�O��6�>�N�!<!�VTՇ�F4��|��x{��7~v��b��Aׇ�R}���Yh�mV�������r���C�R��m�Bd����4 N�2��t����,�&�BB�*]�7��U2"�xmv)BzT�s���������k툷����=5L����e�O�*||����A���ߛ�ɗYhx��ޗ�^��9Y���er� ��0QW�m�F��fAl�!��uε�1��.q�	��� @�д,1��)�d�\1uւ���Aj��N��Y��6"\?�PbV��}���gdޙ�࣒��}��BY�
��Y�M ���*� XD�oq � r���H	b�R*//'��iِ��®�^*w�>��*W�J[��X���,����ͻ')����&���5�r��h��{�����Űe6�Y;J7Y=�������@W��CF��&�c�zzY��ҧ�+��� TkKd�U����u��~r`�)���������:����Wc�w�(KGA��N]�[��������uP_sX�}��NW��_�=����x�ҕ��_�߹D:�������ׯoT:ff��[ooSѲ���F3X��@r^(&�y���G���a._�'�\�r͒������lCCC��.Z��B���W���C�/ �+Z��k�y�,_�/ �Ĉ>V�:g�W�k|l8(���4�s���`���i�V�]��cDl�x�?���n��A�����з�C�|}J���ˀ��d�"""��3��<�t,}�A��H<�,�J|1uƳfE�̈́��߭<����GN�aű6֭Gv�v]����_����T��qtBH�$�}���=)��`�x\-L�����^�8�e�S�C��w�9�����-�����㟼����L�v��x��� A�0>|�Ȳ�c5�r���ƕO�H�(S��o��6�u�f^�!}ma����F��й�s��{8����Kc'k��6w|N���7+��s�Fv���p[����,����e/~� ^�qՐ���:'7H��o�F��$	U:0��C[f2�9{�(�8W����������w)6)ң��8J� ǕWZ�6�ݓ�����#��z���˫�U���^rYMd�˪�.Ğ~l!��5C����g(̄��������=(iN���O�L��t���}��:(C]�����͛�D-2���\��vw��'�Ֆ�EH��d�� ڙ�͜Q@V~��T�����!O��z �F-.2�&����lz��!%�����;�bx�Eߋ�B��o-��F?����.��ս�j��M��~dYU��u�>�
V��ɻ-xr(o�c6��؅���y���Kgr���~�0��{�~Q��d�y��zFa㪕����N^�A�A������0N����^�	��y��A���4l���x����~���PuN`sm��Eg���V}!��#@�}AcE��*����u�����'�����\_� �߷�N��af�Ršдư�v77C�b7�_��;�c��<<<�����ǩ�<��	�u�o�a �]ղ����#��g#�6���/r��TEe��v���>~r������?�%
`aV�]Lgx\����sp��2���p�@�O?"�B�u*ԍ��(nN����R�B��y��s�zQ�ϝ��;�M����DQ�����$=���9�����R��V�/�̲�����CyzE�ϟ�Z�F����;`��u�5 #��N���V�2����j�t�O7���[ic0�Є.�#K|�[K�n��;,s�&����J�[4��6F&�����V�4x��V@�3��D`E�t>]���9Z �5���]C����~]��^�̻	e��-,/�!����7<�T5��1�q�C��Pw�\��$�hJ{CM�+�6�#f�G��H�~H�] P�-|[���.R�M=<ʀi�H�+�}v75������O6 ����Un�����p[�Rd'�>�$k�h��hL�n̰9���;F1Ӟ{/F��7��sdj���#�O\G�y����Z-7ww�B������H����g�^�/��kĽcqa0�����R�ߌE���d@!�{�.���esss�T�Q�����-MMm}����*{�%��<��bb�)h�[w�U�߆�� -�~Rz4~}y|���ੰu�G��.6i~n��۫�nh*eC�Ӟi�L�(f�{y�(?�	q�!M��RYV���A^�͚�͏�'֏U�ͯ�2������&��	�r��v��|4�>��x���%]�&G;�_�lM<��H�ሸ�=v�ϟ?[x2�\�Zdeo��0޻_:���d����e`9���h��y&%ؘ�<����,�'hbع��g�@B �[Z4��'�ؖ���~c�a�p� �_}Cq!!�7o�,����7�fgg���ϵ'�CX�õ;T��z�<Y=E�u�f�x������9�v�w$�eh��k�!��mݻG��kS+rǒ��:���8RJ���Ä�����5�ի��6~�WԢ��EVM����z�Jvv��M����t����:z&Vv���:��J��t�p�>�Ѭu7��v�H�G$����^m�2�� Zd�w�?��r�_��( ���1��e�ei�kk�G��Ⱦ�ۃ�V�u��{���5�ГgΜ�= ���̥?D��ݕ���%C�Q���"���HoH�#z����9Z����**~�Z�1����!���� 
���4��l��SF��W��퉱9�	�Ǣ6�����{qE�>~��(���[W�#�afF��]nE����KyE���PGDF�O·0
+�ϵ�xDn�bH]�հ�-��ND�ō��&	�;w�7�ȸf'�:���ʹj6�h�����c4����mmm��14,��ٙx�H'�������BTDD�wG`����g� j�
�;�x�L.ZQ���\\�mϞ,u,�M��"?��'�t�V8nyh��>@a[@Y7/o��omm�����m4t$'�n�h~6�Wj_��ȴW��G.a}W��(S�yZ
j����7��ؙ��ߊ3�~�s{mZNplhj�ҶX�͑�ݯ<  �������K�E_A��,,���x|��DbP.p)����o	kuH���?���ЕYk��H.y^=VD��^�r,\yե���5[�[]���Tl\�V�p�BB����}3<,�B$���X���0��(q�jY��q�@: �.ǈ:D.--��G%1s� �]ܣt'���'3rs��0�d<qE�H��ً�<=����A˔�4<W�lf!pl��a�0��ǵ[�4�1��!<t�+.�'*��F��n{�Yoo�M0볷�Y%QtJF�������B�6 �:gE��k�8�E��\;��{���smq6�NK6��9���N��^5���>���˟N�t��;-��`�[�ń�,����E��J���ّ����������Ԕy?XF����D4���Y ��Y�_vAA_w����:�ڶ;�
�-�JF!�%'8��e����g�O)�;P���Hȝv�'� ��G���*�O.Lp�Μ=�4mCC�a�wէ��w�qf�!�� R����ˣ��Z�AE\��J�����T�Q�M>'�Z�0H����^�5t;t��O]�0�g+ř�ݕ2��o�B�6�x��2��+��*��L;��nO��Ui�k�[���a.�M��N Ys���F>�7�ࢣ)�#��7M&�@U�]V�o~��礤�I8�����.��[j��66v�y� 	��3H$z&LE[K+!S���;k�&����`��5�1�hA�B�"��
~0��|C���7��#�����֣"�"��"�2�P5����v��	� Q7nj��8 ��H{ 1��5+|�e���y%Cjܔ��x�g*a����s��r�Hdۀ�ɰ�	!��
vȎ�h��1�F
e,ؖ$cVUU�z�+�<��H:������O��o����'�*kL��sɥv�]zd��ࠁaǢ�z�T����_0\���GG�����㴯� � YFn�.3�^u�*_����1���iLL��Ң�������ȭ�5��U���;�?_[�ؐ�]�8)|�������7���MFU�����8L�e�Ú����D�!�x��5OΧ9�|�|
ux��chho0� [*ib�x�"]HQ�c�9�h�0��R (5��K�7�b.�xy���D��tl�K��@F��f��B�����5� ����k{xx|V����HQѡ-V�N-H�j*>>::��Kc��r����Iީ6�����'v��5��(�,�Ҧ��ټ��J�/M�,��Y����)h"׎7�"�
X�}}Z�:-��]`��%SO�Ka�q^M���_޽x¾��ƹ2@7:�6�z�}���+��d ������gM>�g7M�`%ʪ�GJQh(����b\���@������� �k�tq�yc��$<���tt��a����������e���0K��\;�C�aaϿi	��_�,�ߏ&T�����8̑T[~���iY����W�s�wwuu�u�[��k7�̓�-@~����L|��}i�5@.V��7����Ǐߟ������O5QT]}/Wci,��{`)���Ú��p~����g;��NY	Bq�<����z�>��'���������	ۈ� AN�ܢ�����?�[7�kf8���@)�x"���)��)ͯ�>qy�����py ���İTK�Ӏ�;���S��M	�_�Ȟ_�����j���q���1�L0��W��T�5Wz� ��f�g���"No�����_�Va���pǘ�Vtp��Wm
��� �����'o�9�.�o�����4�Y���H�xys�jqN;@G�~}�!R־�qA?�z�#�W��V����.AũdXP\Nhٶ���y��&�.Yx����TE]N�ߦ@��}��κZyX��{���]22�&�eG��Q(}����n�����^�f�����pB����GqS ����b��W��s���d��kX��ӕ�.H�,�~�a���K�wt��&h����/\�մ��}�l���ut���K���j/�l	k�X���1���fG,�;����MU@Z V޴s���0p���"dk��,�	�oh�/�v�_��Ý��A"��sr��h���7A��N�9>���cϼR$[���p�>��w.��z�R�����I�����3���n�KH�f���}��; w����W�D�@��벧����٢O"� �#�4T�Lx8sV�����É=H������ȇ����g.���{��[G�b�O}ɨ���� "�&xW�Z�|���%*}T����3���ǖ��o�ǃ]+�M�^�^a�?�}�}�'�$T����#vYt�xJs�a"��am�{���,^c**�B���:o���٘�_��h �*J���t R9��3e\s%���JN]���V�I�ǶO[-��UW"_�dv��R��}�{�4[0�»�̿s{�j��s'z^]��أ����F��	j&>[}-̗��f��qa�ff7��}�-��� <)~=��>)��%��h�9��UHMP��sj�/Q���:Ƹ�(�r��RWİr��|�����!r���w�L{��ϐ��C��ߕ��oB��� �מ
�����O2,�{ȋ>��r�j3�R�Im������H\�/ـ8=�
��S�$O40,����̉�� �j��	G��<���Cc�IlJ��U�c�\c�/aB����9D�h[���v_�������xٯ+�l�>.`\�����+�kբ>���`����X/��f�F��f�֖����߼��B��,h������9���°G%����y�9��k�7۞��$ɖ΃��\*�M9��oy��=�ϱ�u3s�1k�͔=��J
��~q�k]����GE��=("��Q��/�_�p���|%���J{
��wǈ�YI���P�+����'5!�L>��2+ش���0H�6�'zJ�Hv�42���efb�u� 6����c�â�pQA�CA	II���K��c�ED@����K�`B��AZ��߽���8���Z�zW�}\~L0i!��l�v�^Dt�v+X�ę-���Չptϼ��}���v<%&ygܔܾ	a:�����Mj�!_�����ű���.��Q�n�a/�b(��Jڑ����-Lw��T0�[�-����d���B�	��� �C�XRRM`�O��і�k ���	��g�Hފi�Lt'J�[k�����z��G-}R���\Q�d��H�B��U�2Y~�Mc �⛮<�?�Z=EJ��:���T�FϾ=ظ�,��;x����=_�����A�h]`����*�׹�W'Lp~���`�&���#��j��JRQ�^At�z?�ϳ��r�v ���f�-~�UƼ�����k�
a�.����d��EMtv���:���?�1�o\��//5�Y�ٷ\,���T��U�����T�a݋�Z��|�e�	Vg����̚��u��T���y�D<�� {�5Ȅ.~��R0�pڦ��ɰ��_����¶��)�pU��-:�d��G�7��`Y0��M��*d�������`dˍ+�8]��L�d��/�`p�똦)F����:�D�����u�9���� ��fgw;��N�`�9lY�y���зi�!���{0S�Xd�Y��]�7d]ѣS���p��L��� �Y�ܣB��G������/|
��g�Ye�I����;.�t;/(�n2�~�GiT�r�G��P�5������ wc�����,���>a��*3Y�$E����͌��������nu��ڞ�������Q/�ŗ4�sw3�������n�:�v����7�#E��;κ>��e�8���4���ŲR|y�e�s6���ޔg�R?庞|�c�f͡�gN�ܔ�c�$}���P|C��C�j�U@`E~�)��K��0M��l��\���f��Ν��>�����o=�q����ޚ'j�6�G���7HŗL'~��F�vw~J�R4���p��ЛcV1/b��MAL[�,`�0=�n�"�&}�t9�i>8<�ty��뜚/q�&�eU|f�@ˀ��ɡxG��̟��\���/��M��m�Uttt;X�c�[���B�ҍ���!����7	��-K�V:�Q���g+���;͘3��/�>~1��3k��{e��W�>��g�4�P� S1�kw�`����x��+-+ hB���Ud���Kww��dcN�J��+�|�����z���dRFʓ���mvϿ	q�sFG9��)��a�4��0�ͻeN(��l־��3T�t�ߠQ)�՝Xq��|�阧zbpqJ>��N�Z��OZ���2�DDEK�Po?j��6Л+�3`/�$�C��ni
c&�qV_��G=.s�0����u��v�`4�9��}�a�bj�������Չc�vj���z�ZƝ&�������Ŀ�S83��l+��_x}r���Ҿ#����7��IŢS���c���'�+��^~�u�����#���la�777l�9U�5�i��1v�Vb�V�^����mJWϐ�Aw��U�ڴ���{ �_�[!5�#������$Y�_��$߽\<L_<_�����W�
��a�8:F� b��z.�QvO�����M�����+�O�̎�^����g��݂9��޾=H���3+}k���K���+��C)sM8�T�l���{�M��.[]z�ʔ���뽏�zG�26�Z��a��N��*UDD��w����Zw
e��By����}�#�Dȸ}Ŀ�+l�ϖ7��;%�����G������P �� ����av��$�Cu�/�0b����0�|��G(�y��x&J9���)C��q�ت/污Q���%L��=�S	NZ��<��7̓����qa2�<�k�hښ���a˝^E�q�>X�:�?�|CսU׭oq����va�~���)H���Ӄ^u�T	��m$I0{DT��zlS9T�$�M7?�O�����^fz��
��}�ذR{��-��W� ���e�̩�(e����O�x�I\~���rQ<��:�T*@md��,���k+����UGv�Ͻ�%�����h���'�p'%^��z�20CM�$![��������X�m��/���cꌉ���7��#s��K�X�gSRPR4�Bʄ�?� T�f��<��H�7o�P����������{�_�h��X�}�)I��Z�N���GߏP��������G^���d|�S�,sFv#�C��+L�uP
8^����8Lax�]�du�b�o���G�:͹���@8�w}�Z2"�o<�?�Mu��~�������7�駈a�7A<r�uKO�;A�j����_㜽4V}8�C܏��hs �k�;��P�;D�lnmB���Uz���Ӷ7.W6����c�c�q4_��sf+gO���{�1+KZ��V5��F:��qv�� �{�]��g��ζ4�*9���<��C������b��1���fB��kr��_�/�)j(�nJ�}�E|�ʘ��muN �<N�^L�f$��YK?@-�Hq[X�H�F�,8R���;�~��HN9���BT�e�fw|��ׯc楅76,ŋ�oJc#�_���(o[�h�����ցG�6���#���M�tQ_��3j�@��M��o`3���mB��0�2!�:�$��R�� T�ֽ���Xn��l�����H�䉯4����u�'�n�
Ɔ;�Vpz@��WW�Jf"�5ח##P��zګJľD½���^���Że�r���6,b׽C8̀r����]����Z�7NNf���T����얉X�i�Q�o�U!=��2�l��5������`70c1�Ɓ1�"�wD�?2�~aM�t{ĬuF��p�6�L��j�7ˢu���0>���n�X�)�������<�%���==%��ׯ�|g
�*�_��P��B��8sbi�~���<6�1˗=_srڬ|2��(얞����ͻE���s��V5���Lzd̍�j)ޫ�t+�C_���WY��
Js�[_��������Ӈ��o�a����� �+�(߱���d�h��#�C��;�f���z=Ft���%3,�ɇ͡�*x��!Ld�Z�V����V1d�T��%��aԇ���|wE�/ � �Eػ�U���D������f,�ܛ���d��?�ڨb0	�֫J���#�|p��1�����R!�����?��n�p0;#��;�(�јi�&��T�#mqL�t1����.����o����x��˦Em�� `؂sP<�Oܤ[�����v�3�_�j�D�
�����2��l�����b�
ۢ��9ob9���Ь;>�j�]����쉾��79��W�īI:Sq#I�QK��h���@j�ez0ѷȔ����SP�P�� �k�`�Έ�ϻӢ�A?p9��p�����!1�?�~��"�~o����vw
~�+����$ew<.h�G|�È�����ԘSՍ�����=^��>�wV �Mި�-�Lc�{����[�=d���brO#���ᥲ��u��Y�w8�ޭ�:H̤'�����H�Ww�<0�ǭB�+��z�����=`��' ��^�>�P��������Z��F�L�T�C	�!N	?Ut!�
J �V|��sSp	'��p�殾����������Ɔ��c���]�ۆ41t��k�k�,����"l�U��M[}r�Q�V��kXjTH4�w�uX���yM���?
K��w��%j
c~�h}����7�a���zy�����L�C��2����"��Y�N�S9bA��x$I�L��n�������_�2��nG	�S�ſ5��m��
grKȏ�+� �*m䫩��Mw��g쇚4�]|�ư�W��V�5د��IY��ہ��N�CdNnơ��D���6���ܬ�`^ctx�ӌ�i�F:��y�|E�ʴ{�z�)��P���|PG5oF�8g4����O$�>�J��r%�E�༛mCH ����������/J#��L҆o�E�k�t�c��Yp�޼H%�K��Z���.����;ڂ��u�� ��Ƭ�pfG�Q��M�&,��K�+rU�=I�n�/I���2_��մ�6���Iݑ,+�<S�jqXޟ��h4Z�@�z�T-3��~��z�]DP��"Z���v`������:ң�y�$���R�oO'�t%�ڏ�!�;kf"u5E��]�qe�!b�[�~���E�W`p��}1�ťD0�	f.��<k�`��j���m��%�v�˧�j��w��27:���eԋH�3d��шJ����[�$���^6��O�3���>'�"S�`����xxw)�.<-���N<tmI'n�@6�(N�ް�U����=��+q���#(4�t�U]�.X�%4�<ls��N�|h��B������9=�N2}�J��h-�E�j� P(w����ct�|�:��r}��s2�2��md܃�*7�9�٘��G��!&UB�&c>����:�G�|�<��u���;�����س7��\!�~�N�����c��!Z��}>s�]��oJ�}аz3����&x��͌ ����ܢ�)d&7��-�Mo���*��[�J,���PcВ�������b�Qݬ�b��4����	��$�t�?��Ш�ٽ��K�׿�y#M(��Y_͠�t�iPs����,��9�*�/O#��k��(��إ��0��v�'�eZt��:}��^����(R��2�b��&�=�G9�EC�_j|a���g��z)������g��\!� �y��-#-�R�kV��a5)t4�Iva�����3c���EY_Ϣ�E����M��f+�����!+�Ih|�G���W���v�l��!�,RAO����oN��8O�Z�����I+8%_@ic�gn���DQ"c,�m,�x"�Dh"Ez����'M:��{��D!����m2�� ��b)�4D�ƫ{S��N]�H���'fΐ�Є���t�ޑ�n�v���*�g��eV0�A�~$?[9AEa(��A=�5���Tux`��Up!��e��Nh�����U��E؏��ĬTd#�gj*+��x<�i��yv�U�`&�.-w���/����&�����+&D�r�SO�\��*�����/j7"ݾ�n|}�����4r���� �^��|l�=q4����_<=H�nL�fAA�\||��P~uaha�:�;���PS�E2���x1;�CK}e�5����S|�uoCI�o�ϣ�h2�A�p���8єX�G
W�U��U�h�l��T���(��o��6I_V��5�:Z��z4�X�~�iG��<u��|�8��MU�0B�5v�Q�p�;�����I
��(��CD
������`�>��5 1=_��2*�<]=Q�^�iN�t��J#r�B�v�tJM���C����#5$�?�rj�-,���.|��$�I�R!�8+@�?3|��NX2�n��{fG�������%׏��{�,S������Ͽ�6���G�;����hg4W7��1A�Zd_��˙�9j	R��G>��P�q�k�\��L�:���q|H�V=�����M/U� ��81>ZUKN�e�s-�N�!eG�iq�9�{�;7�l��Gs�/.ޣ�
�wgΎ��꥛}�������6�[�h
|ErMqf�:�<�/�u��8� �K�U�4�1��R)ð<\���������2��]/	{ ����$G�hp���74*�d��~���Tl�˜���$(gb����Y�4�b1l�.�� ]�;�^�r#�ۛ��)��R�ϷV������16A|�`|���C]V
�]K&�Q�
��qJ�(:�tSh�7�)x>��t��+�&L���c�!X¹M��`�
�/��lf(��I��:~0�Eeb���q��A����|َu�2�q}:�A�S��[o�ͪ/_*�!�t��ɼ�����P`L+&ox?/5�
���b�f��|U��"�ħd"��Y��W����Nye5b˄�������a��0*�Р/%*$Ѳ��X�W�Th��TZ�xrx����l^��b�	=�r�����Y-��Z�xi�-�l����b_�'������%�VP69&�uJ�D���m[*wf�vU�2p�v�D1�N.J��� ٿ��@�b/��o�mm��N�j������Սu4�-�W��=lw�7���أ������E��yt�T{��v��T
D���R�e��dTXÌïga�/� +_��zeH�'V-3V �^װ�oY�v���9)�M�~!�-|�N�H�����p*�8:����R������N\�c,��=r�P�5Cg�ۄ=�>�?,��<b@�� e��Hp��?D�]�������xg<?[D��B�A�R�dNEzXC�;���u��{�$����I���O{#������L�i�I�g]7�% * �ga	g3���>�g���ѹ'.�h��E=	���J�񓪔����z{���2^�@��r�Y�EdN.�8�)�[j9&�p~6Azi�ٟ������|���@��`��	�����59z�M�l'�|R�N_��)3?�nw�@���
��bj��[B ?y�o�0��R��Uw	Z��e]��J�P8.�����&$��f��ɣ�K\ X�H��/�?	̢�aR }��ւx��̑�Ң�
�:�d~�2����uw�؍����jM���ǯ��h^�ϛ���ə?%u*b����k�+���`�0/<@լ�>ei���F�Q�v����dH6��.@N%H��ɼ��DX�����7-������<�>\K���'Yc)��	���׫\�Vٓ��T;3�p�;���'�~�0'ҦqPƟ7�$$�b��+���l�u7c
|�#��AE���g�C�'#k$PQ�����헝\#�feO2d��q��u�m4��.��������v,�C���K̜���K��,9a9K�~p�Z�7���S��$�B��۩�����%���R����(~9���o��3�E��5?�.��u�_��>G}��q����W�9ɖ���&>~==��8_F�*�R@���7�Ʒ��2�������-�۽N\�PT.����pv|3���y	���a���F!�%u2��� 0�	���c��.z]������
�d�}\�M�<\�YP�j�/a0j���b��$pz�f�<f]��wNNg,��0ۘ9hv�����j���zkŭ�7�j�10׳>%����<`1Yx3���Hd_���� �f�P���w/�̽�q��9�}����m|ʵ9�r� ݰ}�#u4�x#����9����p�7��Wv��N��c۹�3ot;�����H����w��. �@J��+���ѻENf":W0j�g9����K6����ηL�u��ۆ>� ��s�^��
��%��Wǈ�@Y��^��n�|P�H�lD{��[����Ȼ���`=$6l�H�˘��K�Ԥ�(Rn��n>���V(d���	b�˳�.	��#=��j�7@J@s���%�Eu`u�3�97=����}���@wTTe=�W,�����*E����C����R��M�𺔗>6n�&G�S�{�jʒ���+B�?�@�REj����_�X/�@��?78��H����6(��a��r"���m3l���)xŘ"�x�{�i�:��sÖ"�h^x�<Z�Hҥ�J�>ۏ��&6"��<�����F�T�����Y3-o����aX�Xנ�7ȳ�E���[�!P��]�8�ք��VO�}�y�~�����i:��9��p�v�H���(A�r���X|��-e��������^f��*3���b�K�w~�R���n|}���W������Ne㓇��������m��H�V�`�]�b�:֥�K�7`zO����ᡦ~nY�vS"�'/VR��gF�^�b���4�*9w�G)�!:7Hc�ݮԱ=uHE��T�miaz��������L?%� `k222ԓ���d~dI�MC���X��zE��i�Y�
/8��6pP�nDJ��P�'�ܩe^�l�K��x)�UG�!��֢~�Pf��[ �C]��l�!w�w��pm����ϫ����Z�p�J�t�����XX�-4�1N4�e���h��f�"v��n۝��['I���=�?8���2�.��C�?�|׆+I�Vw�f>�|EM���m[�}����!���{�>�ȧ��'��K�F��F��o��cX�X��7�3���lrP8͏_w(I6uo
~X�sN��
�Z0���L�?W�0�X���2P�si��/�=�\*����_���g�-̝ʴ��Ld]� {"{��MuG���CM-��@����)���-w�a�Lk�X��t�%�8rՏ��߂a���,gRcAO����p���4ief�~7J�g���v�v�:	�d�	`48����e���'�6H�Pz鄮�kun�M�v�H2~at}<Z)�� ���d�^ :�f[�g��W}�UXR�{�Բ8L�_#"2��b'��w�	�5���|���4aՉ[�C��JXҕ=�����n��e?�,��?a4��Q M�5��c9Gk��m��Z7q{�_E���r���OXoW2�ş��xKoM�N�Q,29e�𐺩����;'QS/����[ki�LI��a��cOM����"U�0���,�F�P���W:ŝY���2.�n���Ӟz3�[8C���H��@�ϛ.L��\ի�^N�*9,O�an�,om}z�h����g���ɾ��R(�9���n� �H�烪)|@�!|]j�Y*a����������ަ ()ϊ���/+���{�<��*.U4��8�|?ތ�Fڔ����e���1>�yָ�wZ����o��N��^��+{wc�p����u6\��~�y���Jҹ�wr���f�5����ZO|4����A�Ԙo�()+w���/5�F����Y�����E�/ARL���7�P)^����|_܎j��!Z�W ��;�:�E�Y������be��&�[��Ŭ� v�*���p�{��WƔ)��/�t���q��b�_��C=
��ߤ8�uDf��rk�&l����vz6mUԿZk����zGy����L�fg��U�hk�q{� �c�(�_~�U"��R)��[�Enj�`�_;Z}V��$��>�}]�y�֨��lV������� El��0i�e�A��-���G�K���v�M�|��+C�_\�A�2%���d�������YΨ��m^3i��\��8����t*��)$�tP���Lz�mq{z}�1p��0J8L�����{�k���qfW��M3D�M��`�wpq6$zzzԓ�� Sʹ��OQ9_����<6W�_>�I���u�=Ԝ	����p=E����Z��k��Dd����܂��'���i٫���3e��z�Y���x�X� ࣷ���M�VI�������S�Ӛk$�� ���]=%���O��Rs��{�E�F�/�~��j7*��\��8��Uq}=�~joY���n�*<z��#���-Ʃ����cW�5S���Rm?�>V��ӧM�[+�T��U�
��pz�<o����;DD���/I?�o����pv~��*�d�.n
B���M�?�=�ث��
`���Y�Ǌ���F'��������@��?O%�K��5B��L���T���h�F��u���YE\��&�g�񢗌�������V�at���m�ve׸�� wڟ����^%��"FK���� S���n�Exw�3}#r�i�+�ߣ[ۥ7���˜& m_��L�N(5����"B�i�b	С����� .��ç�TA�oV�=���J���$Se$f�ϵz�#=�cif�n_�(��.��ģ�\`��,�$� ���}"�Y�'��Y1R[_��$��R&A:Y����V�=+��+�����s�����S;
���/��Sr�}��}�k>��3�|�O8���I<�W�v�2�w� ?i}����Q~33Ύ�Yqs��&��`L�e�xg�_�Ɯ���Ǐ}�)�r��W�o�Ǳ����2zƳx��������[bp�Ȫ+����x-�/�.� Z�ń��w����-�3��v9���Lō]�����(tm�[Ϫ��X���d�/�^AmV�0k�K�?G��ud;�Z/��q�T�k8��!�����BppX����`�S�G������3?[- ��N�HI�[�d�UN)��e�Um�OD�%��Y�j��W��σ/�W��,\�����ɟ����H�!܌ΔQ��K5!&��iU����E�4�{�Ͽ������F�FIc@�u�b�D��T"���Swj��^@�*8Ik(pp�y��?7)X�0]���^f�L�e�G�@�M���+**0�$�(���6���m��n<����TBW� [i���!c���P�22�A�]�&��1_����m��V�@S��w�&��ޣ�t��NY?]�5��;�-:)�r�J7����
7b��c(�����doyh���ygR�2@�IC��T�P�;�-Sh���s�y�0�CM�[����DL�1����q؛m���v;O��2����-C�OR���� �y�:��|�eHJd��Ѿ���3+t�#��� t9,�����T�F�S*:���Ɵ��{u��+c�3��X_M���q-<����؝	�Kk�C0�EG���PS�ʞ�d~��\� L���L��V=$um,�����/o�)��h3��a�ʷM�2�F��լ-�,�;rLI;��GWL[�����F�6$�MU�-��N��"W�w(
�^n���i� �׿�M݈ ͙���в-����n��h!d
xoJʭ�����̾�V_��@]�MU����f�*X����o�I��R��5IJI�G����'�.�'b�|�� ���E��=����."�4����za�Es�xĕ�ǿ|&�/ ����h"�k"��X<
䲊Z�����ARKف�S7���e�[A�-�mB8RSQ��|f-$�!I�,vr���-�3"t#P)�r'}	W�Ж�^�s����cϞ��J�ޱ1�w�K.Ҡ��W���GØ%�*��~�Psc�;���S�I��7\SRY%�۝&:cGo�ǣ���*#)���M��������d� s��G.oz'��r�'�x�H �����~�q9�xg�;�{��wJ�:��mi�
Xr5�K�����6�u��~���W���w�8eOvg!�/S%�����|�뢡g�CCC�Ldΐ�J�� �$Uc�h���)�IG!M;���d3b7��ޕ�4ꁣ̯��:���ݔga�&fp��*>H�k6�d�[��l�^�~��q ��=ɼ�>�:õLX�M�������;I�N�Z��Q2�p��I���]�r�"���wK����LC�>��ՙ��'7St|���9[��U����NQeU������5�DH�`����Tu�g�Uљ͕7k������޷n�tD.'O��/��-���+R���˷�6��/L�[��}���`'�^% �����];�Η~<�O��C��	���:�Iß�x7$�w(����S�ː�[Lt\ry;��rT��"v��|���)��o���S��+����U��`B������6�"��|y��V:�"7�	�w���E@��[�UTn�~����e��$��"J$����چ/fi����P�7�D���BYț���k)����Y�w�Qa)�h��{ts7�B62�8kZ-{ ������q����O��)�-F��)��]*�)�"�
=/��~�m��6�=>J����S�ȝ$�ﵟ��>;�.c. �2l����Wg���Nȭ�2�L�X,��cf+�N��>2�1J��#l�q�������c��b�h挕�����z(aސ���z1f]~UsRy��æ�ED��_�T��2�v���h>��ʟҺ�ugu����1�6�7o8I���f�Bv�&��s�s���`�ՙ�D��Ga�m)4� �����#B]xhIs��᳣�Ē�A������QF��aO:/|R���h��.���bn;�?�9�����DA�[ZL�euu0QO�}}�'/��)R�ji2�~���=p�d7�a��;��m�P�,%1�NX����XJ�bTA�ɻ:Jr'�g^�T��Z����Z�e�mK����`e3s�]����i*Je�n�N�f�Bq�c�A�켸u�qRjy�c3�_!Kܺ~� �Q�-�6�oj||��/f��МS��Ϝ��+}Ɍ��!v�6��K��*�T�p%��e_T���)B���R���s���$����墋4:�f}������n��/L�Ǘ��4�i��n4�`��2ձ�O�C��&@]���1�9le��bkkK�1�+�Vy �JJ�l���ˉn�$���co[�w�y�T���[����b�&������1v�7�Xj~�a�3�X>>��6�������Q�l^:�?Թ�a�
��׾���;�KS���OL���UO
�k���ԟF��MV�n̢i"�k3��W���߸wZWL�5��M��ͩ,.��^�3s��~��=ҝV�k]VX�/�������WH��ݎ궀WȀ����~���Dz@��U�^5:� z��-��=xq�S�)M]�r��&�+K� v��d啽���cR�	�x�V���*�� Q�X�o�\�o�ᦈ䤊����HNR��|�7�p��1��A�W�Ԗ���-�i�q5RG�mT�me/i���z#J*qZ�6�eٕ��#�
@9Vb2UR�R �Z�L��Oμ[��\i5N~�������T*���E��zd��>&� 9ϧQ xb�WSk��aC�S�$��@���%9��$9O=Q�:��0�AVo��Q�5e�$�z#�4�7Y�܏CR%[�x� ���G���I�'.(�!B���,�^�b4�{'y(B<0$F�,cX�$%=��kb�=2��#������R��mXB�&��y^���K������I�,�d@|���O��1���UeV�v���B�6��n_�+k��&NXM��1��N���T"�P)����<����3v�no�Sp��,A��������'��.!�G-B�555%�?��$Yt�o��L`c GSqOܩm��S�-�tF���IxИ���-�_�g��J�X@f�̷�9���8���pN�upf8[9�{3��5�w<��t҆�٢N&�,��jHsĹa��J���1�8��I�k����YsHQ_ϔNX���N��*�%�o������r ad�d�!|��Q�p���؋�~͙�Fk2W54������+� �a^rl�I�������X�P`@��	��m�績�B���k̋q�>iw�=ig��Mx�F�l���,�-�����X�������</���c(�*=�w�B���V.�(]	΄y����r�>�0���r�D���̈́�/8����2;���Pk��V:t��`�#��5-�������O��=���#�xfe~ҧ"��a�����J}K=�*r����0��3[�������+��1���*̏�.�.T&#����EUز�N��+��rpp� ҟt�����$�	�@�\�II:e�P�C'�Sd&yBzۭ�΍��2[���FL !���C�������&�j���-t>��]�R�Jw��ʋ{oi�r���ʟf50�W�M�YOA�`���OeGй��[^~��GU<P �E���u���-�QW�U���}�(+��4�߶���-�H`��c�h����}2�%Sx�ppP��wQhW�o`�Ii.�����f�)+�7�i�����'	��&Lat�J�紥C	��L�Ez�WJ���æ���Z<��������o ��T�m��qmY��*'mM�ԏ:�]+^��v�.b��7-��@<��H9�9�8�"�0�S�|�ס����h%�"�;�fz�<�C�@�m��w�3���U�l��{Q�?��Gm���_���!�3$sA`�CK��	����5��J���=+�IX��������|�ᓴ��2�ˋ\Nz��C4�{n�x|�����ø�{�T���&��R-�C,ePc��EE���;#t��Y07蘯��H�SM�6H���Z��'���Yc�?~��vw|�ː ~�[q�*��淵}���R����$_�N�$?�Ec�е ���<���r����V�3v��0�X���;�r��H���m4i)G�B���P�Ǚ�t�ny��|}��1F����1K��|�y���|S����&N����\����AZ�3���������4!���1:���v�o��2ǌ!��M��ScYͶ!
H�2�AB������ZH����I����epP��S�N1�:�^��/��&�.ڃ����7��>�qP�>��uq���:z���;ɌO�u�)x���C����E�� vp�!0S�������������z��(oGhՃ4�VC��ܷ2 ����y&���9N�P��<�s��\9pՕ�������g�_{);`s��ڷ��G�lzsƱ�kW�)��>V5�:4qF��v�8+�B|SLA+<�g���t����)B%���#�O	O����D,�8�a
o8Kf���쁦��iI%ھ�I�G\�YI���}��	W���E=�F��RE�Y,�z�z
���D��^�;��a�mB�f0{��6�l^
׸gc����;�z���1.����&|j�P��M"��JȠ��B�Q���]��]�X#�N�P�쨒՛N�XSc3k�%>%!�̋��*��{��sƉV�N��S紸�ay��G�6̟�z�����F\�G��ݶ�`&�.�j�Bq�_��iU�b�ٷt�Ȝ������j���v{������r���R<�\�����G��m{ӯ=B���d٥�k�m`�"�	��h�5������[���l�Aa�K�򃦅��Q�ʨ(��篞OUm3���Q�a�udE�9c���a$� ���@�K�
P}B��w����RՃ�J*;�V��/��M_7[}C�����'�m R��J{ 9㺮�u
/W&�.j9y��zu�N��d-�/v�U��#+}f����A���S6n:�I.��{M43Uc�B��c̘'a����|8��1k}�+��^���q�������lP���Ycj%�t����H�|�ѡ�'%?�3ir�y<���#۲���W��5i�O���	�xO��Ꟈ����d_�\P9@���E��@����<��mK��EY2|�P��p��]�
KB6��)��VJ�x[�dXQ����ї�����^�G~#jR��q�nl|��^���YE�\>@�z�)z?��on�;[a�Tg�n�׫��[(��|�mq6���>���;cƬ���p�J1堰��U���s�Z�}�O��� S�7����|���Ld��݈�����KPU1�(c�}x �	v���Q�����P�q�\����6�ӣ<�y����$��	�i��ЃE?嫯tehb����;<e}�{s�v�;�\��'Y��~����]�6%�Y��ދ�p:���))/TdͿ}���(�dU��.��
����x��:���nQ2��5�1PE�L�ή0.��u�j�[='M�g�L���� a��:�^O�$-���� �Z���bQ�w�3{����|i�R�\��殺�l�o,-��w�]�mg���KצS/���/?vx�oN��$\�j�x/W�zaRɻ�K4���Ѓ��~Ҁ �ZI#��[ ��/u$�{=[9Ranj��)�Fս
�s�˧���� ���k�7c��qӭ�+	���\�;cظ�軒�+[ޠ�C������i%}�����k���Y0I����	C�QLϱ���6v�N��Cê�!���hگ���8n'�|τc}M��a�Bb���˩�j|�Y���DI���J���v�S�1�	P��$h��Н�{������/�FU��;����g�ff�2���q��H5�.Ս��P�-ҟp%�KVi�%lN�X�͠�>��G:�e�UQ���4=�d,z*
?�/2�j:�}��u�n: �@���&���Ⱦ�Y쾣�N�1}4jl��9������^���VL7R��s9�V7u|�K�ԱGIq7���M��o�w�z����e�O������Λ[���i���@4���:Ik��Z�j}nFS�)�D�D�����Tm+/�#�֜F@f��iN�T�>�	=��!y�v�;�����pq�)���<V�C}����Z�En���ޗ��,�"�!�+F��(�&6C��G��N�}�8C�N�d6Gb�a��-�����$L���w>	��"�s�RD��msy9��yG����e7 R�`l�_�Y S�j��v����[�ӿ��_�|�G&x������@|��S_IC�z��:��|Z�-b�	r)���o$ p�eΔ/���9о�;,#X;)#@���#ɬ9��T[�\�2H��d��6��oŞ;E2�<^j@�1�s]�m�m�/�.�ڀL�7�tTZ�.2_�c��ioOO�9CX�����4�����z�$���tUd�_���)vB����v�Ah,��oR�#�a�YQT��O�U��2~�1�#�9�?�[k�j��j����� �>ї�����^�������B�������Rgҿ�6��>��FBN��%��������?��LR7mi��|�޻6����qc��xĤ�d��N���?Be�c�!�C��sW�����V�BW�NA�S_�S3`�.,�o�P���-#e�N!(&⭌���ﳪ!�����)�I�plCGUS�a��1�,X�=���H%\P��J~�sw>�k	1s��5�g�_8(����������YL��r�z\��$o����wk����x;���ҩ��ɝ�S"Qt��B����J�N����h�:���y��q�Z��nt�
�I
p����6���3�3��Rq�R������~�E����i��6<��O����)���숎"�¸6Nfje�*w׆�o�
�������q��v�����s�S`����4����&x�������{Å�P1h�%��D�:D:�F:Q$��c@����n���o�����k�b13g�����y����	P�#=`�Ɂ���D6Q�۹��w�z�F<�{�?��*WE f>�ҹ��Qۼ�D�f^�}u�H�g2��3�K��l��w�KH�}�}c!��� ��y�zޓ�-��D��O�{���u���v���}JG���R~^aup���O���uՕZsEU�؆"�#6��b��o�Oha2�=�(�o�C���F�=K_{�knI��@� tc�u�b�a!�̡M�v��j�;/�?�m$��|��0T�������j������9ݫh��q�U��Hi~��u+׾�j�t#���v�~v���Q鵌���=��6�'}��~��W5h�#x�~�ޡ�[X����oVM�n��z��*˪�g��[$z�B2����u�^wU�N�'���*�e�@l�	!�?��J�|x�A����@����թ�ї��eKB�)rX��<�{8�8"7�/� �
O�r����]5�����w���[��y5fi�q��h��q�bu��ջ�P�r^��M1[<w��>>�����>�S�/ ���/��?muCK��ǿ�z��y�q<��V���_u9��U�b�R8hJ�w�I�YSkf�C����cJ��h�y5���)��u�����=O���;�.ͥ5BS0uFp7:I۹qE6����P���^��o�5U����0��V��q���Bg�q�2�kbA-�f&jy�?���O�}_b��U�a�%��'6(��W��e�����.=N��_���n���8nLi�tz���/_=9L�D����#l4�a�N|�O���D���=���u�>&�HSWD�JT~�X���a`�IV�y���AJ;j��t�O�=tG:���m.뭍Ķx%�������Oc�78o� Smss9Sr=%ཹ[u�� ���%g��y�ԙt��s��Me�z�+M��~� ?/��t��t~���+`$IEo�ڃwP��fp��'��R3ݯ%qbo�ZZX���}���\M��#�P h�I.�eq-���?��~�hbL�e���6�ݳ}d�%��Z�E9��{�ܝb�KVQ��̩�j��M�k�ۺP;�����wrK��:d��ٲ��4���8�:4��.H��$��{{s=[��KTO(��G���g�_w��g�9_�u��<h�0+�ve��`sW���\6���Q�Gυ�����_�ka�{ȼ'9��µ:TV+�ڂ���\挠��������'�2�!4	'R1�w�*��kz_΃���N+�8g*�z�xΖ�繫�N�7��cO�,��R���,��$��N��Ma:��X�r�3bv��|�v�!� ?��C��6��\�N��L��7�{$��]�(T�S�_����H��g�w.~��C�h=g7�G*?�<C��U�禲���L3K��:X�ߺ�q�/���+=�|}EV�3�y"��mo��0��vn� v�vN��[��ea��Ç
1t�2$	=���^3+Ͻ/!�c�Z=��)����{cǏ:<hƛ�9E�NH�h�u��"���qyd��:5�1Kp��n�4��u-.���os�~��'��jQ���H�@��c��V�"Yk��v{�^r�xK�y$Σ]A �{3Df���l�&����TO�^*.��n�v���>,`��w���љ5W?����j�"��\���lv��s�d�t�ٴ`R��6��g	/"������J^�qr3boDD�z�^�?�N݊��h>��~�u*tȱ S���^J)�����-!�@�x��<���	�]joi7ň����nr�������ٗ<�+�t럤"nl=|]� ���;)����F�ۑ�A���ȉ�I��Jb�v����a��B%�x������~(US���e����i�F������2����#	uA	��Z`��V�a�G)[!��X����q��.N;H�?hF0(�z�x&����>2�
Br���c��E^��wb�]7��hc>Rpf}��-�##��qi���Ѱ���LH֭
��7�'���7��4��#W~�������**+w�bi�ܺ��1{ָ�^���˙yO䪋2/OV����b�Ύ'V��	��	�|�lw�X�M}��Xȟ"��j�S�j�p���0�� �4�u�?�z�����#$��9����nG%�P0z�����k�*��G$!�l���.�g�d�%F>,�h�����G�8���9�܃ёV���I{�/�����:e��+T"�2@�%Q�u�s����6K�h=B�^�����b
�8��j��l���"C�R}]�WHk��P��}�7	�U�T!h�X��"��^�83�[��G���ZFn ���^�]��l�a�;.����uU����Z/a������0�/3����6z��#��_zWaw��sۃ#t��N^�jX%,�C��;�$���4�M��<k%C�P�Zl�â놉��b/wz��nK��'�wٝ 7X�����ׄBS�!�=����+�~]�h��:����Ƴdj���R;�~���uu���ou�%'"E��������S�r��!��\z*uc͓�Jtc	Ϻ�tQE��>����4Z�z=�����~�
1�T|hx
-���4�Qdddm&���r����W��p���4DP��OT��k/2{dتm�%$@��g˖}ڽOoSc��e�t
Q�c���f�ɂ��^�YMZ-�@���h˝���* Þ�_j@�cn���"��W@�=�h~�@9���r'����M������0�|�������蛷F!Č>A7�,_H��t�2r~m�&�5����1�"�LBtEB���g���J]�[=?)}oe�F��ƵA_�c��S�Pe��;f�g�Jb�RV�����`��V�k_�	�b�m��s��a��� �e\��}�׾?�(n���N����S&皌����Dx.F����"���Ԙ��<�4�~��� ��Ɔ%	�����2��8��w��T	�8h[�2G<6
��)���_����;K��J����uz����9�0$��[�J.����5�aSz�k��Q�2PP,ad�?�dۓ�$�]7k6���v���D�����ޞ>�5�e����,V��-f���xIQ`s�З#uc�5_]�3�l���� ~Ծһ>b��=­��A`��t��F@7�$9�L�K�{6=�/|%s����.<&#��f�ws�<��/��n�~l6H�H�%��<jߘ���b��/$F��k:��~mE��n�X��=_���Q,e�0��)�U7���N"W����W>xܭ�X���=���433�w�r*	�#�ۮb+_�ܙNɘ+��^��=��N����c��o�����
��]�}�������S���]�-�d�፼��rʅ^��|}��Ӈ{�CX0�y���K����E�3�Mα7���P}�kPr�u|��{#���O3��0�qny����}���CIT��׫�_#R!&s?��`�Ų���x&�e�2������q�F�SI�
���/��Bd}�����ĸ~zb�:O��Zh�쉙�LL2�FL&)�7��ӄI-,,����T��΍����;M��L�����G-z���Y��Ɣ=������x�|O`R�WX��D�$�`�$i��'j��&&&.1���jͱ�cs�?���2�YKu��J�d*����<���/�����������t8��Dd���x_�LLmp���9�ٚn�~pQ�p͜2����J@h��v߮)wݔ�����CS8�d�2k��� w���-�7%2(FDG�"�Gd��=��%��T�g~���}�!j��A�&��UNZ��B���d�>;����_�	��j�'%?}�S��}�T��������ǐ �yF�����ƌ�ĀoZ}:N����D��Q=�[.����q�y	ON�r a�\�=�PVQy���������5����7��m��<z�����%�~L�ðVcĽ�i��Q_�"�E�~Vt4����ks��[~T[-�@���M������e%U�| '?A!;"Bl��A"��ߋbUK�Yތ�����%�����?}y?	�;7�G&af	�p+T^��_�XZo>������́_|^��۷%S�AE�Mi�+��ݚ�S^�.��Ræ�!��.��5�~U6È��M�B�R����@�4�W���3��B���~Wʹ����sr�z�'&���{]����g��,�z��K7qu�<���1_���B���72鈨'�������ǯ�?&f�P\<�\|I����(	�8SI��|Ua��Ic��Os�EyY�*��]�(��ؒ4�J���į��+��14Q�� w�S�/\0ZE���QX��YFł����Q_�B�#0>�b����b�o�35c��+�͢9T����S;�������ġ,/��G����T��X���n��֘M�������eLbgl�R����U1�S���ʩ�� YTq�*�[�HO�ߞ$�Xg{���B�t)�q㟂����Q�������������o�d}�آ4�L���F�Ǌ<x"�-��:�6M�`��,��W�|Ҵ������-E�JG���n5�'u��ӕ�	{)�틣:>���I&��΅���3���v&ՇD��0f���iNQ��p�U�do,�J5"5z��҇�>��`��	�ٲv�}_��	�̂�|f��������O��؀�_���#6.�]T6�q�ґ��Jvr��6����KqR3�2��V�i�	�??�H`qZ�M����?�kg���%&n�¢����UUեI����<�e�jg���w:��;̢t�ጷ�7&*�F��uYAA�Τ�ed@��֨˴�F�c�;a�`�4A 	�ݓ����44L��wX#v�0�f�SW������Q��� �����U�r%l�����o�FQ!�}:䈕u�^�6���"��P�.1<<`k�+e��#�<�|�S΄勩�/_Rrr�P_:���{ƫQ4�$N��6�Nܘu�+����f\&�V��� ��T݆�R��SU���#5�ts1葉��́���8U$%�P�����O�o
j�����ݗ{Ll/eB�͉���z�d���
����-bjjV�N�tj*��r�>�G	�h���Hy����I�"���s�SݽV�b!RZ�9�����\/'����	���'<�~J���{މ?�����KWA�I��߯�~�<�����ǪYL���H�I�JfZ�d=^˪)[��(�f����P��_�K�C#H(���W�+�ʙS�|m�bA���ۺ�<��
H�K^q�V��+)��q����(��\$VV$�:�?+�y̖�߫-i�L�w�݌-�������Z���|,X���o{G�����X)����d�jG������>��E�^Bu555�&�+�%�RJ#���g}�&�R4��?�)Fŉ�l���Ulm����WX��<����b���f�=���!�:����E޻��/4�
Uq�׍�����î�)"*0,�m����0Z7���v��'��	�$�f�@ �M���nd�
u���ۖR���b�����eo�hE�ⵃߤkOM,,r;c��	�8�I|���x��"��v�fE�>Pj:׍ONF�xi�ꑇaV�d�H�:k���%��6Q�U��!�z�hj��1f��_g��4�2ng#T8��K�i^�7,7������m��V�z� p������<�)�I;�.��s{;A�%_���LV�E����n�A͚n�׾����v�����Լ������h�I��O�o�YTH�TO���"ؠi� �jGp�f�W��<����ն�y�$��֟ g��2�T%���$�G��Åq�ل
jAF�$<޶�>�>�>�[p�v��\��B��$�#�j�`"��e �ݱ�O�'�-"��/��X�PB���蕬��v~�P��>G5��u��h�3e��<����X�vl�������c0�)�������]]��Ϸ����E�b�n��n�r�7??=bfg'lw�5���KJ�����׺|����_Me��Қ[��PU��7:���st'�����Q��Ҳ����tr�]>pD��u��l�>��zF-���j9¥'��T�(����r��'�P�^w�O�)�'N��l-�T2�]�ǝ�ҦL$p�q6�t�{;���T�0�if�5���u�G>�ǏR|
�j��VL&��j�\��9���d��"+�?��{����!�h���~%���U�V�g�r���yE2�su����"
���������ܹ19�6��,�)���%�;jF�>т���I��5ihi�V;.Y��YX��V.�����Gl/�x}L��E<��(-Ws-�k]{�M%S���]�Å��������ӑ����$\e����8R�����l��s���W�h�,<���7��j�x��ng�tPr.�>==��KC�+: �JR��o�i���[\t|r���\����OB����Xܞ�	����3��g��1w��i�s&.�s�l��Xt���)�z�B.�K,��B�+��]�˰�(�����@]�u�(��kW�����'�`u�u/�Cd,��1�+����ڶ��q85�q�k��M{�䫨E���y���)�/�s�h�����UWW�O;�'�^��K��a_	�}uk�u�n�u�:^�Mr6���1Ԕ����@B�G2�z��ݮׯ�2� ��Sj�c�~j޲����Vͽ
A���CT+#�v���y v�G��v�N����H��59g�ԧ�d�p��ob�Aܓ��l3£zYs�r���h������87lL���m �h�׺Q��Cd����v��hm3m�띯M�>�����v%	鐑5��1�hVz�n�B��z�gX�<Q!�����;��P�ƭ�aA`��EW��O߲j��	cdB�]�z]|���I�����V��1ޡ�μ..`��s����>>q��K���)ŗH1Z����8��T��Wo��'���� -��z|���To�]�>��4u=n��	/-�C���5�ݤ�G�q;Z�e ����H"�H;�a���jb n����S�J*�bl�>&�
��u?�J�EYl����>L�}9�۪��h'%`ԇ���c`���!�#m �"���գ��׹u*����.3g4��v�K����U�@B����#_���uA̯u]�H騣,��%�B
-�݉�����6��c��>�'�VV�~��� ���2���P�懰���A��넒�t�њ���*5�\˰���$����|,_�Y��Ÿ�dף���!F6
w��� ~u����S+���d���W�L�%����N(�8r��8�.���m�O���no1��rw�+��&�F_�2�p��(�k�4AУ�p6l+uv�zF6�P�е�Yu"��2�Ь!p���4�������S��d�"�c�����u�������~ϫƏ�J����5��Ӽ1�TH�R�#�����j=��9�q�=���¶G�ȵE�WL�~i��=ަ�i!��dzҎ�.�W���cЬz�b�[;}�%%�e���CPQ��4$�
p�O�>ql��*+��v~��  ���n��?'�~4=-��=��ܝ:U
��Ws��-Q26o�A|��)�_y�~����4�⊿s��$�gړ�n�2.����@x�q|k�B׬�ۏ��}�g�����<�[(7�Q]�)(N��BݥH���y��C�xGk-�XӮ8���7ZÀ�iwEJ^�2k/��;q���n5 ��'�������rx��V���=���(��is��U����0��Pi�#��0ř�MAQ�㪫�6�B�̏����k��?��y�Z���=O�
�as��m��W#,��_A�n�ϫ��4�'N
34ŏ #o���b����ڋb!{4��_����m��Y3�;���q� 7�a�ڝ�6�}Eʅ�	���ڛh1��@��wvw�c	�e���x����=s���c���U]�0�����GS����@�ά{���7���4��e��x��^���X�}oY�n�������D��������|�ͪ�+s�k��/��|� J��<n�{K���1��Y��>���k�(�� j�"e�1�/���Nv֛\�	}U>�.</��%�&.�~�l�kb$V/���v��h�%�`^�h���Z����o�^������d��	��E���͑0�>�� �7:R�9H��naϹދ����4�N�Z�����q;:���W'�ή8���8ʟ^Ss�7\!I�b�|"/'穳��Naȍ�g�v�+ӻ�u�k}��Ž
YȖ��jM������>)�ՇZ5W}B���J��"��h�~W�:;�A�w��c�~���<�\��sӗNݕ��E�ۧ$�����|WVE1��lwb&�n�3�a�JĦz��6T@���U+u�ϱ�c׵�?�}�bc����'����z��H���U�+��fa�=��/�)��ĭ+tq�����rQ�4��˘kT� ��u�������q�2�@��j�F.�+B�ޟ,%{�\�������������,xJ.w���%�N<��*�t�l�S�e�*�k66F^n?+_�"�@���u$�c�;��K��
�7V'^
����x�E�S�{��'=�H�|mH�0qU͂�Jm�I�Uߞ XDO��0b�ᗡw��<�>q�f1�W�nW����c?���ۘ�_�1"'����D�rD*a�i�ŷ��ULQ�Gix��o$v�p�1�0s�6��.3AJ5�)��g�P�N4�5�{����Y���9�8곔>`���_����`ƭ�}%������A��!���w� A�ѹ� ��?a�Hzs�`�5����mZBw���u��_�jOG��kx�N�lΘ��d��V����J���j�䌌lŏ��N`q�8�d��F rÀ�u��}�V�u��P�윗{��Pe����v氩L�}�����S&ߺ)M��
�;[�hf?��VY2}|�G����f��Ft��u��Rx�G���t�/��p;���7gB^?U��5@�_�`ZE�É�Vk�[C-��� B�!��[��9D�NV)��a�i��l;�a�߯�����H	<�J�km4aRvg����7������/ۈ~�G���C�s�Xߝ�9J�?����?jPv�����?��y��UMd�Z�^u�)"��7]�%��:��xK/.�P%:���2E��
�;�nS���V#֬3U�M��F����j��jY����^�}}$<_����In�}�(�̴�Gk��%%%��J�[	X�uf��_��	&{�|b�������&R��YRd��m����i�g!���3��w%4^�s>��T$b)�ڙ��*������� zC]�A6.�H��aʇ�DT'��=}���R\G��O�l��g�P.�f�>
`+<_�2���`�!��b�V�{=&�D����~������6��sԍ��[Ă����A�V��b���e�m�"!�m�B*�^�2�N0f�Xv1�pA�kf^�զe�mZcsV�`���v�IB�\n{��˽sAƅX|�
B[�8��aw���Ԗ3c���饰��@�����,i�o�W�!��V4�[��M�ͺ�<�J[8�����?�ϝF�P��ΰ-5��JMWf��cu�R���"����{�j��5%�n���x����t�P�ꌚ`��es�F����$?�g�!���{�N ��,jչ���gS�V5!G���/EmF怠|he;�GNFŜ��u�c���J��Go�}J�ꎷ�7��7R#���%��U2�%*�*�Ro�{=yN�^+[�g��*��Od,I��(Y���F;�'��{v��'BR����*����ʱx��c��|�'y�@��=�y0��q�&jʶ+�W�}�䍧؋-��u�m]>YXh�io{KT\\X���qg������°���b%�_�Sܖ�L�Y�[���;l�9v�G�"0���ܶ�ϡv�G���_���I�h4V��M!�fs�/΅\ �?�}O��M��vu�1�j��i�����n�)55�����m�����b�e�[�����pY�3�m5� dߝ9��L��ͭ�>QypTE�
����c��#�V��:��͛-�i}��_������;�U�l�ޖ)3��[�,�U��B:�k=��|�lt�!�#ÃGU��΁ 6��Qd��+�!'kl8X;nu������#ϑ�/��R��m����=SV͒�?I��Ѫ?CZ��I;�Z�(����("��&j����#4��D��Ϝ��AG1 �a1\� �R�·��ΐ��@#��>[=�fMxm7�]���V�`RC����@Z���ð���:������y��Ѽnaa2��!+'��WF��[ �YL׺
O��a�0����+�
����g�׵m�iw���}���#e�]I)>n�F�#��t�SA��E��[��nl���Uhf�E�R���]�Y�K&�C܃�t,�?i� ��|���c���#&f�~�+7���=��ۿ ��>����k�t�����t��1YMLL��.���	|PMH��${���90	kc��[���1]#�){S��� �T]l;�47.ddg[��m�ij��a���޶t��P?d0�P8{���"o{OO�!+GK�p�Xci��t�DΫ��qPO&,�}033spyA�g�!�6�����M����uu��1�jZ&k�݉u�yg�Is� ĕ�R��Wn�/���Yw9��{�K{Vt�y7��i��j��>����S�܁��$>1�;��<��~[`7��a0�6������k,����TX����v�^1Ѯh��.�c�~�!B;��;V���ح�K����ݬ$h����);�	d/�_uwv�Y�KD��R�J�jk[��iRvY�Zuu����RT��j�rD`�v����_��a������Z��m_�-�j�A��F��XA���f\�Lj+U��N�X�N�u�u�Vms�)�I�a�x ��K����g����U�Ɇ��6ʥpy8��| �]h��:f��}복L����t���h�֗�Xmg��{*+�]�?�͟ogwZ���Wv�Q�ڡ���5�x�"]�l�x�r�]��""�\���b��Z�Kc�xQ�>�z4���}LÀ���m8+j72�vv�|�%�;b�G��ɜW�e�@�Q;��x�}���6���PyЬ�V�/O?�o{�}w�32�Pp֫"�3��_�^�i�I�}h+$X�)"5�����|fְ����:aYu���<�=�]���rַ	D"4��*���s��{:��D6�VD�q�ߜ���I	,c�|��X<7^%}B�݌~�оfc�o���J��L٘2ˡ<�E>�Ӫ;O4S>�2���n_�=����R=q�dザޖ?�ǃ��7Gև��X�H�擹ϧ���`)�]�fs��#���d��7����Τ]/E�~�w6�}���Hp�"&�*{�&n���U�7���,XV)}$����ۂ8Yt�:۵�9z(����?8���z��~�$-��k6�a�0ʎfՁ
���X6����M�wI���]�R��D�R�W�����ITQG�|W|��� bc�Үv;�[�
:r�g7��%�@�ocZ����3q��?�M�GX��w�wcZ�~R�0�n�R��O�T��\3�&��Iy"^��^2��wݹ���$�?��>>���p��r�⣣�y���q�v�/t�={��y/�����U�A�"��׋U�@I�jY�B�x�����]�U�(�us	Q1��������BLz�vQ��m"�ǔ��!��2��}� Ҏ��ͽ/��ՃIHVꏢ��U㥭�l(]�b�>�`G9����PS5�V\�U[�Aw�ȾR�դ|�l��~ΙZw�`��纠��n�g�F5�8�	=l����6|f6?a>R·��Q���g<�,@�l��"\T��!kl�yV�P� ԋ��k�5A�r�8���6��m-�hl����oT�DEG���	�0Ob�?���j���n2��ٛ�D���X��SQp�~

*s?��Y�8�`��x�ⲉċo�o�	�&D&ю��]�e1M�V�x�e���6Z�����v�l
[4��S�,�	l����������`�����n��j6��P:9��Do�?��{O(���ZT����h���S�j��i��<lDk��d�[�	�AF���i�3���N���6)�MO���9��\�bJ\���,�:�#&��Z}�v}�v�X'��1YW�2X��L}ݼndx]��iIX�.5 �;��#C^�*�5�TYZO���n��Z#:neA�Ѳn*^VU�pȀ������̌�D&nr���=�L"n=p��̾����>듛�y��%s�۸?�G�����B�>{�;�DN���`���iO�S�Fؚ���� )��{��c��nK99��
�̦rջ�@P�G�I+�h@
�z~,iC��T���1y�L>��(����9�չ�Պ��z��54H�#<8iq;x��޶u�<�狻8�S�2+c�֫y�1��W={���7�'��n�0��A\����~^EP侭{3�w�(P!y\�2����P�����n}�U���+N�{�}5+Y�klW����2�u+Q�}x�&����Qw��ٜ��;������;S���!!C��I��P������}��`�o��TU��k@��_d���>�;��Up�*Ga�n�q��T�3�m��*q<���|ox�m��� 0mʺ�/F)~k�`J@
��%�L6{�yk��u����X�d�O�[�	/��5���<<��
��_�#"Ҥ�>z��aˆ�����z.���ʗ/)��\�:7�l\�ׯӲ�bŪ���C(󑼊�nT6 �)J���C�e;�a�|���i�˳�w�)[|���S=���Y;�q;sݗ	W�G:!/{IV�ҏ?��<u_%�A*�վ�@pY�/IIE d�<~��,EZVv`0W5��Wc��F�2�>105'.� �u(��ϣ�t���$���5PNϻi|*o�ݭ���і���l���ߜU2:W4�:�LMvo:S��_���E�57����?���P��M���y_��ooo@1߸5L���Nܮ;oZ~�׻aX�����lW�
��'�M�h��\���������pa�l�\\tQ�Kn5�ˈ�,`Ȏ�!���ޗ�HHI1��������$FCz�*�Y��4�k�k�φ�߉��U���|<�|�v9���<�
����֎��,D�Hs�t�G&�ل��)������.��gk�c���O����^��R[ߦ�(s�9���2� o���Ƭܯf����6�l�eQ�=�ieN=��4cccn�K �X ���$!��$w|J�2���/���JԭF��FT�2#oIKM=�|�e����o���7��kQ�[w��7��?��%!����ǅn�F"FfR���$��sWdT�9�#������I�Ո���Y���*X���/�Źa���VCyQY
�y�?��ڣ���`�m+5��oyV#Eq\���A��B����5���4�:���UQ\ ��d����V��������t�xU�ƾ�t�����d�W��3)�*�Q7�r�Vk��}E�#��t�Z�R�ja4B�����[1�>(�a�#= U�B��m�O�����OA H����&�g��`�{���
�o�2)���	/�/>�H-����:��������n~�
ܹ�J�����8/�۶�5;��-* 3Y����0��2��@��Q���[δɎ���t�\\#x�9�U�qS��P�M�J���{�a�OK�K�/� ��jeee��]���XN0��ֿ�ܧ���2�a=0UT�w��R��E�����꫅]מ-������G���nM�|6M2��e?j����f�N���b�l���O�b��$����N�1�&��4�V4��D0��)~n��ԩ��R�i�R$s6Ai`>�ZQ@H硦檦��Kx��DD��^^���fc�
���:N=B�/��m��$~eq����w8=���`N�k�Ϡ�yKK=d�WG*���'O�Kk��Cβo��G%ŧ�P�D�A���d������o7�ф�t��7� =�<��w	(����4��ǲ���%��u�M���gǛ%�y6_�&,aD47V�~�J�C�>x��E?f)&�+�9��f���rv���v�Q�x�Bph�0}� ����IB�{���Ķ�25�������=�,8�(������-�����ݛd����h{�$_b�Ӳ��s�4*
.?4_�A��~���w�;��QuQ]���ܯ�Sl��X;E�T�ׁ�ϙ�m�#�lر��5_U�0�:ԁd}��u��`Q�O!!�1lz�M�~�{�py;��8A������E@`b����0L@Z���+/�㱘���|r���h��3i��!>�Ob���p��%Q�J��Ȩ��IH�X���~�<���g��	r|�<�k�0-��,�����r��Q>�p�t�>5m����s�"N (P�C]M9J��{��OVl��<�0#�Jҋg°X��z�V�?����˭�ߴ��
�\�`��?���'�)9��z��jC��5��fp�(����V�:�xĠ �$�xJ4��j&̅G�_b�tУ5<�?>K$֩i�5��v~���*�{*���`�{�~mvuz�KaӠ�4���6/c~�oPQAJA?TƁ�2VN���Y�n�^��@���ݡm�L�f0R��ZW�����|>F� S`�V��QfU�&�Y�`���H(i��ܧ	��tu���{���W�免2���mh�,Z���5u����O�D��i����&,}MS/;xi#[хκ��(�<JBV�y13R��û�`��Wנ��/�˓�6�͒=M�_
҄�����+7���~�b�ɢQ q���\V�O֧�&  ��;���N�k�|�s'�>uh�t�c
fe�t#b�$y���8|AO�(�UR�֭ڠ oI-p�5�ΎR��p���o�K���w	/?�����A�|M��}'x�0��D��:��:�]�]���ݝJ=,�m��
�X`6W�)� �M��^_��x�M<�����"�[?jΏрJW���zaqq�p{�M~6�Ǣ}�s#�;_l
��)V�7z�MJi�c�"��C2�j�5���z�^��ZWȵ[W&���:<�>�ޥ�i��f��k6HdaR-��3�d���H��(#m��q/:��s�.Vq�Z�y�߉��Ⱦ�FX��������5�yZ�H8�HMZ��BZ[0 ���hˍ�j�w[)`@����3g�Y�k�ي�`R��DD��_��3�n���j�+F���2���I�S.6���d�u*G���f7t]b�p\c���|}PS�����A�,�n����B�{3�/*���?���k-��q�Z���j�U]?�O�^1ꖬ����� $^��T���k�����wu����3Y]_�H9�e�ʭ۸��d$p"�e>�ƍj����MX8WG���AІ��`��y?�_��ɉ����
��1<d�y�BGI��-��7�=��L��W \%
���'�_��HT�zK|ށ"{�8�3?����7Gm��BΨ[���MyTL��,�����3DiW{:
���=$[7y䈱���uv�ܘHtU�4���q�ٟ�C�T����x-qIMɨ{���;�A�Q��\9A;Rܥ�+�jH�QOQ#�n�g���/�7���gi��g\�'�Zz��ӏ��F�P�G����������~bE�T1c6;}�����+�OF��͈Ř�P�����@8Q����o�پ�n�ٯ�aX�������~�d���ĆYu���G�b�v�F0Q��9�����B�]��跇P��Q�,��Y�A���
����]g��lbꚦ>/|�phRzE���]�0���R�)wϊ�s��a�����0��#�	Oe�����J���r���-��Z��K���?�;2�E�(�J�p�(����y}����zFޭ�\جR��T�!/���)?b��w�!���q##ɶ��1 #hf����X���y1�=9�+��\y{{�%�=�ΘY��Jf^QQ�6����V�j]�<���f����	�P�͡���hK�aŪ[)�!�N�������G�:����Uߓ_�3MPx���a����EE� \ґ����Z� �U�v˺�"�*��xU���	-;�ɨ�1��#R�="O�7��b/��2�� L~��S�!�;�?C��}m;7J-�g���~����z !��۷%s#k3��bj>�Ҥު+��Ĭ���^5�\qʓ
�9>F#��Mj�~Ar������灹f�2�L���� ���_���fH��P蘒���J"�5V����-�����Ȗ!��Rg&G��YNj��������\\.?��d>��qڕ��`F)���[�g�h�,���I��>{�^���̓<�/ I�;%���--/?$N(��J��WD����v~K���fƭ'T���E�v0��^I_�m�/�l�סQ%o����õ��j��F�>]P�f�T���z�	^��S}�oSR�X��] �7FPե����^�2$�޸��(�ïL���˘�;pXxaq�@�3$��5x��_찯���3��\�|��e�r����?����{!MWV�T����9��_�v���@_�#2 .���'a������qF&'�I�~�'##�@�،�i����v�e�z�3�T�9�U���,�����q-J@�.��h�7�47�u%�
 6�L����g������Ua�2�k�o���ԏ���4�ew`1R�B�k��D���r���O�Uh	�-b5R9]�V��8����k4�f��>������ݸq*A #�����{�*ƿ>o�������Q��Θ4��=�C�q�Z�m�.A�y���;U��dde�!�2Z�#򈃃c/��TL�⨇��Ҫ=�E�x�E��������ｙ�x�z-���]�����1�*o�%.B��Eކ���V�X������b
ܶ0�D~���J������޵���-�� OA����zP�[J�ْ���U��s>�t\j5Ť>��Q�NgP��C��oN�KJJ(� �v����) 0l���(Xqw�+�cG��:����D������qhhD'�.�����WL��	��M�%�.JA�n������:7L?��ᆱL^D����/��h�$^��ݍ��;������5MLM�99U�)yY��i�1l�"������Or���?�~�A(>Y�L^�:�2�Nȅ����C7��1�PQ����("R �:�tKǐ��t#��]H# 
H3����- ��C:t�������k�֕����g�O�g�3a��5��$ tA���K�:bS=�,(`i<������UX�+����B��yԒ�\�,�+��Z���RB��{�:[��8r��k��Ltӓ�fЉws���~ܽ5+�w����.G�"��
���S`���=����!,��������wɱ!�c�lf��%�lO���]"����,,�!/��ňoLUۥ��'�iK�ٵaxg��P�ܸL��II�BɅ�����^J�v$��6xl"�BR�1f�\��;�T�9�����{�P��t-�Ẳ����u@L��N��R�����������$Qي�m" z>��ꨴ_z����yj[<\�d&|���c�ewA�.��4�����]OM-�*��)�}�E۩@ǰ{��>~��0��zq[}+H�jzW/��K�mciz�H�>/OX����B����.�Q|�՟�{����2�h��Bh���̄M���%5�l3���Vϙ������e-��#((l{�cΛ��:�?�,8�  �Y���E.8�A-���y�D�%K���:r�q��	�8k�>�p~�A|�}_!���u��C쪧{2 X��}@-�@K۞=q�"����*�l�����z��
��'G�$����XXX�|>V�×��4HQx����g�]����/��xq`61��4zc��0P�&ffV=ь�w�'̧+r/�(��A��k���݇�2��e�5;Eiw�J�N|p_^�@^u-��q��ٟՔdx�J��_�)��Zj�>� vsPV�����,���c`{��
�x@�OR�׻1���z��ey���#eeepl��e\oP�g�l����f�~��oKQ�Q\�����~{>z:���c�B6x�
f��3{B0y��h�B�x�%w��&p[���]������m�?Zmg���u�-
�wHG*����NH�8������	�&���:�A�s�/c���SuJ�[������5��ߢ�f
^���Dؘ[�IĀC�?�n���x�'�β-�جI+m��x�l���Z���Ar�����b}odt4i���ܛ���Nd[���x��$p��8�yX���0�+S1�Ǹ��Q��p�����v�ux�������++��	�A3Jk�	�,5r���s���[g�нS_�TY�V�unt:ڹ��F&���UC9�i\b�jט�uc�Cs��t'�h���t����d�>e%W�U�
mf�����`�9K��4�\i��x����� H�M����&��mN�M'��x�V_��p�y�Ri�ꨨ����X�Y,�_{���B�j�����yp�@�q�U������'|�Oh;�oU軘��ٚ���|�!���<��3H��c���
˷{<c1|Q.��k>$�Q~��fW�(����-�c;;�ң���������k�֫�f ��2��@����:���0��fi'��8i������-0K��w�>���
�pWI�<�-9H���l>I��T�ǻ�^Ui�6��.Ͻ�{$g�G)۫b��%�����Md~�����Ұ�.���,�ZMG �k�]n��[Ol�#�\�r X��r����,d1r0�~1=("g0�^ޔJ�nF�E1��ݺ�ׁ,*�S������#�k1G���1(��wF���UXO�Dcu�'��">�2����@>�/�%F�P��у���
��8�hߕa����{�~1��YGiۅ������s	dOdO\(����K�݃<������ۘr��=(����1�q��@�2˙��<��j��yV?�.A�>���c���	����#��R@�ׯ���$�%��֞���i��D�M�e<c ��W��s)�kڐ;��3<j�7o�B�hwTr�h(������5y��?��%���Xs^��;*�qY��UH�x~�shh�;9����/����?�zl [lэ?����ibb��2�8�� ��z��M�`��}\�O3����?+j�O\�z�g�C�_���JPPHJe�H��Z�뉇�I���I,�@�*y���R�j`�H#�+�+f)��5޸a��'�@x������+*�{'jNWq��Ӽ}`w�L�3�-:�=�R߾�����U[�4(`�� #����c�v����~�H@}۶d&m���U�H�պ"�ۢD,�W?����W��dv�ݙ��5�>�����W�"�u����5Re���� ���WFj/�D�X)���GY��8�Yj$�;q��g������A]����V�L�r���t�����j�������3"�o�w��{�t��҈QF�K�G��ܰ�QZ�֖���S��5����$�Ѭ�80�7�\��?uڞ� ���'�F����ð�����匭&E��Z�1�9o{�~Qz�w��C�7@;i��xo(�v1�`������S��\O?a��4z\��4���T7�K�	���Ϫ=�����"�K��o�V�#�8���i�O�Ԛ�EGiR=��!!P�]���~y��X�	����?�ʴl��?�}1Co6[q�z¨�&���aD�:�C���B��ɱ�PĸC�T�'��p9��Cl��%5��(O�Fh̑�=D��C��|	
��9:����۰�����ez���H�ד��ڵ���*�B�F�YjȯX�c�k"�WBJ$U�������'6M����?����b�aQ{������`
���A��X�N3r��,��(�����m��$�id6Y���T&{��l��AF�`#���e�F\�R#{ňu�='�\&:X�@y������A�~�����o����$j��R99z��hh C�����I�u�gh��B+�c��}*{8�&������6&�$�I@1[OU�C�an� f~�e)��%��G�����6����}z�T�	f��k�ғ���CFg�Q~.)���.peM�3C����x"vll�l�O�巃A�=�_��~M(]usë\5�No���ڭ?�7����p��˜<���$Ә��_}�E�N[L���Q��V���ӳ���5D�,=�Q��+t�,�� �)�Լ�v�p��*�ӫ�`��ZS��Q9rvC_0hn��ԩ᭱�@@��Y`-�U�7Fٶמ��^�I�c�����k�o�W˪��Og@-��fu�]j��F#03շ�R�����:n+�Nx�Z���<�r7��f��`�u�w<�SJ�_������/xrB���@�����G̤�!w�%�z1D&2ƒ����a������:�n㑷wIbu�fh��nx�-��U�7��D���\�ނ	���?�y|��K>��
%{�5a�O�)mi���>�,dlluf���ǃ�6hc��?�Ŷ��*��43H��V�<Q�*�*��N���Ux���|�?m�5�j�*���&�Tvy�GTX~b6ʪ�wu�s������Y�oףM���o�E!Z��:�:�*k�����sX ��1o�`���9��k��gK���~�#��ՓG���+_��'�?�]�p%rb���� OF��Fr@F� �

����Aaj��'��~>.�a�	��ɱ"���OetR���IH �h� �"J����/���om����h�e<Mя,=�RJJ9;�{2T~pRw�x�bھ��k�EgK���Ƨ"����ؽ�3N� (W�d�a�.:��� �c�ǹԼ�V�F�^�&g��-��k.��ŭ���\S'eP��6��3�j�9�(��@k=��@a��<���+̅~ضe��P�[���Mc��ˉ{4fL!p�Ь���X�@^�����B�n��q��SK�����DM_���@0$��G���N�:�p��MzH�DfP�#� x&���~���;[Ϩ4��p 'Y�PE*2�N@ނLv�#o���!n�c�V6��m`:�S�6�����
}S)�<=5�V�A5�@]���55�zr�Q��R߉q���z�E��u�u���
��۪���L�?A�X���[�H��G��wl��+f�ϲ��o�=�+���7�������ez�d<�HP�����b��_��>�^P'X,�$�]NJ��K�V�.
�s���n�Y�mŻ�tf�X����#f1��[��f�J͉!�ɽ��ȶΓ��m��dLP\_���7*����N�2ox�5��);ir�Kq�.��T��{Y6���xu�9MXj:��Y��d�����OGu�Vd�`wu*<���Dš��?̲%{N6��Ȏ��O�\�1BB�,��ʊ��TD ���L���?�ދ$������܏�p	����
K�!�����������
9�g'��aX��lq�5fb�����,�;L�/5E&{x�I�{SY����4l`\���u���cb�|�1���{�N����h�g�uma����/�wDg��r�>oQ�ѱs�U�-��m�@R��v�W��{fSއ��4�Vx��Y�B&뫗�gV.��
Q 5 ��J��׻Ϧ�}��?��g{0b�N��oژ��SG[(�E�K��K�J�B5�~�|�'�=;�ⲯ�D��U�#�+OM֥�(e� ��}񝳲j��"�i�;�]�hʅ>������ܻ�2�*��*�$&x��-؏���+ֈ4"��6Ď皠d�5����z 巟�S��Y�����Y�7FR��M0&��b?z���6�OuU�rit����2��'Zı^�L98{r���!��\x[���9|�@�wދ���Tz�Y�m\'���;R�nZ��{C���ƻ�0�`8ͳ�&�g�;5ǇaN�����_�׷��^V���P>(���A b$u	Ɨ)�X ��AF���&�fFG��Rb�Fy��O�
��g�ѝ�*��L���˲�6w6���p�K2G'�'��J�1S���Q�H�M_�y�^���襷�|~���s����CD��V�|�0��|h<
�_E*�S��9o��Cۀ5�����y��jk��AL\���'�a�����?y�[���&��O�S�UW2���_&(�jC~eS�M.2#ٖd�����n,�7�8�==�]>�$�O�I�Cw�i"u�����_�*$�aWH-w;L[� s�%��ю�ݰW�OCūf�E��{��eܸ�go�5Oan���T+y=w��7�m`��=�s	�>��j2��uy�;V����'�Y�O��PQv��#���e0�,	KN`�i�c���"Q�u�[�,k��q0kHXBb�<�Qe�X	)��dwm��n�s������M����J�'���0�}i��Gs0����a�cZ�Vh�/������C+��v@|�Ϣu䥔9cFz�;=�y�afg�"�۵F^����p�LP*�E2S}$�ş�S�R���3г6q����l�'�;�℩{��0�z�3zg_�<UG#���,�������>�U���?A�?��9i9�c}�7�� e6����p��	V���o���<;̸�Z�*fOi/��q,q]=��f��8o��:o����*1�d|�;�m9��_\�L�ܬ ���٩3�����{���@����
����WNkOS�z^Q��:
��6]fN*����n��W����ʖE0EvG���>��%���`�/�5��8H�U�KF/��;y�1[�X-�%ˬ�?�t#���|������	&��Z
`]{!����,"R�}k,��c�����ҧϹ�أn@��-�~b㷵���}�=ҩ���jl]��>�ٝ)s��w�s,_���D�����Bjii��7���m���Q��V���}R� U���P+�)b��(���yc���?�,���a��4�BU���,���OK�ݣO2��%��c-�BbNO��C�6K%��M�p�/���s9��+Ҧ(`�.r��e&�YZ�䕲�9�$VP+�aRM7����v>�v���}�.�:K�s��X)�8��Xp�7c�eխVş���SlH�������͸;;0�gh��k#�"Z=c#��'�T�ƽE2ǺF	M���4�W$C��Z�~��@4'9�k�Ė6��Q���o��]ђ�[u�2�.���B/�U��!B�{�J�-��S�K�a�zAg9�r�>)���<����WZo�j��
���+�CiL��-�O�@hҞn#����8�}y�1-E��a3���s�p��j&ev{%��x���S�}.nna׮�� ����b�4Ê�p�W��\���H�`%��Ȃ_������.}e�B�H�V�m#����e�z�4k��ީ&��|b�w�̅G܉��Q���u,�gcr9l<�4�+����5UZ���V���Ħ:�X�M7�'ceY��]:^\~�1���߷�z�Vƻ�E�[{5��̞��e��1OQz��xC �j	a��b�~�l�"�Md���8i��HH|ڸC�\Q �W�o��'\a@ ��W��n.}&�k�7�?p�T����u�m6.$ϯ` |.
壣�!\��D�2�hDғ�h׻l�L��[ϧ{�x��_n�&��zt�VU�y;|a��xl����̉�z�@@2{�8����Tn��|4�H�ۂkʀ��Ev:(!�m�!�'b��.ȓ�>4mФ!n&���h 
z-9�b1�RinZq�����ͧ6՟�/�;Xf9�Sw+Xi�Z-��Щ'�Zq��<rN>��m�!�O��hm�.v/�.�Bɤ�@H\�N�^��D8X�˕��#Mnc����T�WuL�^p� }�<��\����F�{7!}��W�yw�^��Y������S>��R1S����(Z�n�]�{Q�C��F1J}O8oA��M��Z�qB���o�<��G�CgbG������������;C���?B��I>��n�_�A�u%�r�T��ߵ�g��^�Z���%
b A�}2n�3my��*Z�&Zz��}�t��I�~xH�~݉>ˉ[$E�A�D!1�ɦc�T���x�-��jv6��ҾRA��\P܅vDa�ji�� ˜�lߏ��J�~��\%���{��㳦hi_�Y�<���q}�0����4���E݅Y ����g��Hu��L�R�ص��@޶�:�����q@�ܾPݗ�+�XS�H���'w?O�>&{���»Mȅ�����̅Z�V46�4{��oxۢ��,v9��zg�H��x�㝲����dֹyx��x�Z�=��s�(T;gk���{
�#���k3k�-u1nS���<\�}�J&8�w���,1P�.Z��kc����͓�:���A����<V��gk]tq�Yim��n@�>���e��!�Z"���7�% �����@*>������x�~ֶ��Gߍ�}��,o�8���F�[E�ە��[\f[;>��j=����;��#{Q�YY��S�W�P��Ivg����dQ��*���IN�_b��@;rR����f�)����!�,m��乲�g.��ҽ<���q3Y��D�ũ��, �p�3p�&�o�fo<fxoc�9�@k��\����AыK�1;�����ȧ��s���sJ�>��-z�����o1�W�)�%�k"�<�,X���Ք3��]K��tj��hi�ku��]�as.������èAˁ7���;Y*�s��:˦(euU��K�v�`�d�A�_1��@Ւ��?�~��=��0���`F�TnH��k���Ն$ c��GЃ�!`�48���)�9�U�`&7�W6��?c	8�>������	����,��UFA�عVw?�g�ȷ��/�D;j�dJߠ�f,+E���q]�����+��?���8A �)��zs�R�31�\ϙDw@�Ŷi���!�4UkG^���1�fU^i�t����/D�=L���r�s��_�	��V �p���	��0d7���D�^T�|�����"���KSl��z|�2����a�"`w��\�=��آ~�� �3g}�&f$^�ҷ�S���ImhY����wRB��8���&�&���|�������l�� H'�u�� ���Eؾ����l�k��i�N��ưND�s~��;�M����$�F�3wt��V=v����r��B6+�3�D�|�fY�=�<�z�tq��7PP֌7���X�^5��:^R313�K�y<QiOE���������/�,z��άi�\�@�Tqy�`�֞T*7�%";�]
M>�;�6t �|��5 ���S��{���6y�`/u7�����SK,;��뾒ܤ7/+(��{��?�Dҡ|��:/��J�B�:�,�
)��}�A��ol�F�d�T�����͠�K[�n+���qU���!�� B�mv�|iƶev���g������=���SFCd]�<	1OfPh����B��j�/o���¤ʭ�$�$k&UIb����m|Hl+ϟ�:2ŀ�]<1�-++�����Vw$�N��&��	�{����e�����2Jd~l�&��5�8�ym��]V��G�j:��\e5�? ;�+�U�3+��76��-�
�鳷��>3�|H�3 ��@ά���e�� �u���.�g��}�@	ܹ�E���c��Jn�j?�&W�I��uG9�|N^�d��:�'�-�s����3K��^����:i�찑n'�R���]�ugt|\2�fصT%	i�O��7����9s���a����� ��X=~?U�>�UIv{Hl|ؐ�Ns�$����D+��Qu49��_YH#d� �̙~��JEw]�-�\��3�w���^f�^�Q��5�YU�.71���;tSjH�� 4Jf(;���ao�pf�O�oK� �Z�Y���ѻYm����u�}�j��L��JJ�k1h�P�3�yy8�Ʊ^WK.�*�(wT�.4�x�N���XU����o��/#G��-a7�I�H>�����u�g�$1�䈴��#K;+>(5�x���&^�4�'��=�7 ]P~<y�X́1�$��C�O������i��mvCo�Rv�\ǒ}�X>�r�}�,��K�C��� G��	�4oI¾VW#i�h�;i�/6$^EG�Ayl̆z�4�{vf#CCt�;ב=e���t��,���&�ט���wȫ��&��;��죨��J ��F�9�%ݹ��][�p��R���>a����Ő��x�
 �"+@�7���?��_cl;�A�����J �((��z�vB�J�,.ug�'V�a�/h���/��_I�ț�Tr�Rh\]�0f~��ѝ[+`����Z�<l�uҔ��o���H"{ќP��%& S:�&��� i��ʲ/ҫ�+NGK���m��7�?���ǫ�Pͣ��|���>��{�,��'����I#���k��`�BsH.��0jHjϯs�[���Dɤ ���b��p�)���������p�]��(y�dj^���8^S풻�Ms�����G3�|���;J�8�vߍ�7�h�*���)�z����r �a�[����Ѯ%w�c~�E[�ץ.�M�0�)CRi��>	���^+��}���v��|��F��ZO���Rء�3`x�;0��ul͞�U�o�~��	���ů;��4���\KƔ"N�2r_��>�0����H��TC�o��'2b�*X��� �`O�^�,� ����;
��گ�{䥺��n\���X�^I�`A���Q�(�,�f)b�p�����H�ƌ�^�g�[\���uu3&⬕ŝ��7��~���z��g>2\��q29G4���g�6���2����2�+$J��KX�'Þ�[��m��7�
���������;�a�7U����g
�9-`2���˺F�}����	ӯ�VslqH�g�7�q�ˊ�+,<�y��4T=�J��^�E�O��$���]T�M&�O�*g��N��<�ip��L���d��[خ� �7]w-����e�ό�ʙ?���楨#����S�G����!��ÂU�!Rz]������� wDD<��y=R"�d�3��c�^'��՞B��)�S��F���ڥK��Mb�^�ǜ"�)��c=|{�ϕ��.����K_���0�ߑ���]���b��_��W��t�6�шꉭ�5RP���tuER!	�9�ۖJ`0 ��e&�*w$�&U�����"��J�"! }���겡88�-~DR�A�#���C�|�D�����q�/X&sdw��s�7h ��8�+�O�ł^��6ď{	L v(�3�6p{�P�6ƧEVZ������T|A����b�>�x�S$50��)�6^��e9��/����k�J��S�Cy�E���0��𤆣A�|8�m��M=��X#(ѹ&����хd�������خ�&m������E�>'7(�y+�SR���8�\n(6A I����SO��~�ų+�����G�!jo�@ n� �u��('{`d�V
����e�uv3�y�O�N����b��u�/a�Ⱥ��	(�*-�L*KKz� ��x� �H��8�.�=��HjKj�(5�Mq���a�\QϨ������Oܶ�Yu�f�$�L���R����M�/�	[/;_-�N)^uqѐ��d�w�T�Ł��];ȭ������y�_��ǖVV\��kt٘{Z��H���"_�M�y�އߨM(�"��y���?ڌiVt<voLpYWCq(}�w�۸��8y(���A��32�h)w���aЫD�Õ�V1rYr��*�r�B��P�g�]�7�!O:�X� �h@e~�G�`���o
��L�vrK�����e��y���H9a��Y�_�C�0�VE�^�����΂�W �W1�i ��N��^�G�x[5�
�ܐ֘D=6H���`s����$D���o �$����
���\�S��� �$�r������6&�����a�㿣(E^(v���V@T�-�^BA�?��.��))|7+�(���A�~�k%|y ���s���s0Y.�[�w�ڭ�RDZ��$k�E�X�0e�;z�f f�Z�?�EtX��G
�!���̌ڣ_5r�۸�ءE���@?@��`�7�R,A1�8��W�,600\���f��?����I+n襵42����p�Y�L�~����U�3��$V8x��Τe=u-��P�M��Gփ`4s�+(n!��Wo�3j��D%���ݑ��g���{�zmY���Z>(���+3�e�9�-=dF&&'#|t�A�u:1���}������!Ԕ������$/�6�*<4}bO4�6સUI���*K���VB�^b>ڸ�:�9;H�|\\A��h{�I� �0a�r���J�qDX�f���1� 8���mK# \������	ʕe�1��k�Qd���-��)
O����?���:�`���y��1}��E,�>���8}.(��_)����y��~9���h�krٓ C��?���n@��a��`���W33=�w��dǊ�k��4��P�o4�kտ^��a���	�-�=�a�j2Dخ�zW;�#g�O+��n��
����N#��������0�`�ѹf�T������B]�)$!Qgt~�H�?�5U�S�x�[�>�_�7۳��y���1�ѹ���4�����Ʌ�z1�W;"^�����^��'���$�M�����ݡ��}0�f	��־���%�q�p��nM����5����í^��GW�L;h����Lv�Ѓ��u��R���R>Q��V2�o�|m@/l��;�cԨ_|�`����m��o/�}���(Op;|ed�gKpAP��H�|�{H}�0�;�7����J��Ҭ�����G�?���bR���ARK��6�7��A`�A�5��彚����!�@$�O�]�4_QTX���h���6V7�~K��zM��l5a1�3�]��U��()/oJ�ޱ�`3]���k3>����֙�h|�A���ϲE�ܟv�YuB}�&$$v��#��K����P�]���$P���|�ڈtdO*{���??IP���N��ۧ����Լ��$S�Q�N^r�h�!�!�#[�V���ʫ�S�����w&,��ːG��x�sIm�\f�׼E�l��Ɯ��ęO�I:�E��y��-��ӺZX������oM��F�m�c��_�,h.ӇE�q=e����T�0�W��(F���WW-n��sz���,��:��C��x���
PH��P�+�T������+�7�����O��K���7u���,O�d��_|���-�Ӂ@�9��A��RnB.�g̿�XK���&!����2�1EOEr�X���&�D�zn�zoc�.&&�ؼO���z�=w��̆
�i��ih��ޙ�ʐ��4R?ٴX9(/��T�a}�ɷ֜%��h�Y��Uy�p>��ߏ9�!�����]�fb�:?M�]�W����xj��(>���40d 1ک��)J4����,7����Z�CX�6�Cq�C|�AF��%���������ah�L"O]�idHa�v��V}}�~[Z��hBt_U/ꁡ��N�)')nK��1�O[G'F&Q�b����9�(�j:~�I����(�܋�ݲ�浗�I�E �)�(�x�&���iZ�s١���f��Ml,��5��,&��4t�;�p�O�/��ls����O{�0�����f���9���:��A�Bs���(|��/I^t���U�[�W�镣"�)�z9)g��>Z���4��x*%�2�@d�*/ɬM�\NN;t�Hw��)��L�1�� ��iu���|z�Yȷн�
�\���E�"IwF�Y��AH�\?5�A�rpD6�7�M�w;�!�򾖢8��:��O/���H7sV��o��:p^�g>��Q�aa�� x��u�B\��� ��ѿ��w��q�K*ɺ󺥑��2���oi�A���+� !�!�p����A�S�B���[��\�I��	�~OM��8�Sx�6���xc�'H��V8��],���g��(l�;;)tDFΈ^���]�c�������mE�_}�=
ՠ�>���1�d�Q���P[3���h��߹ŠJ� v���y�;pժ���,Qn�2�wٞ�(_��l�S/w�8ϭQw��M�&��`q%�����,�����(怶�0�w�W�C�O�5y.vŝ�ɲsD�PE�p�������g�������a�d_��QWQI�%�8[�l�S᯦����'`h��{@���Z����O���7\@�\�A�I$볘�-^(��
#
׷U}.?[ApY-٥#w�<[�7��A���Y�>�Y�_X(!�d�꣘X��X��x������^E)�5��4xN1��0_N�T_�|b���긠6�c�u����O�%�z���n7ڨ7�z�
�E66ɖգ���Z������8�n���a�l���1\���s�u�E��%��@�?���x#v?G�}(x�"Ȓý֕U$���HWnOL���	��UV��1���6���;����v�}�cK��3k���!��j�1W�h=~9l������" ���FK����� ���Qi	:��[�9�%�����X2&���d�3�1~u-�#���Z��@H�=�u��[�Z3GH'�EM�ګS?BX1�������2Ł�������~��}V��PI>ǰ
֔�'�����'���J�[�.��xc��QF���0U�i��U�=��-'�y��k�z��\�߈DrR����w���o-�[�ֈ4]JbkD7��	`�+-P�s�'>�gdI�4k�&�yc��a<���q�_"^�S��Y���Q�{QA�1 ί����Ț�ONUB��@��Q w[�>��6 �I>�M�|�b*���Y��O�v"�2��;`\tTӿ'�f[ke�|��?�x�!\�5��cӋq`��: �;�Rf���s�����	��m�}ŉ�]���M��v0";�d�-+㬝�EqД�P�.B�)F�ã~�qWid$ѵ�������]7Ko)�.����G� )8�)�ܮ�Vey��Z��&l��}�����A xa���_����#�J��h�cT�+v���T��:g�U�άm�u4� MzLE�>�o7dS=��v���ҹn�Q��`�!��؟��N3��^?/y�s2>����?�f���o{������"+���`GWCH/Fj�����r���N�vwι�Q��۟����
��z���������m�L׿Rx[VV��a7���<���0������F$�����&FF���GDY�ܛ�`�Iq�'�z�r�ļ,�� @�j��zL\��,�����f�Bc���/.j����ð b��e	S-9�tP����K�����m9�Hgff��lk��ʶ���3V�^�w�ns����I6���bAE�Ǯ��ζq�%E(Fj�x�{��13xBohB�2�mXY�;
.,�ib�.M��'GCI<ZW�A�O��<|������n6,���:�:�ʵ[�}��y�c���Ob���e��z��w���N�E���.ϧ�^��� ��%g41��ūH�L9���*�[K����M����Z��
����NF�r����п�|�6��E'@K}{��<A�iz��|ʼU�m�Z��	%V����7<��M�/�W.�{*"����;[��T�� ¹���7�E�����T��;$�v�䗡��	l�c��~�%Bz�nb!��i���w?�5MQ<~���*�̎rV��N�2o��#��f�T�妦�jͽ�Bf,^�d-�OO�P{/��k��15l%�3^p����4$�mɍlx'��÷�.�O�I��8��5olll`�?��:o@(w�D��oͯ�|�����7��f��1X��;��CV���)x
[	9�[�nb�_�U��#V��E�d��0'9��q�"�`u���s�b/7���<*�b��S��O0]u�E��o�?�hͨ�)>�n[=�p����7��k�B�� �,�<p���Wc�it�+V�̍R���S+���F�{JDb�wu��V'��ӓ��@���$W��c���D�̞�ӉJ�`�ҩ!b� ׭�m�G�����擗��#V������f�Z։=:�&��W��i�xV�3��H,f?+�d6$|�N֊���D���FR>U��|Jh���͜�\���p%���K���A�p����6h��n�>��Vw���=��r{�����Yktp0��>R7�IV��Ӛr&��{A�Heig�ł�&՟xu4T��.�?��L�T褐�!����v-�n���u�����k�,dU�4�L�(MΏ��Ԩ�QgR��Ǖ_B���0�$�l�P���
(C�e ٝy�2�\��ŏR<����I���S�QW	�8'�d(�hi��&l�~KF������1�Sg��n��7���t�RϤf{��B�P�f�ٶ����i#K\W�9�_epы��^�a?N�cxݽBWY�Ǧ�$� ��/7Ja��6�5��&�)%T�*A������rA�$�]�S=�'�OT����Ky7/�	V9 ���# P�����[���Tg4��� ���!b
n�l근��'6�jԵ��/�dE�,B�U�:�d�*��!^�V6w]RK��3�!��g<�����;y�'�g.���}�o��3tO�qW�Wd0��xLWr`��m[�:����A����������p�;L��x��]zRQ�|���p�������TFyyy$5�Z�I�`bP�}8˨
���9��9�nH0���j��F.P�b�S��`Ӈ�d?X_�m���c�cL�q�6�7���ؐ�ɓ!������ٕ:]q�����R���<Z��'�l<Z�f���+3#K?�����Hy�tR>�L��m�#�^�7Q>��s�D��O��|Jl,�-ڎ5l&��y����˥��(Ѝ�*�2�M�VU��%���9M~P��brf�ᚭ�o��uM���$�J-�\��/��I%��;����F��_�gZO��s�&���Zi�.�߸�j)��9���&$X�C���D�5U�=P���9�/
"3 �F^�8��J��ۚii�=�v��8k8��E�)�/y]���[���T��	�j����jn�|�2��-��A���p'7ȿ��o��"��̞���0i����I�x]�`;�m�tv�f���Q���_g�`33�H�����dc�䴆��Љ]
��ߜ�Bjq^Gb(��Ǧ��EO�B�)��T�J�f�t�h��¿^^P���ڑ
��O�!3�ҿJ���n][D��ms}�H���-m �|��|��n������E�<ɯ��^<n��@�{��$p7��vA�y9���o	�f:�\ܞ6�?	��2ґc��Ԓ� -Z��͔Rl~p۵7�>�?=��aU��߹�&.�hE)u�ܻR��w��L�?��rݘs��0��*X
`!������DŔ�MvA�%](�A�pf:����%��[R��P��ޗƿ�������a�i#�&1.�D��a?Ǉ�=�Á|�N߬�?�zO,n���o��`>V���Kj���c��|��R���Ѝ,#�7O�cs�u�ew
�N�wTthlaT"��ed�8�vf4q�rb'�9������X8���"��z	������i�_[����J�����N�*	���b��X����S�����H�=���!��O�8�fp�PM�D$u�[|�K8W@����v�1<|�V�j�� +�Nb�o��z�''��υ��&@��暛�/p�y�wc��9�ѳ^�Z�u�o;����<٘j����mD�Re���[�Í�������/��?m=�^A\?ms�k+��v��ޣM����g�n�6j'�n��`�=�;�~E��]��탩�|p4��@";Vw�,Z��0��4��Fn]��W��n�����.\"��A��<P��4_&�괳h?iY^��W��vF���/=�l��s?��56���A"��#�`w+��ls��v.,�b���T).��᯸^��y��c\�U�F�pn��bag�-�=�	�۪Wz�JAM��'�4�yuu�>Z��������,�_M�����K�@?Q=&�Y.]�n.�Zb݀|��&�9�7��Ul(��(�~A�#*ut�}��/v�!g�v��|���%�q8�=���ՠ>��`l|��x�o[`��M�߇⁖#%L��H�|3��<G!����W�jxS�r���N��Z��3Y������c=?=��ܺ��������"�X3s����|
�q��+M�Q!��aA�MI��^����,7���էv(�:oѧ�7��?��*����F��Fi�����A@R�n����F:�[���k������_�,]:.���w^�����6^��q���-�ȓ�L���x[�O��rz˸��2�d?2���7~{�4a����?�΍�vM�{s:���,��638663Cy�.S��d��1�mQ]�޲��<U���T�4�A�q��7A��p ����D N�v+>�.��[9R���;d�(�cV<�Y��<�#iM��"/y�O
 K����J]O�`L��\��.���%��|"����~�]K��o;���OB( �R?�
Y&��'$G��H^��u�O񠓕=����I�Cw8a>�H^�_Wr���`��O���������!��=�L�l���1��W0}�d_ )�oH�(ts��ևN�1 Tm��M������~�T�Ԙcj3O�s�������麛銤P�m�i�d��o3i]D�\0����H��z�����_!$��f�1&�.�Mw�C��i��nA���ڑ�_�Z�S|6 ���XGh��&�ԪmA����t�9�s��rP�75�8�R��񈗧���z2�5�m6<��Eظ��j�A*b�=,�Y����UN���@�iX���n��q�U9���mG�o�6IEfϥ���8���8��d5n�Mk�du8�7�v�(���ܵo�%5���i��=#+��_�q����jh��7JOő�Acb�d�*s/�|X<�p�/��n��W�۝�?]��+~��z��~v�s��җ��~�S8c���A�zu�r�l�|xHT�
�f��d@����F�V��}�>��ϸ�_�-���K>B���iE@(�,��a���9�XN�����$F�&WT �ɻ�$)�j9nT*,fx���t�sz�m�i���B~w�����M$Q��%'I��v�E+�f(7��	K��N.���jW��_Mò���sM��n�C��l#� YW ڤ���W�ހ.���ܵ��&gF6�À/W����Q����bc��꙾�ك0��f?����� �j�^$�>�W<��,�s&���Ej3g�/$v��z�}$�y�Ű�H#ޅ'G�$�.�����[eX@�ߘ�۲�̘�+��;�I6�70t�����(� ��m ,6k���
�Tၹ�~!�|(���� �T
o��v�������j�-w��OQq?���g����%�W]Ŏ�p*W-���'�E }��K��#�F|H����z�q������)p}��to�����Q�VqC<o��"�=P�P�O*��C�,�|�t�c���\!\��@���k��p�q���q�1OM���w���o��b3�K�O�����5
�xpB�&8)V���nD�(��*�?f9ܹk�˜MJ���yJ��~M\S3i���njn��w^9?�>��E�L�-%��a'{@󇮬1�9���d�JR��j���+d�`zjΈfJp�f��Dnq�45"�=͎k�=�)�Mڼ�7��/V{���ϕ�6�ߜG(��>�-�g#�宍��������ЇP�ܮZ~Pz#t��OY����Aj�W�����wcG!P���X��ߺj4����-�g: OHݷ�&�>��/Lwy4�X�x�dZ��\��0�͙��R�b��x|?	�q�q�����=9b�<�ܑ�o��fR�W@W��xivQN1�h0�����N��.���	]\���>L�rr��|����Y�w�V��Qqt=T��\����'�N�""(O"��G�`Z ��%_������('T1�@5Gb�Ou��`�Χ������z�"_6���*H�O�����WH��#�����T �z�<'��Th0�OwqD����jt?3�z��V��ErC�+�s�:A�RBZe� ,u��F���4��ٓ�}�����(q����yKѻ���W�����/d/�4I�0H?1}~��}2}U��+Ǩ����t�K��RV ����4#�nK���#V.a������:4I�bv�2&��ݑ��;��Q~����u#���]l,,��6�$yDT�XX����L�]�Kqj�ވ�8��W�|���b=�ծ�9��JK!�h��RR�V�ϒ����G�
C&�o�3��j�y՞���@?@�h.�%�"h-����f���� y��n�K)G�_G��?��0�x�x�w�y�������aB���Kc94ߜ��T���ᆰ�c��k/�����;1��'�]=[K����M��F|�j7�58���2Č7|��sF��^��K��1�Y�-J�w��E|�n2XS�n7KV\l?!��=_�F���F���ʟ��j���2���I�L\�a�����'05�0N��˛�]���f���¢߼�������<���NQ �R*�ǭl�Lι_r���;}Y^��}U�i��q,2������%d`,E���:�m�(�{]0-�1��G��a�'E{�TC�4K���fۘ���Y���࠾E�g��#�-���ŕ޺��s����� ������Jҙ5[��)/���߯<�k;U�.%L�<�}��L��o��0���#����
_懩X$Q+�Μ��&�����F,q�1��(���6�o���YSyyYֿW���y<�F1���*�eZ?1��pgo�$ ��g��G�o�Q����籂����j�V�?v�Ȱ���
����M�}�R�������ßIs+�N>��?��4e�0G���}��C�F��qLDI�O����&1�sF��I�?��~
O�)�wL�+�y���Q�2���Y�phZX9>��Jg}�|�`���P���7p߃��νؑ���R��V5��屑�J>?�����X揟Q��$ỻ%�}��O�h��6��|On"�����x��(aE�*�2�	َ4	�<�XcY{����x�{A����t�e�N=j��Ň���IL�ͣI|�*sz�\펡C�s"zq�ý��|%�|y��~^���}ɟ9ř���_SRR˖5���m��TR�3��IK��ҵ�k�ѧ�����.�x��`��ƾQ^w�{AF��]�y0�*�F��~1h��j���dQ���>�������C{Y漏��v����f�(���2zS�2����:��'=M�M��t��3�/l��X��q��r��\ �_�D)bAg���=�q�@xCs�#a�{�v���_AA�b�Hq,���m����E�^r�-������D��y� �_)�k?��u��s�%�=d�픜6;����>���o��{�<.g��>*�mcJ��.���w~�ttI��5#^����sn���Fؠ@�IN����yE��&v?�k����tէ���C�=h���f�S���<����0��4i"���,�R��e�Y�}{�&�� �9�J�f[s���灯HF���O�kr߯� ���K~;u�P�R���^G�`A�l-~(��22�%i؄0�\�f�K^\|����-�34X�2N:S��GA����V�ߗ���ْ��jV�u����Ӕ��,4��ru��E��=o4��_Փm,p�]��{,�z>L��p�)3
BFJ�S�m�9P��)��Qq����2�T�o/�{u��ܒW�� Hz�B`�vh���M�Q����SYָ�h$M�_8��(?Mq�l�����}_�jFz<��?3�њ奚�j�ʒ7t�rR��I�Q999��"D?L�&Ml�W�IZO~�X�w̮�Tj����� JD���\䫕8�:͋mw#)r5��I�i��d,�����?Xiƽ��i3���m��|G8�e�M��������+�aE�PA!H(���ko��ޞ-�l�ޮ�~�R���sr�4�;�Y�wo����|v*�l~��PT|�&Ud nDig�q�{�1�
�R�h��6�	�`�R�z��6����r��ܥ1�Fln�
�	��ң,A��%c�$=�$�ޏ��B�<Nsㄒ��L�;4uמm{�Q�hF�)����h��$�)�d�;��q�!�j����~TJ�0@A��
O�|�v��c��V�=�Y�0b\k�1��*ϥ5B�h���-.8�;n�x�z����Ѩ��m�e�{�<��	/�񌇚��$��W��6�֋��fgW$9�ֳx?��2��Y_�*�rb�r0���.�ϾE�<Ŀ1�O1j �]�O[���U��ip^�֞����F7}���H
�](	p��H�$S�K���v�����U�2�ù��0V��T�i�"�UK�.VK�tkL��O��j�j0_�WV�I��w��I(w�,��1
�*��EICw�y�Y��]'�R����!Up9��ay�5�[�a�/OG�ֲ�`R.A/w7�UU�.6�!/���>eǔ�F��Y)���k��������-�0I*�^�vJ̆H	��`���I� ��w`��F�y.�������UʀQ�9R�{D�j�ڄ�^c2�B�\[�e�����-���UK^��
�E�q,�$���r�����Wb0�Z��'�[����i�����6�� 	��PR߶��	/�FK�����M)�vq�[����پ�������zŖ��r�a����1���o��#A ����Y_����Th��
�s~�!$D��/ ɂ�}C`tA͹�Z�<dr }ȧ�e?fJ���R�X�V�L{�o��-���.AU���:JV�<p\�+���F��Zr0:nvO����u����Ɩ#y��C�H�XoGe0��D�Pb�f~�ϳ�:�W�ٱ���,((�N�` Mg3��7�s�d�2b�<��P�	��IiD9 :��o��x���d��9qϳq�n���u3��D�ݤ�R���M����!ҝ�.$(q��W(i�[  D���*���^��0����� �X'&�C�4�d��.�*���`ij�u��֙���̊�����,O�����m��A�)����?���.�|�����ԋ�f�Z�(������A\��2��GKY䎚Z���Q4��0@�f
T��Q�
n߮����@\!e�����n1�s���H�����s'��h�1�Y��@����I��ǂ!��%�r�BD����j�]k��6��J�殘`-�n�J��N;�ݍ�n��&{i�M54�>[H�U2����f����3)a�?B����<�w%,�p��y2ֽT���>h���Թz�L��Nl�������{����T4�5tjji��-d��죳�|���A�gV���\(�1F�*Uk �� � ;���\�EmL�?uc�Z�C�������8@9���[��nK�k��Ic&�މ��@w�'db�F<�=m���r+$��-�hA/xD>�ŉf;m�2Dܮ�����v��>�i|ֲ��[�^�~;�l����H�y(�/���%�c��E�S������ejkP0�`�(P>�K������ɶ}NJ�xϚ����;��m0i�F��A��i�|�_���Lq�P L# �o�����o����إ�43ϯ��x^e��4�]4c*��Z�^�ڧ*;y��N�8c5�kq�v��~W=�0%�bT��v�����j�"�����	X������gy��uNB�W�a�7^�++3Q��.���%�[��傐j�t��������v�fLhi���#&�����`�%.M�:�.@�E�	����,�����k���*3�%]&�^ց^���#p�\�L
s��T����9���4�F���� מ���`�X8���m*38�q�e�#�CA�SF���r|q	�^%�MC�K ��N�zbaYFǋ��`�?",�RDk��E��`I�y�]��/{��$�������E㋦�C�@.N@o��/�th_�2��&-��k��]��
.;S��tU�h=a���F�@/ť�Iǖ��E" �&}�)��C ���j�M--cI|��w��P�(����N�ͧ9&��B`L^���nQFa=�|k����[��»@NL��u�l'���~WʓX�$�1�{W�ly�(��Ic
����@A�N��}9�`��?�oK������u��*�Woٰ��|��L�sk�]�*�Ἆ��ԩ���s*S	~�_���m)�w���U0�z�@��OcD�Y�Q�r�Bvm���ּ�f�{E��w�������L�Li��`��u�SJ4�����/�	JƝ�wG MP]V&,*����̪�XW퓌��Lᣬ}3�V^���ӻ�ךo����Rڴͬª�d�L֠������d~�>1v( ���XL��`>*{��n��j���{]ۻ�0�q��9�L�ǖJ�#9����~�q�Mw�L�����.#�W�%��͑�@=88X�u����Z�w��k�@h]��;����a��5�ΦZQ�]�#&Fm�y������,�������eDt�
��ʲ����	諁Z􇬥ٽ.��s�WɋL?I��2m7~��8��y�R�;�}���+���&4F�,�rJ?R�Ѭ�ш���c����bR?�r˹��9��6$d���4�w��O%+�6ݤS\��"P�Y!P����U��Sv7G�d��g%[eU�d[����+���o1;U�5q�����l�0�8������@����f����sٙ��5ũ�Ͳ� ���c�˳���9X&՚`Tm9�d��iĻV�͕j�r�=j��	$?�lREFo�eR�o��O�:�xq��b3�[[����'!��=+]�{�ݛ0/W8�'n� r .�M���9N5nRR�Pu�aV��=t�_:����&j6��#M�į��
�!�WM+c���3Y4��ՆT÷Wq�|s�#���PN�;��}<�Q�es~��7f�$��+�kÛ���h�R��f�~(E�(�˔�ZllY��F�'��>F�{ìc��z5G�?��ٞ"���_�v37�7��6������칰���c�^Z�(��6P(��x����=�R'>��(�ѷ�Mթ��\���2�B%��-����^9��-c�(t��z���˳r"W.�=M���5��
����ˤ�'WW�jL���ݦY���Z�AǕв^�𘲓�3_���������,q�u����������W�C�S��
�ȗ5m)���>�Q�������)1��11ہ�phf�QZ^x�9U���5P�o�i��=�'���1Q"G���Q\���FP�:L��~�3�����C���WyI��P�
é��?Ɍd����[X�����ٲ�U-���� �u�Ar�X8��אC�§3AՖ�v��E�ZI� Y蝇��da��Hx�j�ߓ�FG�BX�X$�3����J̆�<�Z�tI'����A߬�O�*y>��y��L���������EZ���N*��!�o���s+:����kH?`S=3s�Ͻ�jjYEE��XQ.vJ&�n!���36B��.ξ�x�>EJT��;濧�U?���$����k�[���F[���F��p��#�L�~�3�L+]��[ى�);�Ff�}��%�(%�6f�*{*���)��v�U��i(Ok��=�=I''�8�d*�\ �u�}n^��`NI_R�匟~�Y�-����>[.x�;H:Y�~��[�y�V�z���Ū{i;06��F��W��s���X n���w����U��&d���'TSS���c��/�-U�F��T����l��A�&�T���q�WRӊ�d�+��X�o���L����Ϩ��[��
HY���9��9�(1��z"�kᗬU�(�슙t[��~�	�-�R����y��[ -��D��5ߏ�b���i�r��>I�Z��f�j/�})� P�bj��S��5���B�V�a��ϵ]p�����bl�w6&$��}��E�[��#x\m����CV&������.g_��">��2�jW!ny�T��x���H���m��_��ſޢ���돦��`������#��'��A�jʝ��A5z�.�{KZ�I,�_<���ho��"*�5ٷ�ɬ�<ܐf��*T��L��[���5ٸ&�)fՄ������+�b�||��������Qܙ�B���`� T�"�h(��_y��+�դg���j]C�IVB�D�'%2�7�7Z�҉�ߵmr��ԊV���`��31��9���X鸯���J�o?�'*w!�\�}ꩩ�{5�;�x�~�����G��o��)
��@W�.�@��c��#>^����q��A�$��w14�H�[M��<�Кl�!�6�6}�;�sp6q�lR�0��;��D�6+J�k~�-+Zp-���Y
~|ߋ"����  d��,�>1���sqP����>��@Mb�b����F
0�g{�����ԅ�������W'�X�ړ���I�����!���if����'|��p��\���2����s���LB��3���*` CUՅ�$��<K�$ٯ�zjT!�#Ru��U��O�K��j�ٶן�Wp�Yv^wt;�ʓ!*������6�

\��r���k��0�Zi��)5Z`�/��������*NGA��Xs )����/݂��?�bs��t4m�B�d�{��%|�v�3J�(��Ѩ#�����A�qӜ��|���5��-��E��9v�`z�F�ѩ�����]���	����7��һm�C4��R��^x��HƱv��+����J��&K����>��J�BHWQ�E�їq�Z��j��D���b�cnM����1�$����6��$3%?�ƫB���h�����"�u�se���t���)����]$��X0���T���+j����5�&|T����.��(����"q��λJӑ��e��\-N������\֤c\��lKY�ǔ%}�o��Ԭt�Ӧ������'���_�W I8�s�ئ�^�9:]�8���ם��B��ȊP� �>�9����Q�ԟ B�d� �3�aA��q�"�|�ڭ��*�l!NĔ�1k���0�n[����c�"�OW��8&�2W���^:��V>��T�:�Ζ}3�`�GjTu�5uGY�mۦ��,�b���R�6R%%��妺T����B�|ǆos�������{�X���� ed��ݢ�U��17�<��m��y�����T��[����%*6�=���#���9���p�b8M��D�<�e����U{�Q��9�b/�7]��bȯ��-���^�G�W�zM�3	���[�� ��F�F$L�Ǖ�b����H�zj����������G�]nx�|kxg�r�]ʏ������gַX��$�z��ٚ���'���5No-�m�v�	N�m�{�W���^]�Р�v����̞��zVbw��Up�;kY�f]e*�IH�sNP����7�S<��eݑ����|s\�L�� ;����`,�	���X��۝��޾�2�B����dm�s�l�3�IU���� .�=��L��q�S��7�{�)������Q_�%hx_#f�̏Ǜ
�䳿���:�:t{e��Cm��<������xafE$�^7|�ձ[�p7}�8;��'����j���O�G�b��=9���vI^��d�4��8v��tW̷� <{��N�C�G )I y�����Și�������aI7�Pμm<�wOޮ_�â�Yo�ۚ8W��>]K"���:YWW��!����
�nd�����⸃�Ƴ��{�Z�J�m�T^�Oq�[G`�m<F�ĳ����]m�>�R

������hj9��	j՝(��߿����q��_L"�v7����Šva��u��mK�D-�Q܋�Ϩ];�����°���4jW�H�S�S�JaoV��:�I=��!��3^,�����z�Z����·���OR���U�>����6����a�=\p*V;����r>�a9���n��(����]�XJ��N���U�a���#�_@ r������P��%PqaYY0�����{˷2�\�..�����{��N�J����¢"%On�V0�ݯ6D���ܫ�/�����i��|k��$��G�����=0"J�oh�d��/qҽ*�Zj:t�#�WW�]�}VQ}+Y\�`��p�K�n�f�ƚtA&\)�,�����Gy��́�����s~��]�\����AQN���$���iE�����5Ƕ� O�M+�8l&��:}���g�V?�?�ZZ.9H�Q����Q�y> ���U���#�8>�Aw^��q�pͼeqB�4s�F�<�#@X���Ϯ����ib�b������%j��4mi�:�vO/Fs���o�F2D"�,f
�xw��� �(�{ƈj��V֕�T��<��_n>�Y�J���My�!S����
g!����h vs���T^��aLW����ƚ���^�[Xd�t�4� �2USr�w%#o�Z������sK=^���1s��>ā��&x�*�nd��s�	���F��%lv�ǆ�Hî�kJz{����bp�9��GE���I���(z���"��^: ##W�O�F�����ǧq|hs��@w˟�}�OX�
�M��3Wt��0���|�Y�<%jk}f����:����lq�N�c J����)b��
?_�/����x�FH�����]���+��J"ILD՘P����`q�+�J�8�5�x�5H�oۍ������L�a"OD�I"�b�#�D6���n����N�'�I@ϫ�J_��*����
D��hڊ�o!�x?9E�j�S�	9L�NUvdZ���_��B�S�����L��><�eV!CJ�j?YZ2.��B����$��(&��ݻ�_��egSN�����~�/M����cPˬ�?撧��	'B�gX1���% ��]ު�l�����(�\�a�["��Ύ����?o��\�����==}P��TT��ɸ2�fk��OzN�7��Ȣ�����>��M'q|���S�.ʐ���ŕ�.����� 01��//!�^��:��/��E��`�I���*2���V��jp:������g��$"*"[uZm���+�{���n\{��=I�s��6�&1l#ED�&�w�w?�}�߰6�t��'�D��O0 ���Db\����E«�?�Vd����&�1�n2�'�7��|*�-�C+b��tKD,��g�.�OTG��-�����ݮF�W�59�8|r66��\M�}}��?V)ޏg��������t���'L9��"I��X�cb���Kʁ�&�WUWG%$,�_����������.�t���D �(+��/=��h����2�&L�p����k�����+7Ǔ��� �����S���0H��NU`>=Yq*��x�r��#�����B�����n�ؐˡD6�j���łۅ��R��
ɺg�)���Zt"ccq/g1����""�gf���7.�'y]N�A��O�AA0?�1�𧮲�������ۚ���9��;�/l�]z�##�0��#�{/�"\�&'){�>]����������6E����`�d:�h��?ѵ�_o'����?�؞��B�,�>��G������6�]�ķ�&�Q��28���t�������!��ς�K(�Ś$�sr�(��=�e?��$1�=`����~��W����!�&��w��k<���%�2�@#ڙ�_���
�<���p�Xg8[�M�lܱL�b��I�K��1S�x��IK�6X�����&#���f�� BA��]
74t��Bl�[�u�����t��w)ij���vGҀK��ͻ�O�����Y��___wي�Ұ��@�y��N�ޙ?M�ō��[Pn�{	��Q��)�&a�l��b
0�Qh�0??���Ҋ�RNN\��(Gs����� ��b��!@DD�]%Ds[���M�	�	QNN�'�\Oq0��6�D�{��߫B�L�����s�ӛ�1���&r��L�G��R3Xi��A���p�b�����_�d�f�����μ�� j2�N�6O2o�62Z�FR�R�q���G݉��(��Y�է��N��X�^�&}�l�9���5��.�iθ�u"�cb{y�����~�o�$�:�t����x�Ֆc��AFDlϕ�9����C��[�.R�oh�濫H���cs_�,��63���l䉗>�;�Uϛ���!�T'l��FK.��!���c���-: hjkk?�p�
���ÔOb���TK��'��&���峏R|^��B��u���:�K����(UK����%�o�P����%������W�Bn��k,9N*@�����J�|G��p(�a��幡$~`?�)V���2���h�����|��3��Y�a]�*h�m������9�K�H�{���ޚ����T��R�[�v�u_iP��(�.4����H͍L̀��-�1�L��W�H���%�[��U6�8*Ѳ���6��6�ቅ�<�+o����"r�
���u0��%��$ִ�#*��~o~�S�㮢��V�.��Z3��>.�f>�T����Ԩ4�K�8��1���}�wJ��~�
�����"��U�r@Mg�Y{�:}m��1�D�^���V�~�aTho�weC�@0�2��8u��l�PL���@ʁX �{�.�˴�g�[������z�%���$��L�/�������$�RCC������-���t�$�e��D��ؓ���{��	���� �l͝8�T��G���QPR�'i��o^�J��:݂��-҆�To�'R~r9���$���ܙ��鹙KyT�À6���}~Śքc��Nnw���a|7ޯyЦԇn7�5��ڼK=E�r�^��t�N��Lm�
]�Oc*��4/Y���4�Ȳ"���·|=�d%�0�%�S|@��Y�p���n
�Y�����Ŷ�q�w�1�cmr����Dx�\_F�$f��I���&Ii�����uInN�vJP<��O/�7qGGGHY�#����84OP�}�u��f�W_�o\.�yΆyV3vb��J��ʾ�Ђ\j"t�{�]/ƚ�m"9�npT��45Z=��a"�8�*699i7�TWh�r������ֵh�v|��aK�:=FUU���:�{��&�oQ��?��.f��	flH��7��2v���gO����/�z�֑��=b�my���������&�\���SW�5H^�z����7mG��=��5*�Y�܏�}w��M�g���CA>"�xrL\�~���I9�b@�4J����8f�{)�]�c��,���O�ߌ_Ā��e����j����޲��j��Q�͵Ũ� ��q�)-K��Q�o2聓���emO��mH���#���M��
#��^G����X-3�h���O9�Z�Wf�ƭq~���eg2��#��l	��/���T��Q����WX�7��Po�����s�#&{8i#��VUt`i��O����'����ٞ�t�&i� ��o�������c��|~nϨ݈)tM��z?�v��&��g��ED{�ǡ2 [�j�b�����C����]������u"���`\o-bW�(ꛋ�Q��d��ò��Y���%$H�Td��Y8�?_��i��zI ����9q�s���3u^����I7��s��"
�Z�RHk���2R#>�4�&��s�x��|���B̫��Y=F���)l������lt���Z1'���wloiV��X�y�����M iz�c��>=ֵtw�h�N��V�G$�*���+
�罇�Y�ҽ�w�� �IUr���+��t!" 2��bQW����ܐ�g���%{D)�݁G{�u+%_>�5LH���K�6�C�P�0	�T�J㡞�4�Nlx�^:�I��8���O��� |
#S� DZ*�*e�����t���$��d٣��N���Jo��ڱm���>��������YM�F ~|%��]��l%R%co�PhQvPH>�PT|�����������d�]e�	�����}���6� F"؏`��V)�I��g9-w<�]�8|��.�`#�;#i���:M�}T䥹w ���N���
t
����@�	)OԘ���jHi�8���V����HlRR����`D�+��$l��1z��ў�_!�S���*�v�ݳB�#үsn�GY�=aQj�/Y�1�TBB�`�6lbbTߎ�Hb>]�(�1!? �\j������D�꬗C ���^�B*FHQ���}{�	p$� <V���ØW�Yz��?l-�ct��o-]W��|E����;���з��p���'����DQ	f��4�t�
�L0r2������~��q*����7��{VGGݣ��@��XS}�sY�'d�F_��_�� �*{BҾ@�ۂuZ���
1:��{���[�]�����F9��#���:��Ԕ�ׂ����6��r=�e!@��g���98)T��Dn�dJMA�퍘��Y�t�dc�W����g��K8�e~�&���F���A�,rl&��͊;F ��������b�
�P2�\�l"�����Q/9%%^��$�8��Mc������w�HSW0G��34��*��A�1]��=~�T�	4(�eqJ~J齰r��V-N�>z������T(�������E�ߩlήu�5E�{n��7M�+%��-�<j�Z���4�&��`Tb�1���A��m�R�g.$� ����N��eN����� �,9`�I� Ƽ�yyK�mizM�h�*]�T�=�� Daݒ=J �o]�%� �3�6Gк�JK#BZ����X� \�wO7����FQAz'��-wD�����ht:L~��0p��||�����A T�����+S��Ync���{�����q[V�*�s'@bTQa>e'&������qSH�`���}g 	�3;@M���Ke�/���%��g��By��lwy��o�-���<$�g��)�c�j�ULRC|��	ǅ$����5Bkrj�`�u�;�������*c��2�C;$�"��E��?����t6����spppi6�͖� ��J ��/d9_�(t�koo�uV�Xgӛ�er���}[�?�a��YF�(f��}�N/���͂�sV�{G`8�OW�5f��@�&��`�/<��|�:$$���r�3�]@�L7,��t���\�Yb�D�;���YVNnYg�8k�����bU��6�ؾ>i�4~U0*%%v�*
$�j���G J�
�YK���m�Jz�\V�8��<*,Ђ?>j�l�{~}��ď��F����VgR�*"���C���͹R�b+�q�u��5�k��Nc���t�B�~Cx%mJ4V�K�x4��R��5|v�oe�x|����:}P����,a��5��e�a���թ��L�b�P^�KokW�̳Q;-�U��f*���<�~pP�'��_����P�����?��8�A�N�:x����u�xZa��-�Z�j�_��*
����тR�ʛ7�����.�g��	��ZFqq���x�Ąr��!�#��P���̗��	���3��~SV[7�ӄ�)G���($���T�^�t��,Cq�I������JG��֍�n2$$$i99�C�iV�)���Z �rn�9���%}O����-Y�{���J�+sbA��M>u�����%��-�Q�ߔ DJ��z�(x���S�z^
�^�z������6�����:�N�������"$I�a�d�q��Ėw|u;�?�ȁ����5/�CE���|n�9����!��-.1���SݶM�����S�S����N�_���%O�~���|ܨ$~k�ޢ�E���h��0�n�?�n��`�ݠ��G�Z7j�͊8�L�X�
��?�G]�x(�T;|r����S���FR��ed�j�8�-	{���MD�4)�;7|�k�l28TSW7쏦v�H�g�}�}Ӱ��{ٌ�W�<TDϔ���7|c� H���κ�J��L�����K��R�� �P1b:�������&���(
����x�ٻ�,:�4�I�]%7�e�ij���F�I�����v:�pX��.%����7���}_A�pY۳t���`ab��c���x���	k�ё%P��
������.�Cּ �����?�<^����5m�9���e/����?:y9�O�}��L)�����޻�C���d6إ��W�C[6�v�����,��\�c���X�Ts�l��艉4Σ ���
�ǧ�ޅZ���P�j�mw;)lᰱ=R�
�/�.o��h��>?p��oh�����[�%��tyr�t����l�}M���_H���b�v���		� "Vh�?]�bo_'&��b 
WII���6���^��K�E�D�A�|�p�����)�����=����Ԏ�����Ƃ�k�a��xe�Y�|}��g:�5gP����d_���jp0�������_�s¬V���Ô��o�>��f^9Y���Vf�?�P�.�s�Dˢ�Mi�$:[�� �߽;@��������� �Ca�,�9���1x�7��R��0���w�gw��J���M405�Xb&��,zC�|Kf&�o�����\�m�ڢ����p ����Hpۑ���������L��JFp.��,��m������%'�O.�,�sq�h�.l63�޿o求<2���ʼ�h�`�h��g���=�G�M�~��q,��;+��vC���޿ }�)l~�KY~�Y(�S�UCD�D���-�}�)�h��#���fT�狌�oWm��ֳ�W{�mmR�fk�?��n��{�&re�a�(ً�����/@,���5j��̀��sޏ��`��V�C�������`{�5�r�z,��o�rs��q�q���z�W\�*�㪫�H����M(�R��R7?�ys�evjJ�P*��d*�UҀc�B���T�Z�/:����b��Rq&��n��ԏ H��!���{^����u	�����n:MM48|O6�g{�ρ��̳�a�5� u ���pޒu����|���{���YPXX,��R.@��uti���Ǧd��/�_�>|@���#-��Z\*�i���~l,�����ǀ�8��Y�s���?��,��k�PP�{�FJ$dii��;�.�N���.���n���<��~��������33k��ֽ�{�!S�2�oU@12I���?݅z�F�G8�_p�����t�����Ɔl�9��
��ZX �ˑ��E���� ��Ů(*	z5`� sf��
hr^��7`����P���!��_k�`������i�n�ԔU3�����=��������'�M����2�op��|���}��%���J���4��,��J�ʋ!?�����>s�tLE�M$?����Z�}h�o�߷��R��n��ڪ�K/+���ٯ�
��_�҅@���!��X+�d�ԃ`x�w3fUM�""�A�( ^���9N�?�Wm6��Pc�/�A��7TV��'�� ��-<2u�9P?��Ġ]%Џ���*��5=���X�vH�������3�I�����?ГrY�v@=a�����+I�1���!��fv�[�I�j�(-��6��Az��;�d� �a�׶�Bj�z���.F��? N��Љʭ}w��V:��m�j���G''sf�`0���w]LO{�i��Avۃ��"Vr1�����gˮ'�����D���Hd�%qYA�$0��47IIDn������3�W��i�"�L
�GGw Ԓ>�������c~ш��@>����RܰsC�v~���O��@4�G�\�]7� ��4}^3
�â�΍�ԢY:��%p��qա|�l�}�OtY�,��97�'�a����"*�t_�6l�|�>�X[[�E���B�C
l�[�%�٭�EE�f�%�	�2�g��\�|H * ��w�Ua�	q��K��=F^=H�łV���BZP�%�^9} ���t<Hz��9�хZT�dO���ljw��xj���%��t`��zL��2W ����{�7����64��(^�^G���v�� .V�|�y�J����ng�O�,�C�o��e���a��ʹ7`8Ή�yv�E���<�n���_Ťl{:ox�%���]o���@���?S))��0�Lx4򋋾1����K�)���3��XP-@o���^woB��Y��nhUJ�b�=��+ �*��SI���Xh�(t�-�?�}������؂K�:G�l�eq���']���Wэc���OI��m�,�x��7��K=�`��8��E�O�PN �nhj?Z�#s�3��4m��T�����Dҋ�Τ�cQ�Zpl�)�R߁�$���І�'�`Wjў`�V5�#{Uγ ��|	�m�|E.7
s�sg��Dh!�`.������ϖ� M ;���;�P�w��v�?��4��>����� ::�zFñbQ:��ԯ�!�Pfw]����/�t
=aLQ�����$�쬧y��Sv��W��DDK ?�wl�+��f�%dяYZ��֠3>k�r���Av�6�V`jw�����������_����T߿���k���hr� �`�h��.����Cw���З������T$�0���N���&�:nn����]�B�$Z� !((	�)@��7�z~�q�Rf��	f�9��5���Z} �ܔ�|	)�֏�d�?ήo^0�?ӘZ�ht�~�gH�A��Oo�K ��f�P0�$���Ia�9i��)�Ϛs5]ϛ�y��񾟟�]{�#>~ 𸁁@H:�������c!�￁���i0M��* ��C��d(�n� �a  g.�A)QQf;�t�W�z3>�����"�;ĺ͒����!s����)R��4O�O2�߮`����xS{{��8l}#$�@o���yi5��[��+D�U^��E������O���ӥ!�'-j���_G�mE��9�eu�Ѓ�FiH(#c4��NQAauJY���K���A�,2�T(BG��P����@�j�0�����2��.��G���4�T�\�d�Ȁ��,���iI*d��٨ͅ������u*�����K84�T�ї���<�Ma-�Yb�F����i�j/�?��[0�����.m}�̬� ~1H�@���A��{%{32��}�������,%iX5<�a��=Ƞ���� �v�8�b����� 
���Hc�33��رa�/.���X��!�{p�Z111>�2�M'�ە(Vb�t=�$�wQ �d$Ȼ&��ֻ�ʑ��X�����T�@u!!!9���"p�3�j�nw�Q�,�!D�yxlw�N���	-���;0M�{-g5�(����M�.��2ͯ�)!�H���Z{��*�t&����'i <�V�Yt9�J�q��SR�p"
��]Qӷ�)i��J�OS��fTm���� n��F�"J����=�t0S&�̧#a�dTU��1Ol�o�I;�ԣ���%1��f}I�ʄ��d �`Z��X�jP�Y�#A[����m[�By���o����I�߲]+�]� &�FÄY�?����� ���Eu�T�zd@l�ZZ�h�)�I��V�cc��}5��ь���hN���3��u�^�W����`R5	'9��;D�C���m1�tL\dz�)�KO���?*(����2�O�i�a:��ۤ�",��Ĭ��̢�`�Y�|�S���MEB�������-�N�k����%3V��<��fe�--��ͭ�����	}�]}�������x%A�Γ���C�z��2
��Zb�v�S;+G��m�0���.SA�y2����5�6�
��?����X;]����S�Dli~5����YDC#������>�
�w��{����;�/��Z���Z,�\�i�xj��$��l�N�a�h�%�j��9&8�V��s����# d�������T��+��@Y"V*�Kί��L��$������	f��S򅘖�����(M�j0��v9ˉ�}��sPp�?�ں�io}��We�ٸ$kfM�$V��jE`3�����S?��5��Y��ʎ$��bh���MNN����\/1��+�'<d���Ś����q������e������1�̍zY��h���;�&9�3z��o����A@����d�Jf���Pҥ��U����}K�<�},l0e���$2������;���g��I5� ]4T�w�c�
�����O� 9�ڪVR�~Yv�����5�.�R��ӫf��
/*��4���u*f3ʉ��/ň̢|��%����{��7�|��â��2�yڍT��̖����r�������F�Mv�z��v�d��M_�<�;���j�04R�@@	�4`ߖ��������Ne���Uk\b��� '''��n�!���f�J���C��l.�Y/?d��+�-V����{bb�
��9�]>��&���D���MU�2��c�<���=��D���P;SKKq%��CR�����~�ӹ���Ƙ���=�=���7�\�vǄA���->k�ޠ��l|J��bK=J�����)�9{�+.j&�,@i��3�2�q��W�g��p��[x�����[�a*�N���T�Iy��5�,�H0x����S�׿�|�X��7��%�^	2wߩ"��qS��!���f��+���xP�
���Z��b[��ͻ���=u/�Q�G)��9�ǲ�� Ts�(/��=� " w�CCC}}}���.�y��\�9v>q���'��D����'�S�l�F|�-V(q|h��My�E�"1��d��H�ٚN������`��H/�PR�g
e>�u�|a%�PGp�H�Y�k�!�ʓTѥ��:��s��Nw��$g�$���W�S�/Dc��1t��/E�d��A�z��{���)��+�$�)��w |z�?�8�|C�0�K�:3:�u{�C�ͭ��_ cs:�&@9v~�,,Ddg�s�N���.Pb�TT��MN��,��P�� n��jm��0^� �f�\��`RZ��bg�wBF�f��JN�,e���	���c {���A]�^GxAFp`�q~-<�SqC&�tu�CMDU���`�7*e�&�����Y�����$z�¨�K���VR�9�gF�e�Y����x���ZG&,������|�����'D����$�8ܾgJ\��Ŷ��;�Ȅ6Pd:l�V�*q���~���Ѡ�&�F��yvm�k����69�+yWPP�:���ٲ�d}� ���I�|5�pe4��]�Xd�x53~�Ǫ�"v��:'�ׯ�ng��u�Ǎ b��o~����,S�u�������7�mJ�*�w.:�;�?�9�]�߬w�Ձ`RX��,F��Z�t���wPyr��HM��3�tޟ�U��}�t@��G\!�u�["5�_T��y�as��A���V���L��WL�b_3I�uo�c*�m~�����(��'t�9����������L�?���۷o��V�KJ��_IƳ���X��$5LX��<j����VK[���8�� �A�U��p.(.~-.���B,j�G?~�=��m�V��"����}L�W����cUJ1;r҆���[!HL��8���-C��ž�NL�n�?���ֈ7xE٪�Qj�TW8"瞭�v�vL��z�e��IW�[�Ə���?4@��p�(V��=�|��L�����y$L����-p�Fi����<0^��nO�; a�P�]��M�m��fך��L�F��ѯ�d ��ܼ��ݧ-��LMMO�z�:�l�;��~���/&C!P �%�����h7B�ã!�L�<�ե����q��>9
���^����o	ލ̾��g�&.̂^��:�?�+vC��� �M��L�B	e(�����{��-y݆�5�����$�ܿ ���3s� ��k���� ������MJ5tQ��7�e���Q�q|�w�ޭ�:.��UN�\Z5B��A�}%S���G�+=��:�~�GU��B;n�~n��B�5�`���²Z�Ng�">iՙT���$p
S4v��ꋂ� �J
s^ ��v6�s�{����bXQ$1e)�'�����P�8_�BɁ�9�N1q��0�ZÁؗ�V}^yj���oߪ��A�]:Ɓ8�Θ	d��o��^����.ݍ�!�SH�wh�EU��YP_��Ύ�Z�����ZՒAO`�r�)��.�&��H�B�JFE�{�AS3�
%�zt�K���	,��Vɉ/�RF�$J�QDĎ58
�������!fe销�2�]�׼��J)n��u8���3g��ޫj��X��@��<��KyW��踱���-���r�\�����ZJ�oxD6�cu�7xS��\\�C�+]c��'_D7-�I����mgdf
]-ㅼ���n�AT<9*�$N����cV��Vl<�-r��wz�B�ķT*�Ŭ��%�F��o�XI||}��L+X��2wj��\Ep��) &�@qG^j_���f�YGn$ X\���Ϸl�y�'���eddT8p^�z���X]Z�(�p2�pBÌ�:��4�X� N��g�+�6��5_'�`�sw��c��k�ϟ:���@m�k�0�2���N'U)$���}��/ݛ8ә*�?0٪�0J�?�� �ڴC��(����g�gO�S�r��XB���G�]����=Z��E�c8|���1��C���7�l�S�t^� P��K�R��}USc*FǌJ�t'�|�\h�sҲ��U���k���	�z��G�(� 0CF��:��b)2+����W��}�c,�5՞����" ��@Iik��&n�Y`��ꮏ8iH���� ��(*Ieٶ���Q�2�"_>��qw#�,R6��*�ڍ�"��\m��R�Yi=C��7�ox��v�#������X���ES��!�z �Jxk��r���b?��x�w{�E�̬X̂��k�*�rp��ƹܟB&
�ͣ#�s��hO������s�㌣������l\>�+���C@>9�h�Hc��wS�|K���O:	�;���_V�a:#�(�4׃&�\HY��v�{zV�r��>��/5[�����B;�0j�T6��>���"?P�#���{Wz�za���X���5L#(HVi4"nk��'��~ߡ��z�j��=@��2�(�_���A�x�}m6z2=��؈�v �w��=�#�Yts	V�|�44kȬ��rZ��qԬ���\~z��<'Ñ�>��;�'������-˼�ڵ�0��F����;J��4�g>d!� E��RF���9�M��J!��D��5.Lz8�j)x2':) 	��&P���Z�sK�,ML_X�7w<-�jY���CҬ�t8�M{�%�?^ȯ����JNF����<��611ٝ����ɘy~*ba|\.��N"�����EiiQj-��]*����\%]�Á��~WW�ÈY���PU�Sx��%"�����UK��(�Y����l�Ȕ�Q^����QZZ����t�G�ʊ.Aڝ)�į�V~\<���'������ŧ�?��w��
�v���l9L�AL`�/'ť��Fs����������� ���}�Ⴣ���%����FG�}�}	
�w���(D| ֞Nc'��`Ӗ�Ce+>o�ͽ��z�����c3�-�&O�-����Gா�r�H����h��
,,�u�z�ʛ��2	�EZʻqqx�FFT`0q���hy9[��{������旔�M��w��R��(mnn���!�n��~}����{RDd~A�ڕ�דFNI�
!��2���saU��.Po֗�1fv�� �\0U�e�6$E���(�1[��}#|mw�!K�=P�^�|��h�M\�����&?n؁�#�5V��ĳ1� :!��`��%J��=���%- Y6A�(�#��^�m�:��� ��HНr��=QEE��`((�M�󰧦��KK�@�F��W5WB����׮�!��x��׺O7�6S/Sm:wq������O�j��ffh�&������찢����k,����� ��X�X*HE�N:���4�M�N�^ɞ0]��|I��^��.�͘�~�B��݁����-S�^9���p_�����'�́X�q�����Yw��c��3���@�(�y�חj.$��-Ɉ�"u�����/)�x�ma�#�Zu.D��/Uu87]� FF��oh�ު*yGW�@[T>��/*[��_��ͭ��5�C���0��fT:Qo�>b�Z�q���)ތ6��C ����l��ߐ�e�Mx,I4�4r����}�����W����.8�O�o҅�Bp�TD�,O�Qz��RBrȹ�}T���w$(���]�ݾ�LJ�Baj��\u;�N��6��^��-iW�=9'[k��6<�߯��ā|���;#��2ȷ�1�n���M"A�I��n����w%�=D��[V��P�B��Fo~.��8j��D�LJ�r.��O��P���}z\�`��u^eh���lnb?���܌o��iۤ�ju�N�Li��i8ٺ���)�%��Nz�+%z=�9���K�3����=c�_%ݴZE;�I� �ޔ?_v�m'��r���%(�As. �V�KI�_r�}�R_��7��*+����ɗN��Q��:���]R�ϓ���n_x��f�rc���{f��_(:H>kkL�ɪÃ�~g�{"$��A�t�Wऻϑ_f��G�<ޭ��A=�Ji[9�V%�����C���N�Z��q��h��W������Sdt9�d�g9M#LŤ���K*`�j�x���;�%s>k����PO�Zx/ x��)���2bɧ;��}Y�9����vp�Bn���(�o*��[�q|��Hfhު,��;����}�t|S`���n�H�|�$�N���g��$!^R/�:���;���O�ׄ~�D���Gvz���c*��YZ�]|�FHa){������xٳ�P�}�/^��H�I���mGk�=��
����A�+�%6�����;]�^rA�^�S�W ��Z9�=/^9O���s�����]`�>�����(xj�?K��'g��iW�vEuѰ��X��j��ymk�OO��h��ߠ߰�H��=�?��cz�s����u�Fwp�(�а�"'?E�� �gl��s�p��k6D�<]'�>��R�BY���m����w�v��^2Y�\�K�*V�lD��2Z���v�C���4Y��QV��M��#Ϫ���{.�z��C�~���p��{h$y~ؔ2�l�ȇ~ߠ�]�}�REj( B������֞���ʟ��������
J�e+T�P�;�q����)Ԟ��_�&&u{��,;Պ�;��V:�<j	�)���U�x��r v'�'�ɥ��A�P[v��3[��K�x%��+3>���I���oV+%0_F%�P�Nx]�)E��[����f�P|$ݽ����25������ b5/�C������3��=���^�8���pv{���!��9џbX;Q�5����{H[x�O�h������]~A�ax�'��,�WӔ�X�!���R~~�� ��q������)�!oi�N�W��}�������حN���xˠ$o���B�\x��k���}a���5n:����������� �"b��H�!k*�.��O�R�̈́�=Adʵk�:'���KY��O��77���9m��5�!�7�p��%⩏�:�}��U�X�{�k�/�J���C^�\��|��F�wY"�C6UP�H'�>���`ł����`�D��Fif�`Q��'������M�R������V�1�����V^4��隳R�έ0y[h�J������x龟͘�M+����S��87瓷�Ac^e��!���٥�>��
��
B�6�l$xle�Tc��
s�ސ�I�|T�A�qoY�̣���7��;:;O��R�p~�����ڂ�W7cG)3>j.�*���j��d�{�nS	 
=���y4�{4�mX�Xē�
G�X[�[TM�->8<.S���W�H�eWkҤEDZ鳻ϳ�Y$V%�00����Gv�z�-Y���;7E#��t!�
�T/��Sw��g��Ѧ.�Od�Gp����4�M��}mY��ǒ/��e/�?���8�k���^]���=��{G^���m;6�CL9�T���7dO�Љ�u�zr[��%t d��?faw;����7�{$e�J�	��*J|��L5^���9��6��;�z���Kψ\&|Fzt���^���J�b�#�?�ғ��땠�8�L׮P+a^$��vH��_}��p5�;�O��e>�;��jr�~H/���CD$8�/q�Ű��h �M~�i�1E5�o�*[�y�Έ�=Xs`�K�[���Db�Px��3�a�QKh-��ՇX�KN�h��M����\�]Ǽ�� ����UK���xQ�7_�aɔ���s�J���zf���Ҵ?N}�-��w��	��K��N ��̮`q��f�U��������m�{�;)�H�ZC

��M$�N�l�6�ts"bc]�۱�#0ߧ�Vg��g5�G_���<{}YB����LҺ����_.m�����
������zM���h�;ewGʘ�קq�M	GR$�\���L [�\��W7�����W�̷ӡi�5w���@�`���T�*k��O��x�Kv��{�]{K�e�RRϦ��5%�͡�f����H$L@���czǇ�ڴ=:�KVa����k�kFy����M��,f�Ʈ����9�xht�tr5�@�oa��,Q6����E���탉9#�K-a�1>j-`�I�;&�ӆ���_���h���pbxi?�sB��,�t
�{�b��ٌ�9IGu�bX�T�	9]����Z
S�@y�?��VJ߽�RF.��4�����$/�&�;M�s}ynօK�w�;|Qjjᓨ�h���<A�s��Z�@9�w���h�������z�m��9�PA�p(�f[��U9���H1U����}�]֌�X��,AXtL��Qm�Su&�T��LJ�뉥}���Is<u�61��J�$+�`�k��ɘ��ί`>9�IT&�K��7�N�����,�D�/#{K�ŀ_`�O$���4�?gL͂+���uy�\�h����k��W~g��^�gEH�.�}H���o�B�l��3���W���q@�G~*�eV#�����l;3�L�Y3Jz�ЖM�㕯�w:@s?�N���&ҋR�Fe�Z�c�1�mk��*�n&\M��/a	S�MՂ��0�t�o��`o��ef^�M�b�z|
(nBlz%U(�4�^�EE���?��̳���\��ݞ��8��^35��g�t.pwջ&.��{�c q�	P���wtvw!�AAqP���h�	|���HX5��N :zùݠ���?��S p�zy�EY�/�; T89R"�v�fw9��%������ڴ��K랼��*[dI�����/�l�e��Ţ��~~��}b����鉚�҉_^��x��l�(���Ǩ��ax�L���F�oZ�������Ez4A���Lʇ��k��*b�=ӲOw<�]�2� ��qd�}�j��տ�`�ѧy��W����#�� m~�1�/�,��F�uMħO��d����D�(M���{��eO�'�G1jZ���"��.9(���L��OeAH�j��9���R&�p�'v=�#�{AyI,@��0��E3	��p���pa��R2�G˟�
��"��Y�&8�![��Í�$&��Ѡ׸z��b�Z��dF�=�yn�������B� ��N���Ah�bGoz�O��EZӖ��̻�!vg��5��h}ٌ����8� �^�֞�xu���oŐ��Be�����)]g��C���(#��8�6®�g�v	@�4>�E�Cz�:ڶ��n����v�0��ᇜV3]��~I��uD�l���E5�r8�����)�1���� {�Ӌ;"ql��o�xi��(���K:�"{?��7��?R�UӗZbͭ7�-y�O/X�){^�҈s��gƙ��s��y�0Zn'�]��#B2MþH��=�K�Jի�B1���UDS�t�]Z��h�>�n� I��cʒ��	�,2��؁��q����h�h�����1����wF0[^0u��NZYE_���Z���.+�63G�ζMc���X��V��s�o*���̈���_��{Jyb&s[v�3+�8�HZ(c��y	@����0ڷ��v�`�(?by�Lqy\������3��!t������	���g��`��7���t ��������|O�Q���h�<��$�R��~���mSPg��Jp����aNG�:*���$��ށ�k�<6��)���Y�8�Ys㡹��4W77>���RR(X��P�srhE�0�&��pX∇��p���g��*A�DD�3��Qw�D@'�����uJ�*(���"��?_r%����===�z�Z�M�;2..����Y4M� �-o=b(w���f��Lե}��
�9O�Y�HH�-l2z�N���·�9C������9�7�G?���o�.Ś񜹔�$\�vɥ�dH)��o�'��A%jo���k�z`Rsn|�N��϶���Ő]�3��?��aN��y~�1657��!�"~��I�7�����J_�r���Ro��
;iU��])װH=T�d��$�YqbF@�gg}��\���9Z��>�Қw����?�^�n��q�i����+�vΐB�1��%zwۼ�<5N��i7e�5Ӝ�n�"_E�_���;kT���1#.®�rg����� l'�H�^L���a�5X��o�v�C�Ӛ����ȼk-A͘x���#��O3-��[�HQ�+�A+R� �y����(ճ��4:��<\���w�_�7+�`�^��d�-)��[�4�` �c���.}���?%��}[�P�~�F�F�. �]:1�I����[�j4/�z!���eB���fJ�0��͜�?Ӛ9-�#$d͉ 6�.��>>s�&cN^@��PFd��lR�8��<aY9�㮬Ŧ��+P܊�>-䵥���y�X���
Z�@MzWC�_�A4i���K���R�1ܫ!��f������bf�7�.Jew���Jbf�U*�G.�*�����̞-�)2)��#��f�%�7��u��=tcV�jDF^s�}�<�Jā�M�ܕ#:g���0���u�j3�O�	�#���r{��Z��2p��u�b�W/2��pR�vɨD伪�n�E���>�����^���%��5��I�Vr��B���Q��	k�!O��";�F���ժx�N��r)�ޭ6����2��w����B����HB�0�2{���NG����s��i�3���m��ϡ5k��>�g=�V�j�jU">O�5�A�?\�u{���b��&󏟞ꡯ�D�tj7�/0�!/�����_5E�]k1����l�n]*Ux
~ئA]�R��$�s"�$�!�ka}�Qk����Y�Ue̐���p|�>�X�i�,z��l���7l�'c*[�
�ܟ��>�vv�h���8!�B�{S�i��+`���=Q���R�����R2_�[E(14բ�cΛ��b�.�o�S��(��ļXN���6�t�v�������3
�n-��f	U��p��|�>q��� y'FCK��է�����A/fV�)�a�5/r��Q#�+Y��9��!,
ɤ�Բ�/�t�d	Gi&K�=�J�x��V�6�/}%&��C_a���8�"���גZ**E�;+�r
���ό<� G���׍�oBY���^2�R���Yg��Be�Z����8���o�]�[�{Q�99�u�phi�o�#n,;+�I,���!"^���7j��^���>A��9:3���*k�1��m8���e{}�\l�vԷ跾��/����6n�1e:������ ǥ`��]�i�M��'����Am����]�r2��Y��g��c��$vD%o:����;���s���p5�-�x&9�>�^�0�/ΰI���F&U��{Y�8u����~���d t�i@p����z�Ms����C�����^���[�O��jekK��xKF'�)o�0�r5] �g>�/�J�Y6�K���Qܯ4>�1��/�O|��$�������Hӏ���$��*�e�f�?�h�]�f�
9�1�,�a��S0�C���LE�*]-C�ޙD�8f�RB<�>
/�{��mr�fݩ��j>{՞"���d\�c��nƴzw���z�[ͪ�����ZGA42��T�U9
����=�ݤŗ&&�K��.Wǰ1�w�b+^Z5߆�=����<�8T;�]]'/h��d�����s�ߟѢF]���&~',^�AW��_�Y�|���؟��Ţ301���GT�j+��9`�d��e?��6k)kiѣ��ђ����'�G�to��A���n�2���K�xQ�uT��N��l~k��-#ˌ*��6�D7���3��H�҇���ˈ�hi�4U����f!�e-|�������A;�OX�#N��Q�܇���ڬ�]�����j��%�w!���^�܃����(.&a����L�	�]��M���ԧΣ��[8��z�����y�z}��[�4�$(���ξm����J� �a�x���/L��d�=��t@�0���EK1�r��RpF�Cf�����	�N��C+���?�zH~�T���6�����cfg5n��g�m�|ޠz�d���	7�x+KT��C���c�Y�:Qt�;�<l-W�D8Ih�����4?oc*��s�d��9��Ҭ����G�ٰB嫪���_����M�$?p��ʞ����z�<�����`z	�BB����C��{w7?�9$L\]�M�jEH_{U/��v�%��SH>��L�+J��/�&k��0l��ۥs!\���]#Y���7\��������t�	|��Ǯ�AFJ^%�P�.�I���8T�	wB�f�<=k������4�3e�߬E�Z˿�8�����W��8l���������fc�Z*��d�o��%$��WV�R�wXR�ogL�9D�ѐ6�D/�!
B;C����r'�R�"$�٤�}��َ?] �T��Vs���z䨀���]�؊���9?.�jQ��W��EoJ��;aG��o`J��ѵ̺��Єo�׬3�Y(|G�]��$����5��z�&BeO��BV �4�N7*���I*��Mޗ� j��I��yvH�SeaF���<ԙ������X��Ao��!K��z��̬,9H��~��k����
�[ֵm�Ww�ןʪ�Eg�VBmPo��yJ��Ą�ς��'��ɂ)��z\����Y�|�X�gլ��0��6����>bv`r�����UF�h,�/���ي�ٸ~/H�T+|6���ˠ�3������c��w�8#Y�3�pne��n���7t/]�곍��8�Ju
e���Uc�T�f����#��ڂ�PNǳ�Oz��+��e�ŋ������rB�XO�n�ؚ��D���y����<bv�.��l� ?��I"��YׁH��=:*�3�ߨt�M�5�e�;?���}��&Z�Ǽ�G��[�|����i��QE��ϩ��A�q�U|�0���@Tؽx\�H(�{7��l���5��.��q4It�	������ov�]�.-��Y#zⱏY�hJ��ɋ�s�*�q�c]�J:��V�h�|�J��l������-Y����L_h���rm-x�*�Y�Z�@3�ڹ;BzVeYԱ��FR���O��;ǭZ~�|>�/���u�K�1ԏ����i~�x��]0��Y��d"�r�^���B���9�B�8S�ӤW#P�����<wN�ҟ��MQ?%ty�.1��.Z��S�7�9U�Jḇc�?VC����~�nu�n��j-,'g5`Wb��i_��9	��¢E�q����`��d�K����)���ۨ��Q�烴bR��%���	v>�0M|���l�>�H['�"����9o��͆K��y{a�I�t$��\��ǰ���-0�W��|%���н��z n�)W�H�r1)�fѠ�&��_ J��pG��uK��<?�h�������W1��	�\�J�嘻�-�Y"�d��p�ĠJ���B0|�٤iA10�/�":M�%�a{n$�nR��_R0������
N,Vj�gX������MW(���}��S$!���2٠�Ǌ��y�Z��^�e9�,�h�XNȂ����_"0�o�h�Ȳ��x����T�*"7�8��'��.B���z(�F�Q=���f\�e��s�B*�M���5���l	C�B#D����O��T�J�1��[�ߖf=}��U5G��OD!}o(�y]c�@eq���{QFR��pڃ����o@Ѳ�0
\h�k=�N� o��ڤ�+o���~���'��l.̲��&_&o��0�C_T�?-���� dȹ���kI�\Ό���^w�y�\u���f������<b�}�n;iō��«�7˲���j.���hV��^Z!^�bA�Khd|(�`��΀�����1���UNi{&G�um�0��Pf���}���@��<��]��t}��"��U�2#�⒔�	)x�ұ�͵[�G����O����1���+���?���h��x�5#�,�1�{���M��+���~��X@M����o/�O�]���Ц��ݮ �ǋ ���g� �J/��ٮ]�Б����^�����+�KE�������'�Z꾕�y�" ������z� ����[���o:R�!ґ1�hż`PV����u�6�@�|����:����T���7����"�)2��mK�h���O���v�n�o`3�<|G�x�IZ����>8��P�k�A��ۜ�F��Q����X1uF��# �lʼ�'�ȤO��;m��t!�L�D���٦zw"'���s^9�S|�0�8S ß0���k�m%ś�!�+���2(��0S��%fq����Lԅڈ��x2)I�����sT-��Π����K�}6��f'%�W)�a{�CjGOA�X���3E�E�K������|mK��[4����4ys2e��_ǿ�d�4g�j�y��w~���d+tyu��^ �Z��~��;J����EA���`����(��'MM+֊�?����đ�Ԥ �9'�����U��-Bc�_<މO��ru	]�g��KǬ�R�͸`#)�I���e�NÀ� �x���[���@$��W�1��4uOt�*E��/ެ��p9fo���Bz7�:@3�i��$<+?�����!{L[aĩ����Ϗ`�V5�����t��m�Z`�;�S�=�gm���
��W��bf%�f�/V.%ة�6��j��W-�%x�2u&&���.���W0/`�l� ����l��%t�QW)r��l�� ���  �N��`�\��o!O"{�d�.0d\F&J���h��G�`q��0D�3������:rZR��/�1U�_H.�>�:�۫2[6�}�p�8�-}�^\���i��|^�{��#u�p�o�Ca���A�d�{�:�)����LOe?���rL�Y*�r^tv5-_x��m���������xe��ƚ�_f���7'c��pv﯑��O�_`x#$��1�%�r�<t����Գ����l�!�Q� K՛��J6d��G�^]���a>&�3��"�4�NSZ�ȾJ��R*z����\� \��sy���g�`�оh��N����!��[{�ֺ,o�Ny��2�v��À�=~	i�FmEwd�odh�$*�C�"J��o�Z9J�`�I�Q��(aBtT�����ߵ��?{�j66��7�{�k3
������. @�.-��� x/M����cIsζ�U�s����Ŵ�mZ��OO��0M'��a��`M��Ɣ��:6ύ.��Lx����a��=�J���)*%�ʿ�{I(�3�CL��Ї=�ҫe�qA권f[�q��V�����G��������u�Q=W"r����f����}�7n��P�eK��6��J+��a��W	}8��L��\wNݭEÂp>�U�"K��W�t�-$�nX[�u.��(:ff�9Y��/eY5�|�=�Ed?J��CL�L����c��}'>�aa?5���g,�|��l�\��o������
�VUM�&K貉�6'��I}�+���������>5b��-
���4���}`��a8��Eřv�૿cOS$oJW����F�]V��i�:��ڶ5�AET�TP����	(�kh�B�:(R�H'���{G�� @BGz�^/�{ǹz���~�5�#Y�k�o�=�7�\{�A����I�rP��C��%���׼;����O濶o|��޼)��ѹANv��ɬ�_�s��]�۷��9�/��[9K2�]v�(����t�s	u������	���ls߮ݲ�Br6����z�� &��G�P��X>Z��Q��ʹX�mlHi|zC*�䋙J^���
t�|��#?& <^�a��T�q��V��g�&�ᱼp�k]�M����q�2$.�ugD��Ƈ�%�\��m�-�F�$ː�b���2�%&�cm� ��	�ݻ& %y/���?�L�����D��e2��yR>Z����K�q�W��%ߎX�蕧6���Q/�����G���tNwxJ%���Q��W`u�94W@�y?��r�@�j4��
]X�/��@��m�����'+��!o�6#xP2ux�O���rƧ���������ɽU3�W^�g.�_w�����o�Jez�$�tl#b�O�����%����Pzm�VW^����'��N=��X�������Jߒ$��$oF_�{�Hv������A2֭�X���ziBE���h�tha2�V�u�$����%�b?6tN=�&��)��|�tl���^�,*@ccI����J�x�+x@L�<u�V�ܙSUո_�o�����;w��Ü��2D�}lJj+V[e�M\t��(��> ���b�&C1M���N}@0�ԋ�e=�$���k��_`X,�B�+�=M~8��r��nv,��?�����~uZ�d��]ZWɎI���~u2�tU�E�đ}�'A��y�r�
m��>�1ڡ��M����{�Ku�o�����	�#�����G��� Ţ�������	>�濶]�bΎc_i&�^߬ՙ�i6=t�Q?dw[	�N��4��q&�S��2l/`�Wԯ:}�t����rh�[\Em�^~�T1��)��K��?<�i30�^�z�,(t}w&�VkK������T���
�O�S	zΞ@�~\šI*[�|�nЎm���#
VE]��(GF0�H�'�����rU��g���=��uH�Ky�Ö"�aK�d��ZVSr%`I":e�~������XU�C�3����Cdxr5��[��U/L�h�d��dQ��w��)�|�9]�;[-I�?W*gmf��^!*���2l���>2���(���b���k����0���ܹ����q���h���������#��gێd8�(�q�|ÛF=�ߜ�۞hS���"̥����k��e���q 7Z�����**7�:��� C��T��S��}����!a���1�#>L#��'*�?b��!�m�9Ф}�; n:\Ȧ�[M�eB�a��"a�?��T��Ƞn�ı��-��J�9���䎌�p���_�U�ra�����f��`��:�9�RY��ˤ�� i'LD�q|!<�� _a�̒��NV4��	��q}�����1	� ��p�x��7�����6{�32�J�ڦn2�@��S��5�sIٮ�+�OX�9�,p�=���G,y��8��4�&���/4����4�|�͵,�b��"��|�%U��d�e���07���O i���X�M&��
q��9k�ih⼓�=�'_O�<�#٧jpU�j�]}�Fj z D"�6���>ߡەJ�0���ۺ�h��|�桿'����h�e:�v鶼�o�;�r��h_����;�iz�Y߶�EӰ��Ҵۼ��4�#��XrK �.��`�����z׃��P]��V���o/�Y�r˚,V��������&ӱd���	��!|\{���
MUn�5��� i��cK%�rB�si>��|Q�[�M�VV��, �B�!I�b>�^2֘�\?��>8�cG���]1��Ku\ܮ�O�����ۀ�r�����o>k#2���p��ZqnHG���J��|H��'+�t�iS�m\i(�n{=�!H"����P, !!!�u"gs)������(�>A��ܗ�4�>���n���o��i{��?�	l,�~�e#�3
V\�|�|���	����?�8Tϣp�,l���|��}�J�=��E�Iw���![���������w�Y��6j��W��kW���'�Y�`;^��gyy���Z{z�{!��%t'�k>]�P����H�ߏM�1�����T�}�������E
�o��et\"���ٍ�R�sNe�j��aK���lN��#ܹZ�C�;��� ���;���	g#�u.�Wծ?��'\�g�L!�	例?������+�a]]�1ZQ�m�j���\�Voۢl\m��K��,7�
ԉ�W��^����NP/���ߤd����������5q��K�mW����,�`���9�+v��8�~�GË'��l��zȔ����i%]>���R�Jc,��J�v��f�ߢ���/b*?���:圃����1�����&^v�5��4��7H��:$rCg"2h�������a�H4o�4��mO�|Y�SƋ���\�~��m.������s�$��s�4Q�k�T��{�-�����8�r�� ���],dcFQ�����L�N�Mb�@��f�LW+�i�rc�{����,�E����
�(�at�s~��`�`��f b�0 �¼�y�Q���(SR I�>i��B=��p돀3�jS�\��x2 ��<�X���x������D��BS�,��,> �Ft�m�|�?�����m5e�T�MՍ��n�T���_��u���L��]��̓������b_�ZYxw�s� ^�6{�Ҫ�"�A<��h|��D#Vw��y���|
x]��䵬yms1cJf��S���y��f��H���~g���O����e�t�sģ �R�O�"�	��h��w. ���|���YN�[��kX�"YSeW�C��Nɟ��B�o��Y�Ͽ2SP�7���MH^�<Q9�
pI�̂&B�ø�L��D��� ˊ�=#�����Le�mJ$5�ù��h��������J�C�����	y�ľ�/�VbUZ@\�4u1�&��F��Xػ;b����HMd7?z\s�����=`[-_1���2��v������U�Ϭ�ע�|L����ǽ�h�#ge�������O{�vV��|��7p�j�yʇS�V�-2��w|���I�4�Uy�7M��B�8 ���&�_kv�R�@�vS�as���}�s&Wd<�i�.R�`_7UuF�8�ʾa�'%1�K}�����3lbS���~��9f��5�ZNd���P˧oR=�!�{��	 \�OKD��vi��2���-4�{�X�է�q�����|Lv-��Mi/�W��y(����x ��Ch�z�)��EK��J~V�*Ag]�ɨ������FUËMh� �k��Nն��קE��O��'��;2�ދf���}L��<z�>�_�'*4JGW�"|h���4ګK��|�.��՚�_�WmHUBa����/���49G:U	�ϯ�|�
&HƬ:tb,�\d����<#p3�3^��`���S{��d�	y6<�QS���y��Νw4��}Zg7vʑE`�	 ��!��U�ۺஅ�q�^5��/��B��|aO��+�?r�="CZ�a�J���)�d�0��Q����B5���hrN֝�Ť��I4r�$2��2btP��z]y���� a#�k�`�fYc���)�e�Q���(� �����d�>i[��v�V�m�Pi��-���ϟ������+3����3�/�v#g�d�������Wm'L��H�a��YRm�{��fj����lël�H�O&�˾صj�lu�DD;��_�5�N9o7�1q��FB�ţi�w�>�i4rZC��"N���#�f���:��)�c�m ���*9s�-��_Ea% ����Rǫ�r]E:Ss�z����%�K�΄���W�V?�)J�Ə����q��ow�!����4j�i�|PO�ux��!��0u�k0G��W�%�ע/ݗ��X�O��\-���2=1��k��ҁ����֗y��n�or�wM�bKQ���?��a�/1?�\v�1Kg�3�����l�;[�����fq$�}o���4��rm��k�*�*_;D|`̷�۸����1�~��MQ�WB�rpb�Y�)���� e�]���v.=f�sek���+0?�ZԊ��Z	����������H�u\r@�V�M�/������J�>�#hƐ۟w�&n�JD�c,W��5�YS>2(;��D�|�@{��PԶԦrR­��;�1Cf��[�I|�����;�Ǟ��1�ف٥����b�^"��N���u��
SW�����T�fJu{��A�b�:u�l����H�#�ol�~clD��	�NFa�ۈ�§��9��eO��W�Y��i#���s����s>td%L5j�b.�-�?+яPUn<Vc'\� x���aP{ٗ��J���Mf�[�p4�^e�U����l�R��!���n�,W�����d�������Y=1�Kb�u([�ː{Ӓ�f�lly���JFu69PX}�C�X�>?e���|9��%\�[�na���rY�N�/ߔ��N�Y���PͪD��ee������c��������g���$��>�x�G69J�/9���K����K�F�hF��O�NϦ�}s1�$�i�J6o��p/ɤ��N�lG{IKd�=�m��m��zZ���M5M5����ke�bpͅJq���JN�k�a�4ut�
-p�~:{��-��67k�̓~9���YOhz�4��@��t[��*���e�@T' S��6<F5��@\@+3��Fs\����T�NKix��r���Y4��k@�c)aa����Ϧ��t5��hY�i-'KḪJ�$��$ۍ�sn�O̪�庶m@ �?M]�E[	�|�������\�H^vJ��;��s[��h�(w-M�$ϩ�-"��R��.%�M<)V�okd�R����Y�ϱ@��h�ST2�땻������j�PZ�I��ˈ s�E-r���8�.�bW��k{��LDl5�A�t�#h5h����F�	%Xڵ8]���Z;�2�폋I�TD�| n܎a�4�l£*2��rvbF��~�ڡi��MJ��8���Q)���Se���6n2��O�xo������N~�Uh�U�HIL���@�_�ߎm
X�y��H*c�W���9+�W� ߀Z�/��J�)Z�W^�Sv_��}8��=쌔�=���;�,�\אN#Kx^`�LuMM��X����1G�4{dwfw 5�mѫ�x�Wd�c�����Wi"F9==���Y5M�r^��R���9��Y|_~�m8��bw���a{:����l�,m�+�}�r��HB�ʗ	��+�eOU�7&��~8�c)���ʬ�s�t�7�����x� �y� ��13	v3�7J��ر6��E���6π���/�k	⍁�pvW��pɍ��ޞ�bA'��$kƃ�Puˣ��*<oU���0��`���I������H��g�;%�(.�8s�X����dK�E��39/9^1��'ץ���fR?3�h�2���hw��T�ҽZ�I���LOe|O�D���T<�`o�SA��d��3#�r͉�b#"pâ�"Lq��ql��;n���y�"��/hz�|&@�7�-ʺq����;��E����[��%�Y[���Q�6g�!؀e�� ��$��*0�_�C�[��^�/�w�G�l�J*7�5�m�sIt?�27b�S���F��B�������D2�_��0F����`��n*˭��Xr̍�����@o>̖
;�C���:I�1��OI�k{�� l�ם�o�C(m|6�!����mS:�Χ%S�zNdg�=��֯j1�0��_�`�#�S�5�y��7��
��xWzE�証!hz�QJ����X�����;<�f}W�I�k����Y+��;��yV��T~G����:V�ީ����ű0���Բ�Y_�����n�"#��4�����=��gk:��a����G]H�+`8@��A�Y�+3o޿)�+���e3��t`ir��M�6�î(�mU��� b�îg�X�T˪4%� ���8�����qN�ĳ;��#^)�ӛ�Jrn����s��)QeYjNLK� ��λ������)��7{R_7e�A�G��8�pq�����5����Q8�r�fZ�^�*�q�d ^[cFy�k)��hK7���s�
�5�r�S��r������5�?vbs��J�􏱙�D_ҁ�vL���)�E��������yd#8��u��ƠH�ïx��X��G�lu�B�\0O�{����G�+��Z�Ŧ[��x*jX��>/���&��m�%`靗�����8�=Z�t�"� CK��T �μ�&�[���DU�h-��<��:\�;���(���"�B:O����[��u�����M��}�p��J&8(�B��Oi�)Ցl�H���AP9@���QK�2C[E��S0�YG�v[|Ǧ�$֬6L���E�,�&����������#"�;
YcSD%VH��8��,�W�W���-��#�j�^�ۿ��M�!-|�g��G�Ѹ��}ts�:6j���:��Ie������.;�#��D�(��6L1�͍�t����E,���6��E`av���5�^(�lE��=���p*u߆d�1�����؀���x�5Bs(�6*B	��e�r"���A�zr�z�2@�T4(P}���������B�݆�[�Q(�> �e�}��f۟w�;���¬cF#U�H0��>�=���TZ���H�H�Y��Ta��dz�5�t-�/!]��<Ѝ5��Cs���H�l���<���UN�ѱK�H�S]"_����  �WV}s�"�v"�X��?��;J���:��I��|ɴ��)��L_t��ӡhi�#+�m�6~{���Z�D.�DS�{ҋG�������y�Z�u5�hظ�]�.�5�����E�mY��$��:�!���̯UC+y{�
]"�N��6����*lz.������ݳ���bn�߆ږ>�5*H~��w/c���?]���2��+�q:�X����3"m(�p􎏹��v�X�L`t$q�)I�X��]`qx%^��-����M�uo�4�q�D2�{a��l�Ǝz,�.V��9!�3Աk�̵�����&f��f�ƅ�����m�7q�{�Nry�S���$�96C��); �c�\�e��/&
Ӓ�}�*�re� v���ۆ�8���6���9
S��E8�����:蟏��C܍:F�[�;���>Xn�Ї�,�B�H�{S�e���#67�� ��Yz"����&���~w�@�X��D5Z�P��D�bS;{����x�dlԋ���w�q�*����ؤ�%G��C��˜#�g�,����l|���϶�O����٘�G#���Y5�%����8s�-�yH2��~?ݻ}�>gi�'�x�8���A�HM3(��b���`Ј��9��?��QЯ}��0>Q�J5�'��8���vΑ�!-oe��K\�wR��}z�\�W<��f
I�5� ﺨ�ɉ���?���U��U���}z�&UX[Q����Q�i��[���V�C<7a:lJ��~9IB�%��$�a$��gӻ{�������ע����'b�H8P1���o�����ط��/�Gh��s��f������Սc;���L����r�
R%o��PK   p�X��
��� � /   images/243a459b-a2a2-4803-9716-552aaa3859a0.png 6@ɿ�PNG

   IHDR  Y  �   �ZN�   gAMA  ���a   	pHYs  t  t�fx   ]tEXtSnipMetadata {"clipPoints":[{"x":0,"y":0},{"x":858,"y":0},{"x":858,"y":422},{"x":0,"y":422}]}��U�  ��IDATx�佉vɑ-h�a%��E�����꧞���9�{�R�U,n �#���{��#U��o4���	0���nnv�m޴}���RN�_�S¯��E����%�i�N�Oڏ\m_����+e�?�+�{����O����}�����>��UU���׼����@����Ux���Oɮ�2������2�Ǘ���������p�õ��J0���2|�+��u��nφ�/���v5NL�H�����}bֆ�j��[V��$W�#�E�3d��e���?DR?TO~��:�����Ru�%����T��J�4�x-��L'�2ɐ�"��s�'#̒n��o���x��U��k���~�1z������nK~g��2/g��o����jʬ��W?��G��>DV��4up��Ԝ*}�-��^I���w,3#��k��A��hi��C�ь��2��P+��C�n�A�WRe�1&��X��Y�{��7f*���|u������x���_�o��u���;��m�������;�V��5c�F�������K����g{��it��I�����Ϸ��ǐ�������?Q0�Y_���\��k����!����+|���;e3������_���l�j��ڜ����o];���htÿ5�:�y��:3��ܧ�,��d��2b�w�O�6�W���}�_%�Е��i��Z�yD���,@��!��Σ����ikf�����L�� ($f1i@��;�� ���O�5�������N�m�b�F�ݺ]v�#o_;v0�^��Y�T�7��[7�y�a�J��x���z��xAo�ڸ���0Z�i���ץ�r�ܶ��6k���=>_��%+�#xLΣ�Y~&	e.]�Go�~�0���������[�h��=cY������5�Ð}\���h�ӭ� 6.Uݭy��(+���������.<�@�㮾�ጧC~[s�2������.5��^K$XE��f�J�:Q��;��fb4X�4���-����1S�/��l�����׿�x.�W��{���.s���T���3����_���o�M�I�w|CU%	���(~������/�TU��d�������sT'i��Û~��z5ү��:�2��2���-78^��JUQ�rQ�I���cs7ec�!�o��ݐ�������*4&D`ܶ����kdPj�S��Žs~��a
K�VU��g<U#ŝ��q������Qhs�_�:3�Y52�>_cei��ބr�ԗ�b�d�xx^���a��6".���9S�ʮ����e��x���u�����:º@��ac����F����T�� ����A=�m/�-�7�S�0�֮ϭ��sh�ڤ�-p3���o�K�8��n�m���L������~�+��*`��M*ʧ��U �n�+:�!�*F��V��G�sa������H�덪8V�\ma�<���ǧ��gFύ����޶k]��2G����=�4>�/�m��L�C�f��^���d�?c����gS���t����F�	�;m&�/���`��N6���{�t@� Tz/L�X�@�7�V���o�o�S����~���z�����M��l>Uթ�S?�u-瑟�	�P|�7�=J�(4SD流k�s<�N�
�	�o��{��z��Z��^�W�o��	����׾�6:�<�5]��z-�T�Y�.ج ��ƒ�n˨�5L����Mn��6��Z����C�Mk���7�Л�����4��tlf��=��e=�ڽ�Y��x��QY�N��� �k*��i�3g���7��������o�7ڴ-�Z�:G��j����|�<
]E|�}��t-/���ax���d��U����j^�:�oU�rX�pgz�ܪk3�Kxn�f�g8�����9BG�YF����RZy�	ޱ�v#�FO9�%e���ߡ��5�|ZO��Cf�Ɓu~�g���F��n0LcV���"��*��Zs�\�m�1[.-�V���#�Fm�G�����77�k�eff��tfg6��>�y�(C������u5�^7e9��+��ɱ�r�1�7RाS����/z3<d{���e�v_�fd�PV��x��1*�)ckx˸���_/�n�g�*�3'�wo����?ĳ�.������l�����AO��ha�{m͠��<=�z�:�ƅy���xB�j�BOT��,T���_�������6c
]2���v؇z �2i�X��j�r��5gx�l��M&�2�tK�Q�ہ�|��[�8��?s�ς��Ua\��Ѕ��aO'���?i�Sq��9;�P���h?� ��L���q@W���d���"V=�[s�F�j�eǽeɨw���9��WB>�wW
�W�������D}�G���4�Z��DI�2�y����$b_V�,�m�mt���{u4�r�8��پ]��4�G��<�I7�X�ny�9��6��6��І�">ΔV2�p.�4�zW.+e72c���{�ОT�U!�}6eJC�b ��}��4�߲i�GyW��*��,��F)WA**�XUn���y�9�el���A!� ɯ78l<U���Udq,7U�����'��U6��W�ʯ���値��h�QI[!��%c��H����/��2�){e����%=�g�zһ�:�r&U(g(�ʍ�};��\�C^nyϝK�ߤ�E��1q{��D�)����IO����~����e����c�@�$�[��I	 �lM�+���f�6�����b:�\�>.��q���lu�֍Do��M�Or��� ���@�Hua^ ��$�}����Z�^��cf�Hb�������^�n&�p��3ڹ�m��'�����ǘ�[�<1�w>��2栧.��sy�@1��2O&����ib�@���F�`�������X���kn���/��>���	߇� �4#cBmΙ��ɠ���M�T|C��lep�ޢ( � �S�T��R�fsH �m
��ovԛ8>�y�����8�2�S���a�v>�z��1��.�+Y)��T���ľ����@����'��_��|�\WN�!���9�Vei�Z���J�k�2 �����kB�F������$���4��{>�Fu}ѫR�g%3Ȅ��W�ŝ�A��ER�� �&כ�RA��E��Øj�0	H��I�@�d`�U۵��Dy��g�ҮpYUF�Ai����5��+]#���o��`��F�(+�@������*X��&w�����Ƒ
����k��7� |A�� z-֠3�P�lñx�6���s��Z������uV0���ӫ�^���2���ڕ���a�6 H||�Ҵ{e���IK����S������=�$iZW��L֚�n$�ح��;#н,�S�X���Q�B�����	Hf���'v@{���ռ���樓q���h�{:4���u��l	IK�ا&SL����QҾF��g4	����z]�)�K�2�s%�-l�H��ρd	����[�k�����3a����z�	8F�cN����..�+|�|�g�ڜ���/���b-�1\��c*�s��C��"0pҔ�vqKkΆIel�!�W��W�	��gz\k'P:]|�*^'l,f���Dd�l��)�a�}��k]��~� l�Q2�8� Se����hE�ǀ��Xn9=�W�������,�K����6AL#��NO��`�C����zaF��~D>B�/���J���h��2�b�s��k,W�p��>z���	��1����4�Pb|�*���M�o1�}�ђ�xo��R�xݦ)؟G(h��$��tE)RY91lj'&�:�@�2�1����=��q�dF	�v��.�p ��M��7���hk�M��2׃�j��T)�Ir#��2��4�c�D,����u����T�k_"Aq[<E�Ƽ=��� !I[�7~�B|�Hӳ�����!*��Tmr�ݶ.Z7p�,iD��gh��&��Wi�; 6���" "��( ��»7��o=Ҕmn�<�s�?'37�8㳈Û���>-�!����2����f��!���q��l!;����@6���u���־6�%��fc�Z_���D�۵{:3�s��+�R�?]smaqZFٌ��;�mUÜ�����B賽�"���u�����B/r�k�����l�3�l���ʄD�10�srkεҿM�#;�ϸV$)񹦳N_k�|0�S���u!�Ie2
۷٬IL6:O��B�¨��}f�&�j9G��u�/:�<�}q�0����p*쩵�����X#�ս��Y�~�uWd����Z�{�\:��p�Fw�*(�m&���('�r]Hǝ$F�jN�;�ʍ�����d�K�c��~6�o�^�h��@cQ�JX`���-t���ۧbk�M�:� t��[�ߨS�ì�g��/�/��dี�ŞX�����8���� 4 IvS���=ӽL#���4ِȘ.��V�Ъ�"�хJ��U�v �^|���,IVD1r��E7���E;���f�2Ss���X�#��vloo_ǿ��:+�o����
yż`���T�=I��u�bk-Z��?Y�T�Nu��=z�Z2z�Y ��(w�U�BFN��K%���] ���	��6�YU�`ٰ��.�I�o�j��E2,dv�d<�C�5�{�&S�s�>	N�����b���V�~�	:	�k�yf�{cJ�l���`�)�6�D��e��&�a�oY.Վ,7#�kD΁ɤ�=�i�����Ȇ�{�ۊ:���������@�W�9�+s��-�GA��ǝ�7L��nF�0O$��i���:�Y����*Nd	��sL��>�~�EeiA�]���/\o�zk�t%E��Hxp��ޘ^v����N�$���w�p�!��PRc�_�N\�K!Z�����ţ ���G`��>z-� j��Xo
25`ԁ�����"t�,�,^������m�HSߧ�J�g��t�sA	���5HT�)w����r��KcF��#�zָJ6	��F��&5�s0�����t�T��k�i˃B���}����(sc�c�>���y�aۺD�]�����%���r��ic�ʟ^����+�L*݄��n�3=@}e� [��̈����#�p6e��ez������ �JذxvR#[��n�^���Gu���g���8<����PHx�܇ǱW�[F�YQDO7%0�K�>�4���Tú��A�(�ύ�'� H�ZZ�8�5"jxV�{�'zrj\1'^�&��������	}�����=�`yjQ��~ ��{	Ol3z�ނ��w7��x���Pm]�#ˮ�D���	�$#�	Qˉ^[��5fD���\ؗޢ� m������u?��A�:��9ȏ��vS�5T�TN�1��y̌$�&�x�Y_0�;�Pg���U
�X�D`�XO[�e�;���Fܯ��JV���Ή�y�����T��2J���םE�peDk���c��ul��۶��rd`m%����0ð[Ze���(��R���HOz�M�"K���sg�{/.���N'^�W���]��k#*����S}��M�ib[~pj Х��bQ�u�!�X(4	O���m��Y딭& ]�	R��p��S����K��]g���,;ʈ9�*��s�=*�y�='M�'�h��ֲ$L)�R�m���G�N�:c�a#T��
�M�X�!�6��$A�1O�<M��KE��=��1_���D]��4���뙮��u>�� ���Y�=���Ʋ�q�5!I��ڴ%J`+�2�`�/u?!�����+;��]�rM��(P[�ޮ #�Eq�~�^]�=WԡW�\/$5 ����΁�F�1�)��sp ��ҷEv;`���N�S������[*D��Z� ���5�P1ʴ�t���%��L:s��}!�7�7��u�����m|v�߭��\,u�r ��$��YXs'̙�����,�Y��L&��u&�m:��̱c��L�-�7���ฆ�0	s�=�&�zK��J��|>#����L�K�)���`�� ����{j&R˂�H`!~���2W=��J�XjdQ�4DF���FdR����*ө�3�"�a����9����U%�+"�creN�ʯ�`��y�=�����w�!}n�cו�z�A�>��B? �d�@$dT����9�	�*����<�YId1�iI��Yd�
F�L��\!Ud�o��%|5��X�Hx3q�g�?#�v=���α�X��ĺ��O.� �̞`=���ҕ�D��ڙ�	F���q"}7G���F�RL����J�..��f%*�!+Pk���eOը
i�}��"� u�8��y8+g��B=�lA�x��$x@F(R����iՕhP`֭ �@D��AG)L��4�*�bۄ�~�4&=�;>g�"��
��Wx(��R�� Yy�-ϑ	`��9��#�J�!��O�Ј��Hn��!|u��Vi��ke�l"�gӹ��rk�d1�Y�H�7��/Lo��֜����l�9¿j�APڪ@��E0��{R:���±���Hix�� L" P�h���nd�R�j1�	�h��ޮ��$a�A�1�K��R1"Yu�ź�z(�l�0�yw�{e�)HQd�C�|x'l����d�,���!�*�Aʵ�H���)�E�LZ~���:�I�8XP�Խ�>����j{*z�G�G`�û���l�.��V�Ӻ2l�`HY��7�7�Y\�z�o66W ;��14$kH�}�fH9!hH���2%�{�[��\m�g�H
��==i�D�Q���%�%xB�ϊ�%I�H!Y�Zg6w����5=�)2	�L�Kv/a�3��@j�f�BS�h��V�v}�)�L�h��A"�J�J���`pl0Bτ
��Z�⺸/�Q�fT���w��1�>X���u�TP��!0�뾝d�+u=�cP��nX��b�l��攩s��޽�$%�2��(H��5^r'�$tC�n� �D)kg�H�úTn�x�:O�څ���:%,��؍ j����Ե���|6�$���S{j}��R�2�y��/P�y��(�Z�	:�HL]�Y̗��̈�T*˓��.皑��e�m����=�桅��辮U>��i��}hL��kH�� ú��]%�9Җ��4:� 8�j��V����5�I��e�EQc��R���t��e�7�Ӳ��Z�d�98f45�+B��Je�l���w"�nЯ��N�vE�I� B���=��j�Ys�;���vl�y���Wv���kV�?C$��:Zsrt���<�S�А5o�[&�~N�XA-"aH����Jp-�X�)h�k%Y��a�Ĉ�奁ڳ�,;�iS>���D�����fZcO`�X,�==#}7��ru}��H��#%ē�����0n=���h����憑-ڮ(1s�>K%*��&45��R����f��I���#�j�)�$\�~;d	�1���\���fW��n����m�d�z�1����u	���D����E����K��i&sx��5X�:�K�/uJm��XWfz��,����D<��x��闺&7\|b
��=�Z�$�,5I��֪��	u]�آ����������X.1��v'@��c�H���;�{#jàs�E])��H5� �N�ˌu�������-�d3�Q��5N&#�dw�Dt�=6�bZg]�"�̲�Z'm��tR�/��Zv�=�u��g�.n���^�/^ʻ�rv�m��r�-�&�lo7��ë,ԁ-5HV=����g"ZSH���-�f��ϱ���{`[3�%�G���R$������4 'qE�����"�`��1p�uFV�i7u1�ŋ���˟uf������Hu�B˧��2O�b1)���bc�7�cà6R��v_��w�H �D�u�R�TB߽y�!Le5j���3��B���0X�b����ɦ"&*#U�^��<c�x�R�v��=��A�����bg�g�{��}��� 1�S0�s�as#�E&˯R�$�Ǎhx��N�(M7���ƪ�oӔ2	��K}�����G�� ������4���#��tb��j?���9(�:7R!��|[�s�'�i��A<wȩ�p5�����+�)�J+�7�J<�8�x��&C�(ӭ\���q8}J���)SRQ<�Ϯ?��y���:�pO!cBC'R��䘯���	�8������뛕�jɰL@u��Ŝn�_Y~�U��37�S����Z.�o����&�+��T�M?�g3Rp�A�L�s8�ϵ����҄��d��H���#ɽܐ��tf�b+K�;<<��wt�;� Ui�4�ݩ���U}>��\^1�����ܰغc�P�$�!��� R�$cc*�@BO�a=O�	j6�2XR�<���Bc�����D�y������<
$w��Xm�� ��w�7���S�W9	���l4%���D*}�q�;O1�ݗs<{�D2!ԢE^�m�ZǬ2@}��N��Qץ�ό����ޛ�$�+�ĭ)���d���t YZX�����Dz�<0��:#Ő�:ى��/�m�Jj�V�����}�$���z0���aQ���Pk^��^�=+&:��Zq�h�jȗ��#۔8֧��J�g-���J��=��w�#{�ٙ1� ��>D�;�ik�&˞
�9�~��Y�|�M8�3��^nn�ryz&oN�q@��?��룮j�$�gj��������.,�;ܥ�7�������)�I�ƒuZ&��I��{cMz�� Y �h�4ԛk:ڨ�lj�CK�s����^R@��i���#���j]���cZUy}��ǃ4E�*8��¾�yUnz�������j(���$�2b�Ѭ��#��%��1���}�-`J�X-�D��um�7��A����	��1����=љ�3�܏��и, ���`_\^\r���{�m8nwOn"��MV0_��Ret]"B�|T2���t.��,QB3&d�w��� �����t�l^s����i8��cK��f��d-�x�)u���c�1���T�������6�fZt�y�M45�GA����+Β�I���M�=1����s�'�;:S%�r�:��٥|��K��_��/�迭�n��X7��jEτ�V>��ۃ�F��t��Z���@���j�yt^�3D�L�:D��o��!ԩ�LEW#�8c#�G�W��H-
�fE��
6�kt)�s�OtvJ[d*o��oM��FJ	�T)�6�5%U�x\@�$�1�($kT7ƍ[�%��hl��S���� 	�*W4C�C���%���N]������.:��o>�f���t|m ����0�,L�D��4�1�
Rr�,���Yl�����0"�]�Ec�j 1Q?D��X�4��2÷ՙo�˳�̧4�m8A������G~t�)� �e��X��vUt��k8��)C�Zԧ���*�p���Se�� �}ldt��b�ɴ]�5.��F{p ӣ(dۍ��)N��ac���%w���@��78<l^��F��*:�=U�}�P���T��,S�Zy����{�t��DnV�d��a�d���=�=!��pw.��ߑ������G��P`ݽ;�7���/���S:ȫ�h�~�Ƣ�3�ֆGz�D��K'�}�&9G�� ���$y�i����#Ll�U�e��O�����ݥ\.�$&0F���ۧ��������K}��͛wL�BvER# L� F�_O�NR���bZf�k�Z�	��2/�1��J"J�r	i��׵X.WL���Z0��iD9M� b�z�o)�f�'wsn��|�@�����,��G纁z��\ߙݠ�ځ�9.�����G:t��*�����A�7Sq��v�bցg������kѤ�}R;����d��-u+���&�ڸ�U�r+�@�۝�1B�N�=�ʌA��C�GiB�H�=��"u+7�����d�<0�X������t>4�R�DVR������Od���<���4e$
�'�f�Z׽���5� �^�����2!D�9g�dSD�֯�������$'���U�Zs
@wT!��B��[ɇ�֎"u�������5��n���O�F�X����ق���]�z�k�و�w�`#Cs�\���c��G�l�>Y�tc��,�����"Y!S�qx��h�a� ,����A�����>� 0��H4����s�wĕҐ����fD��>ZG�T���u��BFӃݑ=��}_H�ךͦ�ҷN|H���6�����)؈j�P�e�hL���g���4#}T�'h|�qg��	ÿ��7�[����F��3��y!�wx�6Q�둸fЁ�ϵ�%�n9�ǣ0�oLg���ұr+�l�9�#�j�E;B �ތ,=q,��&2��ұ�xO����;������ޡ ��D��2�7�������ݏ���9r�g|��>n4�y�F���ϣ(y �cE�2U�<�"����t �~�:4�� �f�G����L~�q�E����e�8��� �JqejD
���E��ݦ	B��(����Svͪ�@lC��MƑ���cr��^E�!l[*�5:#Z��(D�����x�^��/�pP@/��Z'Y W�@B��F14�z9�@�M2E=Ȓ}UNBj_ϊ@'��IT��_̸vb�`�,c�P~����c��2��!�҆G]�kaS�;��r�@�F��T�_d8!/D�w��X���-�<���Q��@���F.w�J*�Ĺ�z&'X�ƅ�8�ޡax����(�y��<�C�GJ눴��2�ﻁ(GS�����p�>��R���{%-]a�U�E�jw����s�kA��Ǐȝ���%C�D�W>y~&_}󍜼;���
6LS��-ݶ���H�ܝ������W�4���L���k�G�7��rrr*���/��b)Hk�)#!��,X�E�V��K���WV�U�x%!�-%���&{�ʺ=�Xհ������<{�X�=�˚��|�z(��`��NX?��=�^�ʫ7o����_��o�gÀ����!�
�٠�qm6歬͞`ݖ�ݒω����]A=�5�1вX�
C�'�mmX'�y�Hr�g����$��b{�ZZ���G�A�Pʽ��Fi�]ou�]�UnlXM�(��:*Yv��at�D�˂5�����C��0��6�o�h��)�b���d��Gg�`%��i[�ފi��:&�V���A��X�c �K$�N�G��8���z�#�r���Z�_x�[�F�R��\h��ca�6i_�ޓǏ�ѓǲ� w�����]����ӱ]_uru��Ԗ�7�?V�x�_/��S�4���mwv�$WJ�nV:����}�^���9=?7XY�A*$�t�P�YZaK�����w.MV���z�ѵ�0�֕h&����2��I�:��0���+�E6�i,S�(�S�ű�D�Q�u�X��d/Y�S�g�{�3�������9PrDS�<r�C�5�{��l�3�eoX֒Gӹ��n��:Gk��S��j#���4�l�m<���cjbt0���k�
a��m�B͑��q�V��	}���_`
w�4u8b#:o8"����'`p�4���7�lj1���z"Q�����ױbάOR�a��Nk�AqAK�t��-gs�6�*�NХ��ۢ��6�xt�Kg���#�L{�=�����V��׺�/U\oP�a�=}:���F�����뭿G���2|c�k:�sg��,�Y���@�̻��g]�"��HO_nT�b[��/C�,"2&)�J[Қ~��^ ���K�L�,?������4�%9nλ�^�mL`��6T!�^��,2���hsm�&M�&���B퇭X<@�I��c�#������f�쾕y�Ҳ0��e�q���d���a�vyH[���X���0"$�EJ4��J�+�=�*u�h�܁���g��J��ʀ�(�O<�+��`h7��Y5��aʻ%��iS�đ78��"�����s{�[o3]��p��@~d�G����C��q�u�ޮ��Rw��gW6����(E1>�ī�$�D��ƥ�._}�1���>�8`ة��Gw��\��J���SwW�Ffg3v����+������E�Ux�P��L��Yׅ���J�w&�3G3�'�h�=��<���)�Z�Zu���������5�jf��ڥ9	]1�R�8��;�!H;��Gq7����&֠#R��wi;�^���������GQ���Vɜz��H�x~��$��(�Ł�A]c������FEz�u��ܬ����5vr��=����+y��9�:�g;#�"�K)����#�$#� ��[�䆹��>X��foj�J竪q6��,���2�*����9J�ю9���Z��Kѭ=-�S��1�� ���~g� ��=ѹ��5�[ZV��W�dk��WLQ4ǒ�y�C4+;GAj
{0&Daqn\�Xj����ݶ�}��$-,���洎uUA���o�4Ǩ\i�@x���,�.���Ys$;{����GJ�>��c%X;;�0
�F?�W�uyu#g7�HTY��r)�X�C����rg��e)�V����{��U��J�wvyn2C���3�p�ys �]� UCw<?`���s ��ƎuD��/��KkyO[��-MI"MS<q�}HGi!����a����;���ΊȽ��t/�� S!����s��>a�_S�����5�_X~ ����!��t�5��YP$АȏWq��c���N)��"�*:��ɜ���w%�c5ȃ��)v�ܛ��<��g�t���`����x�L��m����증�gN��ӿ�)D��%n�#��ě�uv:���^��p���1Dǲ�-��J��R;A����e+�hy������#��$�|��� ����1}�� �g!tH�sg�ǎ#`zsekM�!F�_X��ĳ)�ܨ�ͬ��^Z)���
r�0]k"���#zU�ɂ*?����Ɋ[�CK��^F7V�Y�[;RW���B�M�Ж�� ����DA @I�E��Q�OQ�����H�)��A�aoS�5X����WD7��|��
��� �����q�l��L6��d�R���=�F9����ps�y��pt����c�������jdh�Z�r�P�� �kt��R4��-�8X��M�Z����	B�i����
��&��(Ma۠�����E����?��U��1�w�?�C�9�ͽ!U��_[�q�E�07y���떷7��}x��hkx���R瘬YI���F�(W}��ܫ��v��- $��<
W�$�!>w�D�$*�2t��{$����s᷍J8/��X��k\�!2DU�s�Z�؛�\�v��=�@�ù�M�#݅��@�{{�'-mdo��_]_�ۓ�rvv��k��9k����kF<�10};#H���II�²�nbg�CB�^�r~v�&+�IV@h�"��#���US�w�
�䩻d��X#�$��E��!��N2ݡ�� �c�;�[�,oNN����ՕKy���<|xO?���)�@E�.;Sie휑�:Al�"��]�m�#��3�gEyjH[[i :���ή<x�P>��W���Oyß^��/���,��A���Ү{;��#WHC�4� ƺ�u����vei�USGV���W������+t����{GPk-^3FJ�)��|g5f��H弿��g~	F�?�6��l����A�LA�>�@JY��u�,e��#���s5�A���d�~�[<F�@��H��xK�늻q8�hp�������"5��G)�q�H��?��UaԐ���$S`��Z�!��m#i��5�Fgւ����O?�'O?���9��{W�"Z���L^��I~|�VA׆]�К���b�v=|�������ɖ.�������#�Ƿ_˛�'�F��:OS�Ȣզ b۷��Y":�A�6`u�����.�L�2o�T��9H��;4��Z�Sb3oT���֮�:�z���r1)l��2��*����%:ej "����TH����%
��v�N�$&Eڥ��G`�ث��R�����d�Yu��'��z$�ϊUx�M��T��/��T�tAۥ�֚LC�Fc�d�ds"�&C���!�q�Xo8)���Y���-�k��lb`9��>�@��W^׏����Eo+�&H	��;�m����.<�:)��C�[�XĴ4��-M%���A�e-�ӹ��5v��ͣծ2K)�Y��r�P�7�I�`�0F�<��N��2a�[w���72)�|��p�����HSD��Y�Xd�:�RѬrӭ�<Z��x�<֖&cBA�����u#��C�ۧ��)/K�ѲF�[�a�]��x⑩H����>*�Ô7O���a�Ѭ7}4�5��"ׅ����mj��@���B��;̅�$��56����X��5R��]�1�F����Z���iʣy ��u���6�!1E�.Pr�a9p��=���$/H��  1�=^�A/�b�O�P�D����9�u[�6�/1���*7���٪�b�%�9�b�{���x�����3��F���c�(�L#Ńy2�TBJ�	�����6���`�
�������Ÿ�ѓ�/�X׻f x|n�t����P��f����R�:����J���x
kG�^�X�G-�j�/��i0���)
�'���GA��gK�+�>�/�U"�z@�hܹt@�N�B�����#7�/k�Qz9��~�׋�3N�������q�ߤP��O<,S"%��������aduAon?�I�fS5�s�+��ћ�L��c�s�H�
4ή�@��P߷PW�Q0v؂�ݵ�]�����=9�w(����2
ۼ��,��2�I��Xmd����s�Hf�KU�͊�k?�ke��J��<���z��*3j����q��P`K��1�0OUb��ɫӷ���/�����O����9:��ݻ�L�ژ��R���tG��Ρߗ�s�͡T�=v�����,�0�h xa� �l��^�o�h�H>~�����N��o��J���������)]o�s06�6W�Ԛ	��΍��\{$�2�`]�
;O�sO��f+���M1B�[�Ա
�J�.ȩ�zA�,N� �3�*w�Y�\���]�=��DezBr���@�����z/�Gj�bg!�Ǉr_e��,�_����� ���"� �w���Κ^����i���m��=��7bw14���T�԰�?��zgJ�x�;�Y�Ԕ�M��`�w:�[7Lz�Y�'l����E��7�E{1�م0�BDvL* 7""V�cz�G��,ekvAm�h��@w�ʝG�d�h��7�5�"7JX�]��W�'�����/߱Ex�i�0��9>�#/NNe�{���/d�P���T�Zefq����W�^�d��L�.�2��6x�	�82 洩}2����!��uF��=�h�{���p��j����N,0W�.G��xY�}^t��9���>C���~����w����{g��W�L�rq�����8��? �����V���s W�Mo6� }1�a������aP�6����b�:s�����kA�
�k��l��5��Z��,�u\s6�!�Le`��C��[����uN��s�{8��\V:<��e0}g���~��<�-��~�U�m��±�yy��kh��V<��R'��5�{��õ��g�!F�qlǦ���>�����/�[h3�yR���or�X��%�NMH�ʀ�r���>��:dGl����9���b/OѼ.YԖu�8Ƨ��k��,�*������HT�H����V��#+�8iGZĎ�T�����<���XwƮBc��w�r�6�3/�<����B,�z��J�ElU�C] S���\Y�$+�'����0jy������N�3��0�x�;���-���� m�/']�4��	ue�ʣnL"�$����	,Q���0��Iȣu�p&Li	�q��Hð���1V|)���0H��ę.���#~��]f�?ad���� ���:���in�#���i�u��v�D"��Q��s*h���"P}2�5*{�b9a(ڌ.s8���C�v��@�IL��������r5��a���8�����į @�Eb�k���㰴�h����7M�C������\"G�t��CG�q5��kx��N�����2�."��~�Ӑ+���r�)!g9������,1����[��ɨ~�
�vx�<W�w���j RC�G����/�h��O#=�N��Z��PLT������`ڵ��iP������Oxs�7<�q�����ٍ�+$v�<�LYS(��LK�?8��[3�v��r~q� 劎/4t���'H���:��=���+;x{M�bQ����_j5�)-l�s��w��!��F�u"����w1C�s|&S�^(�<?���J��y���>��M�n]MK�#�/�^ۙ>K3]�����f��4����������4~8G�ѣ{����J���?ʿ�_���]��9��~����ˮs;61�~5��LVЛ�_�9\<29�sw���2�����$������0i��[��Z����ᗖ�inQ��W�H֫�荂6�	f�:�V�f�����0M��%��6ܹ����"X�g3�������S��q�jek���GA6��u=��{��n�\vp@o����_)���`�d�g��S���l�S����>�d�A��5r�w�b�QC�6�[��i}F��1�^��@��{��*2�a��.~�hW��k;iMK%�+�8���_� ��K��_���|����Ӊ��T�~v�{z��_�Dh���gO)� �77��Z���%�
��G
̙�֗�f��c�o�"���9Stֆ�!����R.W7r��#��gv�6�֩�OL��2j�yݰ�e>kd�~�G<�aN[:o"%x�����Grxp��{zv��CM�ңm�5�;'٢>A�j�V3��~�C���PGK���ct ��e�bs�)e��c�I����ruqi7I���Xv\�&&�%pJy��wvt ����>��}nG�`�&v�%��CV]���� ��f���^��F�l��9��.Ku�dQ�H;�Y�]�z����1e�3���cJ&v�0�@���'�}pg�)�7�V��\�q�2�QX=<�����,�;hoa&b;�0��|����*W����|C�lUtJ��}��x��>D�G�񁨱�7��.����,$�Pdg���j�F����Yoc���d���o�.����t#l�W;��xp$P�����r�a$�0�7���<3.��`�'[�;w4(���Й���R����y����@��6���v�G��y���5 hL�:��~�>���J9 `!Y����wZOJt�^��vmW<�*��CX%��/�;"�c ������8�rpmc�ƾ������ ����u�m����S*a�ډqɧ��� u�%��4���e��(�b�(��4��i��S��+���m,�%Yg�(|�R.������J���Z�Ax���!:��YO��*�Vc K��AȘ+���b�S#�c2����o7?��x1�H�x�U4�H&VRE��aM+��ީ)
<�DykR��v�(i �U���%R��Z_�
�-�sh�zo��E��)�}��}rCٖ녂�h�[���q_2�6�47��	��Fd-��kU�g�;�%�1�Iְo�Hԑ��o$�GN�<4$����r~~!g���sWA���,ņ^ԝ]�^��>�����m0n��pǄ��;r��C%	��lU�Z�0�=y'/_�b$d�
ʺTY���9��z�5u��u ��X���/RW./���� 0�������A�¼�s⾨�w�꺓w�O�͛7Jl�队��oS�\�lO]����� O �ZC�r49 �a�����٬x蟵5G$dޱ��ǟ<������_x:�<{�@>zz_�����e����tK��RE��ĢT,��������R�ը9�������-x~<�7�K���4e��$k��ưq����h_nְכN=���y���Lm:٥��"Z�tU�;��bCF���:ef�ଟ�����F�P��\a�t�7K��->V����&<�5�l ��ݙ��֝����Q@������������+�sbj �8L�^k�{��-�-k]�d�9A�:!�<g��^���f���v�gg$������Z��$IyO*O=������0��͵�~w"w�Z�iv�d������/����_��Z��ᅼ;����INYo����g-un_�y'ӿ|�Ը�Wtf]_��<A�·o��޾$��"�PM�eI�yÚcÞF�g�����#2��\�9���w��u}OTg������%�#��j�����i�a�b 2^y�"�����{��ﲣ�t>%��`!j����ߓ�����ށꓥ�|5�Cr�cE�\^ܰ�8jV?l,	���K�T[z0�@�{�*�;<�#a�T�����b��Ip���\^\��7'J��,�'�,��̸U�q�������;���\[�V�2�x�f�D�����stH�Ǿ�ٝ�9w3��ԵCD���Rn����j/��\��s_�ry�sp�d�������ñ3!�j�L�Νs�w��g<�
������F��N�fM�����y��X�=ƌ����}ϥ^��~A��3��g��ݕ���&E-޶�8��I�;&�� �0Lӫ̱O%��v�|��1B� Q���;��rdK2'�Lo��X�]��2[z%k��B�w�L;�.�u-�KZ�a';Gփt#�����x S�>j<���l��=��Xuj����B����+K#陇ٽ�]�4&�pK�Q����w Z1z�b)<����=G)uq�9}e'4�2�E:Æ9R� F7�P�I�P�(ܧ.�"����R�N_D`�-�?|; �W��oR���V�4�%0 �2����!H���F�8�h\4H]��m��s�h-o��ҭ��r_x�D$`xm�5%�����,ŀs^E�Q�q�gzZP���OP�ʽ�����;mE0���,���MA�[�̾�B���{��`F|�Y���yaQ_E%kYQ�ɟ��&q�9u��9u�+-X��m��Y�Xx�x0o�]�<+WՋÃ`�Ϩ�)�
"1I�H������
��_�H�~ʂR1�Ld�̵gN���[�i�d������̾����ż�Ö��6!�7![�S��s0���[Goy��d�#3� ��HS5v�����W{�3e���@E���ݽC98����Z^�k� v�}���z��ʟ��j����3�J��|+ ���f ��*���%��Q����;F}��V< ��](��-��:�����ӣ:�;a*�R�)�{���\����Ts� \�()���7�0���u]���ճ����ƙuw�����s7Sy��<W�ut�K�ho[�������=���Hί�t��{��J�ֲ���Q:A7?tKg{�;�Hi�g������=y��<xpW�"�x������@�����~A���z���
��<���siFw=ը�V�j�D���|���Ƚ�{z��
x�|�c <�  ���[9=��7v5:8��`oJ}�&#�b���~��ߧXkf
���PԗVQh����z;��<�$Gwv��h�]��EcAZ,j�ޝ���^��Be �{Φ;
�j9y�����/�I�&̠���� �n�mwm�����,a-�W��G5��9@����Wnv��TE/�t��^^�듷���A4"�Hc{q&���|��7��w?(�z/+�Y�|(#�tޡ���Gs����╬�W2���a�����8/���Q=D����$�-Vp�AoN��s��ܻwW��ﰥ4�'����=�w� �MR }%�'
���r�<`�Ӎ�w'�����t��S)d]�tDz�Nf��O���u�(�9�nA�Y�	~wv�z�����c��rY��4��C��ְ'''�мU�s���BV�g�'6�h����sf�x�Q�u��꣏�˓'����#9�������>�q�l1-��$��J����B�tޜ�gE��]��F Z�ߜ��Ǘ:/�r��P챲���JX2�����g'�O?�D���q��y(����7+8�T�����w����R�J�^�P���ky�sqq�bd��M8��,3'�L���h_��y��^i�K9}��x%?�x��?1ҸG��ۓOU/�淟ɽ�wU�����H����e������Oo%��k:
q <y�|�^t�Tt��F8�(�fQ"�=���\���5�2���J'<.��z5����v:��ǆ��١<۱f�|dBu�@B�CFg7J�,��
��6I��N�M��8��V?g9�m�>�d�f��bB��੃LU0�a�����W���=zzJ��Q���d+�.YPf���׌T�$Nޢ[�M��h����e���z�� �B'���q�:.���v����!{��h����n�%��#cf*@|.鑖��F�[���GB;D�JL���PQ���:�k8�Bܰx:�����g0�n b ~l��k�.�{�����ɗ5���qc��~udFfᵢt����A��rmDὰ�z;���_�N�VY�v Ȗm[��+(r�K�Q�BI�1F�Bܾ���O)t�GSEa�7����+�~�c��$��7m�Xl�ۨe9�6��W�
"{jL�F!�٬gIa�W�$E���5V̟F]Ҭ)�L��˕��H��e�$�����)iY��[vF� �����U��J���4��������.(����×��z#���J��${m(�
���^���T~��'
�����k�0wo�Ōq�쬬����.�.�g�����9��z�TB<8R�6�����y{�$����ZY>�a�����gJ�Ը+y�`쐭�-@ti] Ch� ��T����M����7�	��Y'�?��4-=�-T���x��oⵂ��''
&�z
���u�
���>h�q����%Z+���k+ �)MCP�no�>�t!��C4�_���<���<>>��w�o���8N��ߗ?��g<��B��\	��O?����%S���sؙbR:vn��*�=�h R�>�����7�ȧ�}"O�=�g���T�(xр.�!��O�f��ݹ|��w�����^�����MӅ���F��/H/���l�>���F�<|"�<} ����X�\p���ں_�x�'/^�P��8���X���IgH�Zлr��W_ɾ�7of�m�n�́� )���*����f�}������|,?���S��m-
&O��<~yHy@
:�`>��y���o������]|���|g_Ƕ˨���X���s���K��Gv
3)�jƇH�;��)뀬��ˤ���M<�c_5�*����~���^����S���HnK�I"�k���^�~���T��P{J$u�t/�&�~�h�OJl���� b �k��.��#�w�ۄ�Vy]ޱ�$Ϟ=���� ��}^�c� N���N�����x�i���:�o��/޾�����J���nk8��q�@���ټ�now��dH�BT��ΕX�M=R��ݷ7��ֲ�����}%f3Ց�J��	�O޾����k������˳�JHnH��%S�Pȳ��p Μ{������o��L	�G���1��"�4��3�S{�.T#d��z_�ݱC��,I�ԅswJg��K}��K�P����_�ܯxx��k{�I�h�4��+�<}(�����GG쮺Gg���{���38 6�^�wW���NЉ�����/�ȗ�^�z+o�Θ���_`T�7D���4= ��ݯ���?ᳮ�W���/�?tmo���8��=�k}�_�ꉾ�S�կ?&)�[D��2�>�7t ���W?0�����Ҏ�`c���Ȝq���f�|�-�{�di�9����Tl/�I40�4l��#YmN�� �g��6v��jE'���Ӭ�+��qSY�Q;%ñ5�Y�N��-�,тs,�1<Z����6mc�i�j��)m�OMr�mX9[�>;�8_�p|5	�j��!y�J�����)��+>x�J�{k�Q�u���{=�Ȑ3]�?�+E(��)Q��_���kH��4y�2���k-ԧ�C�xx�88�m���N���tNUy������؁78 �Z�䭳;Π��0ÿ}Be W%Z�d����+���g�YC�ո�����X�X�BW3pvm��x�~T���A�1T#^}�-^�@f��w���C���sl17%]${��<��4�R�BלmR)�#R+�R��F��Ȃ�.��������MԺ�������\��.gq�hP������[���_]'�8|�X~������qAAE]L=JA��FU--��Yδ�^���M�Ѷ�"��KdBGG/z�<����9�&Y{�W���Ĕ�]���-6��C2�k�0) �U��+r�Vd��j�a8'D����8�<���@�P�uyy!��LyA:���B�H��ϵ��
���ѥ��ҨC7�KX�CK7j�8��^ɻ��D\�ݗ=�C�7��8CѠĚ��s��a� ����?�/�����g
�i�� p!�4�!��)�o޾WC���Yv$Y��.��;��7���{fʃ2�|C�`ެ���g����)Id�_�c�lH�����&xށ|5$Y-��$t��b�:�)P[�z/�o�)ƙE�|�����ik<�
��^���| Ȟ�T<~��x�^���AD���hj�iēa�	�(��5���H�v�>H�'��\>��?z4�H_^�(�ە��{L�`D��&_�|-���shþ�a�S��9��Y���w�k�R`� ��]��˿����ӏ���]q-�8�c��l��΅�́�;���A��.������k�����û�BI�o���6�e�\�M6�\��&��S O?���G����J~�ґf�G�s�6��n�={*��H{�߿ù@�u�U�<��ɻ3H}�1���;0�_���c�K]T�y��5�%� lD�z����I�@Y�h�v_������W��#��B:*RWAbpF������U�Q��յ�7�y�bm<�H��z�{��9�A�';��D�;R�@�q/6�@+~F����/wq���J2>e'OD�vTVJf�8�&�ҵ+�Ҟ���H��)Yp� �5A���\ޟ��a���g�_t��N�|���ɑ���'���>����r� ��x�K�ab��v�����������w���OD�.�u��
��,�8<\��|i��6Wl a��vl��̿���/T�>����K`G�T����s����ߵ�ddZO�	��#sB
���>z,��kݯ˛F��;��$����)���|���W�2j>�#�����@,ʨ�KH'ߟ)6>�tH��O�G��������w/��ﾗ��NO�*{k��A�w�#��D��~���)�<�n�t�d%���ߙq�?z�L����ٯ>�G:?p��y�zt�k����Yf:�Q�������R���E큍������ '��Ą���:;FC�Ȉ1gqc�ٔ)��1���3� ��8S��)8�ܱ���voxHqσ���/X�f;��ӏX�`�+D��_��;���V����b�M'F�,�Ϻ�#�f;�ڎ}�zw�͵$ݿ�q��fK���x8�*� ��hypl�'Qo����s�Ar*i~�k��Ҧ�\�h_ι�݃e(`���׽�$��ӹy�;	��Y��`7J;ߨ���	âֺ�Z���l2WH��6�B:ۄmQ�v*����Q�H���hl��5�܊LE����Oe����`�4Dk��e�ء�p1ƷE0JT�C���ϊ�S�b��m��9����!�Ԓ�{�q�Gl�R�бF,7������8.�M�V������d2��M�g.!`����9A�1��Q���|c�6����/v�La��5EM��6gHQ�w=��DXRL�F� �@�=�>�G��?2<GW"Pɣ2�g�8<x��E�A���0�].F�1'81���%�r�h�B�����v�6������R��P���ĳ��.Q���G����*�W�T�"¦����R�5h O;<Rz+�u����"X#��us4Ei�x{k�띣H+�&�6�e΢�9�h�Lg��ry����]ZJXۛ��������� ����L'}�A����W'�����j����A��; w�_ۚ/W���+�`�1�T����7�?�N>�����l�s��,��g�Y�׌���|�1�uzv!��ߪ\�P�0�&Woau3l�LDgʄ���+͕y�2�Je54�t�Q�\��հ�	=��Be�2��/����\���]e�F��̈>_A����Ã�T3�[D�&�Ou}��X��߰U�	�����=��9�s�������?���?����+���G:�s�4�TA֑���������7�Y�weg���w8�u9�o��A�S`��j�I�����gp�����Q�tW�����_�����TAٽ�s8O ��q��(��]�1R� �3�y� ��u-�	��|B�~��������߿7�c�6����\e������'�o~����w�˓���33	?&l�		�>ǡ�ό����O�==yxOI��؝�G���߿����7�)wJ�f����c��8H�mlA)C4�Y7��<v~.�Z+����� �t̙��x6��Zë���N�NO�8ܛ���>��x��>����S���N��l>۬z��I�$�?���F����`�X#�Y@� �b6Qb���ޑ<zpO	�#����L���h��f�ؘ9k��ِ	Rg�4�H3t�*�3�|�gUD�Wz������L';{��Γ��#{;���G��_��$3PL�5�-�$�x�x ��7A�&�TM���s
l[�F<J8���ן?��6����g?��{%?��J^�|�s~�5D��O�)�z&_(�����ӏ�3}�(�!:�^�_��Պvbo��3�����Jv���l��h�r��w��z"O��X~x�:�k%��݈�<zxG�={�H�'�<#��S�8׉Fg���Zg�iy�L�J��Zc�bH��=%������'���G�����_�L����t�n��:G��T�*�>d/ ��F��X��7J�v�[�3˱���{Ǻ?���ʘ��}�3��}f࠺���ɑ���'��)Bm\�j���\�n�³�:sN�w�g�a�C/�f�w�l#8L�gP�
��xG�:G�V`����J�n�/���./����w�?Q�3%�e�uSԔ�z���yF2�nϦ�$Cf�72zx�^��9b�����9��/<rU��ʧ)y�������j,��n�(D8�m-���E�J2�t0�#�R��82�5��_�b�V��H��ԃQw�8$�G���o������ �`4[�|�"x[�s���}�*�0��P���ut󓷙�2��ZMm�X����#h� =��r��u$�X���&YJ�_ D4��Ϊ�D�\@,����指
�����<yKo����5���Řؙ�f7��:[,^�>�3����Ľ�eg�عg� ���Qc�4���1ԾFh$D��v�P����yh� Y@����g܇��[;�xS�އT������χȖn�m\A�H��F�mjk#G��3�1� �����1���<�6_0��<¬��>��(A.���3�J�0Ǎ�ɎY0R�`Q2u��t��]n��r��ᨹ����%�$�H&;�."��7i|���]�B"-��A3�)�8�Һ�D
,���ժpM�YKDxhgom�Q��&�ѻ�ڽ:��s,���v�"�����=HT��}�Ƅؼۦ|�\��:���r�Ho)�C�皨a�{|W��]z|1�(~�S`���%���U� ���r����n���;�]^ޓ�����[�>E,�׌��v J p������	���g���UFQd+Sc7�k6�0c��%x�
�',�7G�ru������}��������FCz]��Іr�������"�	N|t�;ؑ;
������Յu��օS<�À/�\-k�Pp^Ցڛ؍��|��8�]��NAf���k3;m�5H�C��g*��'�8 Ҩ�� k��)��xﺉ���O쨆�ԏ=��8R=�H��V/�Lҽ;�����+�S�mVrW��'���T:oY�Ĉ<�HO�1� ��`W>S@���-��/��_=�;w���8Ev�p���Z����>A\rߞٍL0���<�P���h�[���O��䅥��8��?Ps���?�?������'ϟ�׽���x�ioځ���Ab2G�k|�O�꾹�?�˗_�Hߙ.�Ņ�U��<��>�G�l�ؓ��%R?�4��w�y!^�)���(0���)*�;u2qt�AD���Wr����ZrdG���J-JKh���4�ͼs����p�l�(��Z�xn�~���O�U����us77�?��n�%�{Xϟ>��1�D�@uE
t����R��x��K�WT�g���͖	C�TnP�9��b|�(��᡼y�L^jb0!�}M�ё�y !��l�I)��P 1 4�k��ڬ5�=��PmU
g��ލt����4vM��9k���������K9�u?CA�p�")~�����r?�f|�$2���vv�uZ��M���ݞז�y��������!��H�7<���w��� ?��Gy��y��X�y��S�)P�p8�O��r7�L:�{����. �b˙kt��Tc�d:ѿg<�:�mM3�u���%c�@}�E�?+��{����^��7aLaT�L�hWm�1@_�Vz��<���k�y�hed��c�L�r�!���rx� i[�����f���9;}]��bΏ����^��߫��vP��ya�T&O�%NaG!lMv�U�yV�-uХ�f���W,��l�!�[7�7D ��l[��ɒJ�����f"A��#'pВz.��E}�+�@9�7�����ٴd��	�1gN��<6��5Oحb.eE'愈�N��?�.����YX����͕[��8	�#�R:`%�s�Ȼr)�ɢl�CZң<:YT�P	Y݇8(����+��c0�Y�$� T���5Z8��g���S��`� 0nV�i8���%�PA��(�E���%<��c�r�d �8��V�Frm]T�r1����"�E&?jU㬒&��N�`��ܫ��%���)�ě���!<���n�mEdnҡ�̜�#�*��q���u�4a�@���b�NB�(�4&�It;�BB�V�n�V[W[�!7���k��Z���5�!� �	^; 9k�P�|�a���m�0�f��@ �NN��"h�q
*�1*�=&����9�T?�L�+>(�� ��l��u��D6`��Éo������$HE��b �1���8�Lx��"-�<���p���k&b����H��Q��ˤ��ǽ�b��R9�iK�*�$������ ��
]�hB�?�Ӥ��Pכ�R���%~G|�BQ��M�&˼��&oE�2)i~�{��M���KO� 7�۲��s�:��0i1�u& ֑AB���%�pnE��c#.�nwQ�"0r�"��!GAR�G���/� ,�K�E�a,��dE"�`Q�"!�n�j�L��� ܽ�}?u~��|��݉����#�@V䉟��ֽ����n�@��S.ޓCt���2���
ݜ�ݮ�������W����i"rD�!��r�3�[.�Dc��B)�^�o���U�z� �9}�#O����y_C��-8#�y�7��K�aƃo�*I�D'���fh���j��&;;ݸ�'\7	�
�c���7Zh��� e��	z���z�u�h�ѬyU4%%��.(b�B��Pc���T>��(�g2P Z}yH���F�?qd4�u��P�qy����>N�	��:W`���Dvw��p���t9gx�lTC���~Oz
lzH�4 q��v���Ɛ�,������ʓ'�
�����o����}V�Am�|�Ro�"����jLv��D-��y�/>`'u�ܠhYo��{��*x�Z�з~n����S��&��ˏ�lq,��/��z͋�� V=c|	� kRl�������di"�$�������"i�C858����
��8�r<��c�}��myEޱB8,�ƞ0Y�a�����h� �����r���HNK�G���N��`�k��Q�[ ��7(�/�gH£ʊ�q�@ʥ�Kpw��;"�Ȋ���)g'ѹz� @k_�f.��`]k1����5�:x߽�CJ��w[�"�<Ȇp�u��� ��7��tl���ܡ����˹��.�H�;�������MDs�e�!��AF�/*�iaZ �v&����g,�i;���VG�E�׏"B�֔-]��
.�]���?��~�����P������?*p:М ��i���u?�}������{���� �f�T�&O�P��Ç�|��vv~&�77\;�������~��{�q�:�:>ړi�������t��BJ{�����'[b��u�h���s�l�==�8�k�j)����*��v&ݭ��P�/�Ӈ�\_^����8;S�-�u�q��@����ּ�D�� ���AJX��B"�3h��7ry}'�يs�&2Qg�fl��f��̰kd�����6��b���9� ��{�{S瞏��>C|M���*���&����;�Ma7�D���z�
�K�n9)kI2��9�.�G�3����~�'�V�
3�։��	���y3���:�
H$�9���d��]�z����V���{�ʱŧ� V�[�%-�e�ɾ�C ��ϡ�Xw�ӀPP5DKKҸ���eO�WD�vs�0G�^��A2��>��屧N�C/�:X�`3����ht2�(gY�����A\濓��TܤX8�̧?�B��(�D�]�҄X,�6��F �D'�p�x���D��&�B��ϝ�jY�G�1���;�i� úQ�Iу��mN�KS�אzE@���t4��� �`A4b� ����'E�D�* Pi�n���EU���ڠ%�6C	�|*4���\.���͖t5a�B%]�je`��r k~/x���Y�z�7�4�2�n��D��z%�y��4�K$,�<k�wF�*�XӠq��3��h&h\u>��Z�\�uH�v��Q�,9�o�֥�����V����
�&�W�{���֫��|�����y�}�V�y��4���QVV��8�\���5�|��+��� hU����)�����'} �S��uO��b`]�&;�
>7�\�6�|�hi���bPP��wY��%���D�[A���D.�����.�x�*p������+vʠ������ _�!�V��
��ho�NWv4	��=@ER��S]5Q�C37x�U������*3t��s2f��,���DXY=��qN�5���ѡ�z�D^�:U��Z�>9`���1�P�XA��A�9Tmq1��4#x����RL�1#���IJ ���[�ΗT:�@�a�D��.zm Zsr�!�0��ڛ�)����\O9����̅ᏤI[���c��I"�K��Ϣ����r� ���3^�r9�՛c99���ܠ����ş�d$grvy'o�}fR��-'#7�� ^1��8��?7�ji�%�U]_]˻w���otO*�YLY�����gO��tM �jt	׋�@��
�q��F,��DT���;���ރ&��r}}#��}m�0�h2���KM�~��޼��&D 0H���&��cv���d1�QL �x4�S���{}Mh��vI����)���fhQ�?�$�}��;��'�u�+P�g���pC���A��:���L���+@ۖ���*���]9:ܣJ�I�s�edb(��z��Zq��7�3=��[������	�̓ �;Xx��mO������*����Dy��i���OFT� ���Ãc�/6WE5�8��Č	Y\Xgɤ���K�# X����r>����#y��^�פ��`O��Xӭ�- �|��|D��/�?�׫������zz�n5ܫzM��p��Q��<�����
��X��罼�*s�6�Q��#ɬh[��rU� P�\�d�դq4�L��K�#9W0qH���w�<������'�vmA$����4t�NO�����
Mܙ��J�De>��"o� �C]���Y�- 0C�Q뉂Vv�q����!������?��u�ϰ�ݣ���/�)�c!fwoK^(���O�^<"[��u��z��;��y<����Z>|��q� ���������r����
��z�@���|����P)���uF,uL%����� .��:1��IQ� ���3 �w�?�
��F9��RҸN*5@lE�$6
v����T �I=�̕��c�zJm��
L�qN,g���ǰч�e�s_o9Y[V����S�֒j#H��X�{'v9�<�d9q���p���XED��v/b2�T�.����c�kYTE)�����L]��5��&R��T�8�U�F�����q�ع��U�P��D���CP$��	���Z�`���:���F����,l����^e#��~EU2p�+�;�>�2X"��1Al1�'VF0%u$O��*T�7�����5����3p��|b��3���"$�\P{YNEa�4����
�&70��.�$�ݘx��0;!����U<8��8"�kJ�VJ33���j"�ј�,�|,������ª�̺B����ʥnL�����ŧ�y�/Cb�Ġ�Z��ll�yt�(���[�����\��\�'
�fz��f�)�S������Q�no���Zf�+�|P)O��L�ID�U�qAЊ5���	�	���L�EDzhIz�~d)����ps�͋�$���K��P�*��WcKh��$%o9�(6y�N5:TkZSI	�6����G��3S�,�+�krZ�m�� �s'VT0 �ׄ�����҃�JV�;�;x��*%)+��jD?̀p����uX%i�O5i3Hu����y��-+��6�[��d�A�������@�,%1'�5_���k`1�5���1׋���"�h8�
��N��sMP�M��o�0�n��+�Q��U]7'��P��{V3n8=V��l!���(��ӻgR����e��`�������;H�@�3A���%�1⡂,����]�ҼL껀���-��"�O����TF��Pe 8Ei��+*Ai����<��s��Y1I�2P�&�4u5�:�������+&���M
$�쪉F��M��ۏ���g=\x /A7�l�&Q����SA��@�ݣcP�z(=�`gO^>{.�7w2�̸ؐqi��g�N�p��@�t-�x�,m �!���.����ŽQ�zk�����C�X�0ph�@������G���P~x�L��������3��k�����߿����r��>�����U��ʙ��Bࡢ�1�]��D�&����T��o����˵>������/����NϢ6��M����=?���铺�wƃ{KA�|.�ݺ|�ɯ�~f%�vp����n��7O�/�^�����Lz���=�V5�܌�j���;�m}���{��5@����阀��ͺ&��������,�f��آ�������ءI�>�CM����O�y/Ot}u,$A�b���9�4)��D����d���B7l)㙂���U�^O��k���?�Q;�Vf�TT޼|�@�\c�ON�N�:#�M�J]�o����U��3��*�}��2*K���C� [7,Dh|�"t�j2]Try��g��*`M:�E*Q8DAC�OA6�y�Q�f�a!�M���It�`���ic
��d	���i��Q���7��{WG���^�9�3?��n��˹������Gvz���������T�pw��J��t�*|�c]K�2}�
���~jupx"G�r�� �3h�o�eW�$h��O��J!�r۠R�֬�u4�Mi9���E��=�g���<�Nd��g�q
t�I	59+��~G�J��g������\�XG�e=��w���������3��NGϤ�އ�
�z̍2�����J�~�{��BA�-��Y_���g���d
(O��u$;������ٱl��Cxb͟c	l!�O�L5� �sd�����\���ļ��%�~i��:(�ʦ��Y��=�՛�{(���
��k�ΑV�Ti�8��te"�5��$�y��� @�dy-m�T�*3��5��v%���s����`�d\A���<b�mC�l�1�AᏊ{+D �xi�Рe65F�
�AG�tB�Z��X�/d���k��I�܌�`�ր��+L��q +ƫ��=�{S(�D5&�%��� P��f(�b�2�s��zZ���/����@��?3N)	b�(�ƅiX��Yj��c�CI���gY<�nJ��,�6���K�d}#���2q���C�R=*z�&,��������%�B�����H,i���� �Xُ���45�����9��sT+޸8��5g���b�*�*�Ea��غ`�e7�.�
,��t��	�h@��\iR��Ć��tS�)�`��IF":��&�+�!�4UE�*`h�	E Ό�\Ę�#�L�U��+T2r�-60��@	��X�
�z��M��(,�OL���Č��	ȇ�B	�st�p:@j'Σ�wrg�1�M�Q�ǥLZ���&��YkA�p='�{�Iy��jgx~e�L9-a�qJ3��\��~,�Xs��A��|.l����z=u
߂�4�FhuCN�$���}AQ 3J%�����{Ea���,�x$\l]����������	�Lv�E�4b[�@��(�\K&��^�;����f�O$��IQ��G,j�R�s3/�]�>���Uɢ8�W^L9P����"����@
����_j�,H�(���L� T��x(���������^�~�guv��D�����@ǰ��8�lA)�N�Ry�ݻ�U�1F7���K�Kղ%�� cJ�[��f|H�m^�^W�+���f".����O�!m����F7�ꕞ��ր	q�bt���-J��)5eq���ߵ�%�h	�N��v�����qH�4MY�@l*����U^t� 0��M���rv;��qν8.YI}���������4���㳴����vv���0����I(�ˀ9$鵉^W� ������,5�����a�ϻ����޳[Z^��/	v|��(
�x0�#u����<��՘]��Յ&�C�529zr ��۔o_, �<�k}?�>�*�𦙣C���:��P�7�=>W��Q]{����h���X��bJ�&��\�4aCRA��ق���m&����k���=����!�Z��ޫHn�������Q���`<99�C���p�TL������������ ���4�i�) ҵ������X��ݧ"bjo�m"VcN����`����u��%�ǧ��{��
ܩ���}���+MT?����v2�M�!�<� [k4�?�}����<VG4?���s�`�Dv��4!]3I�},}_z/qq�IK6s��$�0I�[ɕw�6�����x:>��r��b^�Y�/_�٭�s=}rHe?�@ДMp2M9sE�0F��f��n���i�=9:T����`8��lE5R��q���h�8��%�L�Ny�B�t�0�����������2o���9'���'�W ����~O����x�p��M��u���j`��y`*+�5.&�<��O_>J��%5�=:�dH�O�-�p�XG7�������!
�P�KF���3�iw�K;���`�[Ø7����
ߛ}��}��&��8vY�69��L���A���71c:��AA�DzOG�1��9�򄪣E11C�h���Z,��3C��P�[!g���r�CM��|�0�����{u� ���Ls�9���)tm�~O�x����4,�=�����r?x�{���_p�g�5B�v�)�~|�	\\��D;@p�!nr=��{���ʿ�p&�wC%3��Au��@���)y������_�xG��0u�p��>.bφ����/+Y�6l/�`��Z(N8M�k�AD.M<r�S�c�k ��ܺr�ќq-vR�C�Mxe8#wQ;Qa���G���"�t�Օ��Sy�h9]й�v�<�i���0�PC��6����${��Sq��Lb�qHTd�X
R���Ng<K�Ib��R��P>{�䗮�1� �`�֊� �pmH�ᗂ� ��ϊ��m=lN���H�<��d,���N�P�N9��פ��@��\Y�U���FK� m;\l.U�O�Z�t
�2���jT�ݜ��f
]��P��Zw�Ò�2�EA���b�f����4�;�W'@>3�{ܲR����-gi�Y���t��s&�P�A7,�g��1��LqɂS���'(4��D6��%���6�1�:hX�,t H���T�`v��z�n�	=��+�u��b���c�q�u�wBm���ې�Q�L�q8�!�2a�EXgk{� ����d���� r��D�u^�3���(�<�>MM�
��LA��
�w����`3Bk&f��J�:b7�NJ�����!��U��[qI!�L%�7��П�4���٣6 AeE ��w�֐6f�0�/��sy)�&�I�:H܄!���j.MfIK����8#���y��Ƕ�H��g5=p������o��U�P��x�7*ͦz�b�,�0�T���>'I�-R,&d�V��M�v4�$U���8U���e�q���T�誕8ИU$p�6�vjk��ڀ9��@!��8�C{�c����c|~��
R��R./����>�o�����'*vA�ԉb�U��E$f�us�X��O��Z��z�����  �>�J���,�?�ipE0�ne�����)�W� ����_��s>?,F�h�t������9�B6V��La���@t�`G���m_��MƦTm�'6�� ��˯r�I�ln�2��!Ϯ*YͲgL(��%���`
Ք+21��1c6��n1�8�ej���S�~�$�J��Ӯ���H0�mR���ohҹMCW�Bܨ����4JO������ӻs���&��^>~�Bzj�hl�-V�Fe���n[��s��g�H���@`CRT|+�k-��Ge�������Ky���>���q@�U�Q�sx-����RϪŬ��P<:�����o��ړnƺw�CTT���Xśt'
�Fm�U�T=��o����%��+�d��]=��)x.�ލ�sy��g}�c
a��������j��2J_����=����l1��]�\(�*�J+v0���rtT�3�����;6�KRC�}�[4���Z���p8��|�g�l�Lp��o(v���q�^F9&��Y�dN�ԘJ�x2�����b+�
+��	�Ld{���"胀�A o�$66�@(���GXWTQ��淵�w�o^=���J�gT�.�:FH_���%�j��:���|���A:4
�)���޾�։>�)�#c;����]��Fhjpn1�~4������)�$zP�кD�	(��{"��,r�+�H�}�,]�~h����; ��)��{܏��a:X��]�B�����F�ק���^��%D�����Fd<�{�����4�O�>r�,�Lr��s��w��|:����a�=��Jj��e(�"W��#�x���x3+�}��ý�]���f(�X����½p�@|7E����k4��4�:t:���s{)20FlL!��)w?*#{��t���ͭer��v�q�ȺϠ]{>�aÈ�g:6�|f��ll�d=;���U���O���P��`�&$��T�8�N����XI����F[�x��)ܰ0�
 ��
��jb�ȥ��m��p�������%έ�7�Z���Һe���Cƹ&ɏ*!r_�Y���Y���̙��4�~r�/?��'/�Ç!h��pe4'\�r������5M8��mmi@�0	��9c�����5�g�M�� �4#G�a������ݑ�[Yq�����k>;����l���а����Xy�`>i�T7L����s��%���m�%�V��I�����Ti�ֺ.�ԫE5R��;��#0cE�Z�ilp�������A��։jPI-K��
(^�����M�u�1� f��N�b��9��jS!I;�=>���D��y�d��=���Lf��v;kX����z��ݽ���)&~�Uk2&L��@� �tcDT�G�:���C�$UT���؂�@�؆~o::�s��R�3����0+�z����Լ�h5-	
� dЙ0�?�D��K����v��e���b��A������0�NF�J[(��Aǳ�Ȏ�lmt��!9�ý�X|���I��O�d�zC��������1���?Tk��;T^l�e"�G�"����dx��"�`F	�`�IB� ����Ʊ�,�X��j�fPsQ��̡6��҈ ��<�l�R!��Fs�A������v|
���DYI�PGG��t_� (L�		/�/X�(�L�cL`ĸZ�C@�Eb��oo�����|�x.��J��c�bϑ�Ai=� ݍ��.�����s�[ݔjp[��lo�^h7m~tWRB��S�Y���u�]�s�� u���ŗsg���{a��&&
`t��Γʔ� ���(��c&Nb��{���?��>�L��D�H�	�&�n��؃�^bUHS͵!�|��능��T�@ᙀV�PN v��r&�U�8Y��&���$k��5!���z��i�:�3��9˙��} L��U@�L�n�
b+����w|T �����hN*��qN73�/k�U�A�l��s{^4�w�ܾ����x��l��!���
�J*�U��DG�������
<��3�n�q�&�ؿ�irvk:[�#�z�_��&TR�=Ik<�$x��M��?�a^hx�����_FЉ6�+
�����|�L���A���H�*P�Q�U�RZY�������z��lg�ma�iG��N�����{*�N�C ������O���Z���t
B�K����	@���3�;Bp
�)����I���h2���M2=Z�ڦ�4�c��"YM�� �$���V�̵�&��k͙#(2�����v����Y��T�m��9im |8�@�ì���a����,u��G���'(��Y�`�J�����*���O���99�������5?>tײ���n�k����,�^��^��e��f#'���<vf|�����N hx�M'���ۼ9��L�Pl��^>�������=0�@^,�I!��W�7r3�P�a�ߒ�~S�V�k�ȱ>*�5��y��9VPq�V�� +`/L�A��������������9��uɬ3���P����X���/b����x��a�ʔI@���j�樋��%�m�*t���X�]�<a;Yp��,<��
�(Ys�@�N0��U<@7���7����%�����f����	��]z�,�(}?����'@X���1��| P�`@f�˪6߷?�1�b��.6�L�̈ӋԜ7�p*g�rs�����v�p����8b���o�k���3�ׂ�(���X�4�ϱr$&'n�
~��=�� �0��S5j]�IN�fb�C�S$%��=���s���/u��ȳ�1���6%�AU�������k��gg����\\��  ��������:u �n���XeA�p����W\jJ/�����$��N_q ]@��/}��ՠ|Ik故�y����s���ȣ�j�xڝ���qsY׍C��n��{�� 3
c���qp�����|1a{�`����á�k��������%)G :��:�9����V��ʘ��j͍��V�0�$�T��(Yei��Nt�������]l>\*����z@��Y���O������J	&�b�0[h�w2x�a��ς�n�	 *p8`�҂�(��C���s^�|fE�7��V��`�N�2��� �z���7��*Mv� �E���	�����~J���4Q���חrA�\�a�`���s�(Tmk�*����s%��`A�C�
A>?�~ ;�Zo�,+e+.�[��#D�Δcv����XxNH������	NFq����@c݅�Qt~�>v���|��8��(���Ѕ�,�sF����Z���su��W�f��L�!�B�-h������dt@�����`b<��]k�*]*���������*�7�3Az`���*a�����>c����&Aw5��t�~��Ԡ)�
ЉA���z�p+.�T��A��'A�{���h(zO�v�º��U�)��@GEe�5$wc7>]s���G� �I<̑�g��ݣWP]�2Uͺ�Oa}ЅP�S�㊳��[�X2���|�A��L�w�X��u�L����u������3.�2Y� ���g��	� 
���B����^�WM��4�p��f�`̧���5ά�<W�:���LF�Cx���-Ίԓc�q�^�P�Al�ޢ�`[�%���|�}��`pw��7�g�X@�>H>�>��5ku���b�����UgQ �������"Y�G1�+k\�Ӑ���P��DS6SR��h�#lP�Ѫ�0��])��s��G2��ߣЅĲ���w��QY\�?:��)I��`gc���x�/cj�׺���}�Z�z��v�.wO'�'�P�i_�k�?�&�O�zN����8V*(�~��p�9���8W ���6g=����π�%6��n�Zc�1ju����/i���r	����0�sꗦ<�!����&;>��8Gnx���*X;P@5����̊���[]��\��z*�_/)�tp�-����A������xex}�
 !��@���]cc_�|�g殼ze����
��5�X�P}=�ܓ���ԯ��?��=��\�H��/9�ys����"+���k�b���s���wr��V&3PE���Ἢ%&�����s[
���Ŏ5��m�ts�{�`���BN����ua4��H����?{�yćO��_��/���wΨ����f�6��.���i݁��ҹ� �Ŀ��c�9�{^��Nb�+��s��>���_��:�i��*xV��Y� ��MdϺU���v� �i�����ֈ�$6�8���_Ì̓��F��U	p�7	��I�h\m��G�|D*t�xOȪ�����yg�h��W��<\�����qءU�޸�U��O7�7$=�V9��\c�|�U�i/��c+�f%����c
%��� �1�u./��7U+9,�|f6H�B�������Ej�p�)zP��T�hx��׉��0���p�j.��a���k�z��b���RM[rx��j��F���Ɛ�HY�5C���W9���](mA��|�����=:��0�v����}�u뤆!P�� 0�/�!(!y�tzf(�$���Ni�ZT{��f4����7����"�G� k4��ה��=(ʹXm�&��
\��{��A�\���2E����u:�,����X���� ��	���uFG��z�$	�b毐{'��,���\� Y�mH۶��O��%�F�ej���@�9�ܣ��������G�&��drX�; hn*��¾E6���9dA�c�}���n�iҌ�
%�hTFHp����h�͵��w�����CEs:���R�������TTD	��r��\Gf ��A�ܳ�{��n)7M��CfK,���� :�h��$^����fC��ٓ;�zT0�|A��e	�%12��>'L>@{�vxgaV�
���葁!r�JWՊI���L֤��X���U|DL�ss@̀��8 *Qm�V��(��YGkS�[N����k����<q*�'�\?���\�7?�̙lQ����y��F��i��}�L�d2�k�s��s[i4k��4���Ip  ��С��)jK�^�Thй�6	�$�_x�ļ����G�T��ݱ9J=y�8ׅ*�|3�rJx=q�.�uq��h��ঠ�����l/ ��M�a���������뫯
/�1����d�uΙ�<&��}Ib�����n�����|��b��=��9:<�ӣ=zf!N*����_̴����ťQ>�5@��o�9�}�9r��������u������hib������|V��m�(4��/�(�V0mI�F���s�5�Xd	A�r1����{v�����-MD5�,I=�b�U����|��+ʹ[ ��a���0�o�-�.�̑4�5�m��
@��q���<�3�G1�����dIh����8}pC�|�8��@VRBy��8��[�#p�6晏σ�W��tm]��^`��p|�b:z�ӧJ/
#~A.|t�+0�����/s�boC��^w�f�,eH'�WhJ�9�^�k��y�6�Q S��}ҷWT��	��;S�l����i�(҇tB�m ?���w]���ݸU�)������4柸�0����3��@O�|(� k�P�a�jEYyZT��lő�l�p��M�TVΣF��=���s)�\vmL�� w�?�s�ۜ��J�h6k�����׻�)�q�W0?����i[�=��3#�c�}J ��nEf�@0p���B�}F��f9�.�ـ���F���k-r��pTE�+�i�R��(��9ݎ���}��6sl4`�̐ójAK�?�}����P����f��C��Қ lF�jkD�����˃*������nƊ���/Թ�Q`*�㱏"�|��k\�$���4e
63ޡ�z��4rz�3��7@,�����]�	f��0���?=bS��Ҭ�AY��1��am�G�c!���$�dE.����&�[���D�f�<x���RC'*��$2Ie�,�8�t �3��s����m�0Ț-C ���I�I���lߙ���������y囎\�U1SP� �
��Z�Z��_�p$V2�Z�='�]y�����NJX+i�!��v�y��T��x ��,s.�,���_>�t��E�G�֒�����I�w[|#�j�bєe	OGևF��g�q�BY�7J��!�t1ș�{zط��Ψ�G����&�_PEL�	��y�B
�w��es��n7�G�)*a=�[&-�*i��bե�Y�bk+�x	�c���H��n�����?����n��9gf!��˅񈻝:_��6
L8Ȓ0��;l�&]K�O�����=��)��$v�#���zƙ�����z��n�q����g����
�}]��NI1q��)0���h�NB�����-�)!��M�9x�������hb3�0:�k{��у�i��M3��/��2��p�M��`�n_Q��A���]�S�Hl(�홬V������@�	J^x�0�L����zh���#oh�}k��V�?��1)+,��Z���GE7���1(f-@�P�[s��^�'�V�L�=������S���;�]��(�A%wLJ�@0Dc�r��������k���_����'���KJ6���k>���Hn4���V�5���v��>eL�p���yph@���O��̧k5�u�VN��ld�X9���r��k�A`�]9�'�v��M1�{E��`D�f�@3\($��v�8��|O^�x"_�*ؿ��B��)�u��,�M0�Y6�	!RR��KRD��P�آg�vw�LH0�e@���@kz��� f�r~�k�(墓��3fM�����t䕞��{���b`2���n ��BLdL��E H�ˍ�
�~݄Vbɡ�IR��t�9���QBװ�2�4�������S�-�i�/xA�Z�6q��ʵ�EG}��n�*�H�[�ܧh��)��I��z��g���s�|� �7'��z��)�
dIQ���88^��"�`���H�1�����;z��
�ZR��X\	r�Xc���E(�����q.�oq�&���{�^*��_l�+�Y�;�
O���&��E����@�b5��D'ne�{2���o��Pc�`-�����RO������8�_����c��5��	� x(��yފWS�U�%>+`�`t���y^k\�z@�v>[�P������( ҕ��5�ĭ�LۺV����n��p�v[��Eu>D8q�Ik�y(l5�.ϩ��������h\���cW*��|!��ڣp�+tߗ,�,(_^��罯r�����Zש�ԅ������S�{2wL�j(�Ġ�g��a]s:=�t͡�������ɬ���%·�ҏF��̗�Ǉ���1�0��|���m]�4�[���gTs�ӳ������� �H�NS������'��;�c���"��	�����
a� �t��ZG�F��d]����@�9	�'��z��m������g�i��G��>rŐ�G�2+����~�c��A=4�'F?|܏�k4�>j��
��آp�*�J/��0[��	��/t��/�������m6��=q�+�����#����2���6��9�(D��AL�xqLb�r���x����{l�#ky��S�%�����_��M�ҕ�62�.�Q���oUK�3O�M�p�qz#��k���̦�Vq���9#�^>��~|C�����v��b,Q��X�*i
����)�bV5ʲJ�6�$
�GċES9ǝ�1�L/��'�Б��U�$9���F?�M�^(��@^>(���[��-����X��[�޹'��D�ٴcvt2���&�,k�>�Qu�(�*`FO�ɏ�W�ӇMk��9��F�a̅&�S�-��ڑ ���e��h�L��\����7�MD��!eu���sp��=nf̱soM�����7�[��
��X�jhT�y&M�;5��>n����Ȕå^Q���Y^kz�A^ q��P�y��  s-�#��-���9m�YՇ��~k*�,y��P�	w�؎}�Y��em U��$�o�CϠ>��R�zh�� H��T7���wm�]�Ue�ssl�'���eC���(�i��ú�%�X��� �3+���Q���ԓ�����K���N��͝\(88�J�K�m#�Â�D�x|_����TPD������~�HU��1n̓ʙy5�N�.OO��y#���?ɏ?��gOO�\�ἃw?Ⱥ�:q�{{�J����2��Ж�z�T>~:�[�y�'VL���$��|y�y0�t���R'u����vON��ox.H�Y%3�H	_�b��n3�%𛩪�<}z���P>���)a���܏�<�`93BB�l�֪(��[�����=~�n����YG�����v�M��~P���������]��j*��P���<"���������7��`F-�E�BL�B-v�YaĊ{xt 5T���	��L8�Uz��~[S�fцQ�!N�5��ɉ�m&7ibq�cP2���aB5�-	ޓ���Ok���J�]	;?{m(�
�! }�I�t|"���r�e������ڡtT���F���:-�
j���u�8�ą� �J�R�������6���s������Ͻ�9o^q����I�o�xe��J�	��N6yQ�/�� ks�H��^��\
�?������� ."�F� m6a�b���>v�󗕌W7s���nweg�'�[[fUPZ��
�2}�V֥�(���|#X`��BE��"�=o���(�jE7����`�A���^�������p�2ԯ����3�`�l��I��f�ۇ��M=9����&��xbL� �;|�bA�*��`����Sy��EvZ0�gV�2z�Up5v�*6����w�#����W�J�+�� ���,�[�2�(bA���Zۗ�~x� oN� 0n0o���g9;���_���u�{q	q��`f�����BahM��&i��>�Fj � �L |���NNN�5��m�Q�	��[�In���c�<[�n�@�MAk�:�b�/�2 ��U�����`-0�F��p��u��aF�3u�+iދBMe-����GVKF�Y��� 1���uGQ$.\��96r�؅���
�� ���(h:�a�j��:_T��3��Q����0���|igA�u�P��,�yp�3gvѸ������y��Է�?�A�c��E� ��]���o�7h遺z�,4e��L�6�4�!A�F)L���=��AZ�kD�7򇏭�0O:Z|h��H6��&#_���Y���0�uV6?�{w$�R=RBk��۸ %gljz@w���:}�z�L����&<$�9��s�z�Ip�H��  �>*���"y$O�^'P#�)dӒ�u����'
C��{c����	!6ɗ(�:��/á�>-�9�Z���N��[���UW���%����d�Ō��Cl�f3fŊ���+�psU�^g������K\兜]<OdVN1��E�>�k��A�̰uz Wlz-n��(��ґ���C̗<PI�z(t�ޠÕy���(�+x��9�Z�mۼ�Z��\�B�o�֙��zw��ftʸ�,��ȧ��>VPi�����(��:�	�6f�M��^�~H�[���#<4p�"���� s`Hz0���k撍z�f����mp�q�Q����H�fV�R�`�Jv=<"}����sM�TX�=�D~2�������TW��z��l^���%����)� �L�p_$��G�:;r�ua�)T�ؽD�.5z%n��%I)I�ށu"~�)���X�Eԕ''��D��g��kK�����@�a�V"�g��W}R������Y����cE1�=���޶&�/�?��o���gv��4Ƕn<�(^p�"�>��'�O���5����ى����דf;#��F���l���S�R����5I����,%�:<ܗ��)�Ll+s��I�9�� Hf�iE/���-v�С�����IXTS�B�L*{�p0G������P'�h0N�Ks�������m99�����l�IB`���⌋��k���ں��h�O���o���������-~N(��H|C�7:�8�$2oIRW���8Uegc)������l�Y��}~��<�L��vܶÞ7$��8ZU۔GyV�F��Z%;������ �*�L��J0s���|����/�[�ON��ٳc�����-���)j��hA����eeF�H�ҧ����@�G#ڊ�?X� ��ZG��}M��Y��\ι>�y�z�SU� �ҷ��op���z��P���� z�	� ���N��ӧ�7�Wr~����*����sV���(��l�\�tQL)����Վt]M���07�\�g�����ٛch����q���KS=�sT��a�s��k��-hT��=����L��(H��X��םI����������뻧�f�!|�������{��x��1f��C�£~�U���4Т��8�.P��v`��W�^r��{"%��hEp��b�[	t�����������z6Ayp1��� r�^�k
�����v��W[󽚭H�����HF��o�������~Yi�b�zg��n4
+��-x�t:v�w��2�d���Ŕ8����7t�K�]��/4�|��j�G'k��� �б���HL��(��_(Hp*��n'b;b6����Xg,��l����(��UnP�1:�D���Z���KP�s�����E� ,6e�o�Ȭ�ې�¿��:! ¼�u��si��9٘��D�6�����(H�0��x"�>өj������Yn�}����|��|Vm�5��n(�G��-f	8(P������@뱠��"��o[g��+PCݻ^�; �r�j.K���Ɵ5��ܗ$$DQRΣ5�D�iP��a����8~���0D� <�[6���T�@ eͩF�6bF��%+��9S��	Г�#99�Ʒ�j���3LfS���� K��ki�jC�W�Ҹ�n�?ȸ)x ��g!�:q%\;�77?���G�s҄b{�����-�`aI��K��"��<x��J�#	�?��w b�����	7�Q�l���3W~ӱ�&#��̙����:Ws����}#h�s�\	��
,�sVm�,��|{׆I�̪o��ӕ�9����F�	w����Wp�ͬ�9�����٥||�I��m�~�B��9�; i1?~�L5E
Z����VU.co����91���RbO��J#d�{�Xw�\��<q bM��	�7 :�$+tqЀr��d
xAEgU�^��of<��� �:>:�D�H -���nD�uEA���zu�FX7ir�k � Y������{������+=Mޑ�%���P�	&�&w
-�9a���b2��&e	��-?<����36����r�	�����H�k��@If�Z�AU~��.�  �Lf�Q㡺2����ٽ��T��K�S���I�C��9a}��l��O1��*�m*�Ӊ�-��x���㺷���X~��wM��I��{ʫ��I���Wz�>Ѥ�3o� 4��B
��E ���3s�Ǉ��Hy���]���9�/@�P�q�%���[�ǜS̟���u�8E�� 0OQ�'��i�ߠiFF˱���+����=u�e���[fr��l*p~.aNI+�4.�d^&���@���-4��v��6�۳���D�D�7V�i��Gb�&�#�r���������~�N��h��-H�?������O����0�/֌�c�O�ocM��Ln�+�[@{��G�%�VY0C�]2��8j5S����&���Uh���d[w�@se���ͤ���j�k��2��ܺO�dF�⩛~�M^o��ǂf�T> �Z�I��ß��,H�C�ʳ���W�z�o:CUQc��Q^�]-~N�6�o�T�p���@�<����u5�M3Ŀ��|y*�����

P�y����1$��up�,	�@�稲į���fkRq_M���{����ѩ	7��P���2!���@�fp����x>a."��f� �\��"��\�9�0RH���s>hޒ�k̺�,6~޽�,��
�V��v�=7�m�����Ӻ�~v�
0kH�+��
�]��&�/K�Х}��	gN1cDS]�a��
���@���ci�ʠ8^�_�Gp6jnt&Ϟ*��XW	:Bq��'z�(�����(��'2�j��ǁ��}=K�q6�}x����s�4����O��	����c�ܨ�1�%llf�v����/�|+XE�8ـ/$,�MY{�H�@�^���"�Gu`���]�V��nZ�	@6��Y�]AT�,.@,ř��9��R���J.@vx�s
���,Ź��Y��	�Z�֞�G����#h��>,;HQvFE�0#�y����)��7�օ_"O����� P�]Q�W�U���ͧr�iP�i��-7\�Y���,P �@�`�` �J�5Wώ���8b)�"gU�fP��ͧ-z�!iY�:Y���uo���2�Q��B'��B;�#l%���Ԅ\G^�/y�o�L�7�h���5Y\�}Y��#I���:w�%f�@�	:8CpL�sW؋X�7��h��qÐ��b�0	J + vS�q�������FJ� <��rJ9O����ډ`�j�!���恙$�����^ɻ�_���-WT���EU�J�����6�끛;�B%+�M������\V���T��m!�T"ʟU�I�kMWN� :�.$��/��(�}$�A2���+�I���q��2o�@�A�~�_���\�'dS���c�6}��m�ɄPM������k�`�<���4�c�=�<)�[
g�L��������I��ޞ<y���A�	7�ى^�U�FP��v�T%�K$W���>�hT��͍������)���G�PY��q�8 ����k���� 3T�D�~tp�σhg;e�A��gOh�����-�.��A%�^�h3s� 3�?̽���۱\���-C&�6�ݾ���;v�$EY�_t����J3�1����SJ����S�m�l>/�����}���}� �>{��7������*@�ځ���D>~��_��|��He�gϟ�R����%˨A�A��5o�V|F�?����>)3l@����6't����4��Ɣ���)��$��	EI&z4�n�!�Rh%&e ����XM1�]+��[���;G�K����p��@��o*R��VЄzEsH�iK�R��ئ�Z��P��w��|Z�����}�G5v������p+_M5n.�CC�vvt_���? @���O���ҩ�6���HЄ�:u�{����N��A_�۶�j�Q�\1~IP34�� )��9�hՁ�ٌtIT	���']�M��g��)a����Id3EP�T@��	��U5�S���m>��ݕu/�A9���d1^�z����D'�C�]���P�+�������U�C�f~��Jн�0�d<�Z����w�|6�&���4�v�i1YA�q� :/�؈�]�Ğ1��ڶ�����ק���S9<�"؝,׼��&�6t����+����Y8�'��� i��0Ca<���ҳ��gC�=���.����
�[ s�����џo����7�V?#�I�@�QԌv�]�Ͱ�(�`���dD���zI	}|P�1?�?�`?�FT��o���^[��w ,� ެ*2(Z�΃>��ƭEAT� ����gm�B�8�����gЇ��?(�1s��m�;r'6�)n[��i��E� ��S쳙L��N��oYW� 7�*�T`qrБ?�p(�ˑ�yu�bUg̴�$�TYřk�T�*�(b�&���)mKF���pЭ�Y�5��sMj�[4q'�ɢ�ͅ~���hd��	�T�T�|�ǯ�/�h#f����<)��2��>#�!z�<��~��x�{��U�"�A���@���b�ב����@�]�<}�o�p��i�r����<I
+��͌9\�÷����@�{{[Rkf�5 ����j�ݗv��*�`]�l�����z��
����^C�`Ȼ�(CYs5��X�XiPHع�" B^�Ad�*�����6�pS�g~Ԗ�����n�x�%?������~򎴱��TAq��B���l5:d�to�Y��K4)�&���4�ל��睞�=�����-kN ��8�^���ߚ5|�4��d��~9������Ҩn9{9���e��Y�Ydj $A�O�&#�[0�P�F����%�Qi�F�jK{e4x`%�����؊j�ߙb/
�ȋ ���fj�Y��&RQpe /����n���Me���v�ޤun����a���3@��t�} z�^���\��Δ��#��Y:'W��O���k�So�.�����dfa����Ty����X��e�T]Ο��U��Z���d�~�9���q�+�@�&�;��hyBE&Z'9�g��tC��j��.Q|��,F>�4]��h�b���6v�m	�$>[��D�2�Ve��|�ڒ:к(ɎR�v*�
%��	om?�sPQa�>fU]O(	}��Y�����|�D������QanQ���1 ӝ0��P
i�RI�n� �7P$B�d���!�������noL��A���49���(�C���qտ��'7�
$tx���Ϻ10�C"~����/�h��D�9��(�a�Ƃ�~ss/WW�� 5 ��l�|D����Uȼ�l�{6����y<��k��z�JF*�fw ��R�+���5�����'��R j6�ى��+�J�8���+�Lh�g�6�00܊��C�o=$ �
/�/_�l��c������w&����`�����d��0�B��J-(��@<�،���Z��5�~���o�&H�?ؕ/���ݦ)����#�w�i��=D5����m�R��f���ϟ�������ω�L/�$��a,�.�mTPR�����I~���|��Ax0��h������W�V(�V�|~��;?� �*]�"��TC�^�ٽ!�F���x(���y<�T̈́��_M�)f�ń���עG*r0>�|@�.�5AK�w�f�s�@�b�-���4���)���MvH+�d�ɳ����H,��d�����P�Ov4f�4O�X��=xt�+��R;��xB>; ���/��S]˚������mq�|6+X�������'�ǆ����#N*�w���P�=bZ�7��S��NhBÐf���1�u`�����6��NQ�DP�	�d<��H�ҚJ`ww7�	��@�m�L:��KR@U��(̇���N��3wU(36�ܔ�y\�j������"�3�A��"�1�|��n�{J�?�A<qK��Ju�mأ������Iq����CA����\2�!^_�rmG0��%)�%�y;]Pwvh��,�.N�ȭN ���,�Fv}\}��j�ʾ��5u�qc[>|<cWe2�2슲�y��f���(.�\Er����L����}M�	0�Բ�|`��qp@cZ�'(Vx�.Pq�B�@�a��i=)),p�� ����i�؁�A��i2��E\G��ٹ�h��k�f�ks�a�(pm(�M�	P�*FA���5�`�қ�x�S=��f�b���\tD0���R�ɩ&��7��|K5�����ጝ9�C����?��|:�guzr,߿y���sv��tx=#����K�s2k���� ��������,~�^�ᳳ3�"�쿾�`�>J��Ln���v@�`n(��FP�� 	T��]�{�p�)0����J�>qm�T�H���5�ك�H;F�jIkS�#�������>��sIl���{Z�8��hn�^�J϶�͂��K�>��añ��� R��d&/^=���O��f�f�,N?�%���aq=�
5\��:'(��5`���l_����Md��Z�1Ss��˯z�"&���OKݟ�[�٘]d�����g8w\1'�}�"̦q#�n�ٽ&��9�������*g}�p�JPB�i������#��e�2��be9|�^u��8��VlsI�Ox/�}�里������q<�Ԥ�b`ܿTȣ�>飂Ϸ���G�\{�tA�8�������߬��rX6p�M����H	�G����]���󾽁�V�����Ax�8��� I�p�y���M�������XG��c���P�1�2�-(WImU{/7?�EUy��_x�Ea�8@*G�A�"uM��a�y"�v��e�Fk��+&8�	��!�����9ݜ�퀣���׫y������#�PA�����i ��A�hb��cnxH ���5�,K�A �P� ��8C�3Cp���rMdF����,N���c ���V����7��{��]}}���z���{*Μ?�a��%~���R�/b�����r6a�[��q�~��J��wwwD.��/;7����!�%�`�`xw;�����,�P�4���eA���w��LW��뻹k ���� ���̙���yq�����f2Ś��{0�� ��{iL:#�	���P?���a-�Z
�`��{�_

��u�`�@�^�xĠ�^*�YV&�-���~B��4�a�| �����!�Ʈ��������>@:���Ӭ�|�"a�� ��5��(���ْ�����W���:�5	�g�H��y�\>Y��D����A/�m#*ۥ�>?���mw�ב��!�&<�f��u���P�N�����)�Yp/2��NJ�������O�hǑ{��L���ߝ���_�	�}t���1���I�E�����}�M|�6�^K0����?����n�X� Y�5�::D�$z��iltS
D8���맜�",��AC�u)L`�y�*%�g4Z곺���8a.��H��
 ~��e@�*q�����>{v"/_>�
]q�{�`׽֨���Uu���h���w��R��i�{��j3b�Ui���3p�C2�#��x�v5;�sSOdӳ���%A&�0s���]�$Hsd�?& ��cw41��Ȼ�[�[ήZ�o��G�G�#Hɿ|�	$m0�F�2e'��",Okv{��� �vaM�(OO�#O�����o߲�����h��=�5��-�z�+��t-����@l���f9�4.�3���&_�-R�r�N�Hc됾����� �Ϛ�C:xd3t>P�]�mM��ܓ�A0JtJv	�O�%+������F����b2���3�������Xt
�c���G����l�����g�I�,h$YqT�4��N����ݓ�p"����[63=�npZ�Y�`�j���}�0R��BUfd������*�XßON��o�ۧ��L3R̤�0)��s�ԅe�XM)��Iݬ��N�I��rV�󛠵�ϰq>F�D�� |Ji����E�c�ݰ�$���ƆGY�C���ƺq-<z|���o�<���zĬ&f�11�����`���!�>M�YH�c.���<�Tamx_qO%p0`G�t�ϟO�I=���F�Wv��xFB��l�}Ft�a�=��:�7r�p���sJEn�C�'���R�I=�'.�5pu��E�R���zq��g�L(�'�+&�3��qnF�� lQ@�l���h���a��U�|k��3}>7�v�^�[�.x�b3d��X:5M�:�:�?�y�ӆ�v���J��ؿ6{��Q|��YNG��;�g�)Y#����et�r~2�bs�ƽ���v�X@Ц!��55��'�B�|�y*�1~��Q���� �����P�&w��߳�b?1/��#XP�\\��؋KA�u���Nj��А��g�g�1��XXoQ��i5ZRЀ<8�H�WB�q��c�2���}�0��>�P5��<��yL[t�u|� ��b���\��^�o%*��\E�����J�J����.�K��΁P?����0�Pd����;��t������?�@oz������M�x	~;K��,����,[���A�CV�
��Qy�MK��:�t�4ar��M0�/,��)�\��ă
8����������P�&CT��fAþ6�-]FB���"H�>��uC���\��Ԝ����51�;/����T���3-�br�1Y������Y��9�J�P�8��S��':�I��~��C_lZب��D�k=?�9(��@���,��\>h��\�����U�fĳY�K�Ko��5U���A��Κ�~�ȝ�c�����M%�Ҍ^98Hr�  O��a��eY�����U�5��?�RE�e'
�jF��>A �8^]!�_p������0��W�Z�]	ս���"޻��Ʀ3��6\r=����I�����>���A�ڋ����YL&�w
&(�(��	~>��M<f1���,�������jG�8�����~�îs��C>�$��Ku�}F k�u8a�f;�a�1N$����p��~R\e:e���d�������-U�(B��~@z��y.vR�݃c��'� ńh|@JEAq�9�9������v��n��{>@�Y=%� Y�7�<(Au�x�YUA>�W��������#�w?��m�np���I|�{��0�nZ��b�
�GA��sYd��^�5{j�����˿����/��Q����g��W7�`#�������v���74��=���ȵ
�it�H��>O�~����~��{HeAP�I��h��7A6���u��ݨ�H��=�wo����p�í�5��ݡR�����f�س��$��+��^�k���,��'�E0���x2P܇�^�X�׵~7������d`��Q�ν�R�de@<h�f%��A~ wl�$%<ce�<��쏭�m�ۆ��ݘ|Y��*]ƓԚ�zH�1�9g����˸����W���ή
/9��
��>|��~��{��||�xȄ����s�N<�2�����9�c��S5"7 Y�c�a:>9#hd��A�服�ac̓���>9��������w����)|#��@r��}��b�o|]t�K�v3��)Z��<��tJ��c5\��Sm�;$ڠ��)��,�Y����hW��.)&�����ͦml�L);���E��ɮ�]ю �A���9����9">cOMc\:���#Q.�nÇ1V��:":Q����IP܀��xm��=xHn�8ҷq�y���2�W��g���l0�U6P>)f2���B^��o <P��,A�JI%�3�[/h�{	j�Ѝ��k����fd�&U���\�Z����:�`w\�\�Ȱ������C��;�v��pYjV�H3��5��=_�"��a����m�<O͜���X�)xmg�(0\QmtH�\|�W/�P\��'K2T0G޿��=���a|�螽z��^�z��:~���=�x���T]�La]��6�����������_ �Ψ��*AL�܁��Lʔ���8@ـ�_CD����/�����*+K̃֒X�P:��_+�+����)�1�Ub�I��(~�{\�����;X�Z�||�^��V��dĄ���K��gpd�B��]�y�Z }�q?��VΔ7I|E��X��L�׺pR�q$@�=/U&\ޛ���fYY�H��Dw��_�D��űE?G��r�Afg���+�?$!���d\8�4 Kp��������V� ip�K;.2�7L��$4)6%���:�X(��xY�՚�2�
�,&��Wq�]q��3�9U�Pa@�M�U8�t�⍃���;U/��u�ZbޢM�==X����!�� �jV�!䱈����:^╒��TݥT1 Ii��|Br��%����bU�sU�Nk�ز��h�����.���`�{>w���'����Սr#$���0__�1���WsTA����&�"���<Pĉ���9�peP
 Mڥ������b�x:=�I�?6k��� �}��$B�
p�N��\�������ZL�����Ν�6��6��b(q��XO����>X���ݽ�M%[u�������� �g#Xz|>�Q�g�)RI�@�5�������l��E^2�H�`�:�%�����$�������#�pp���ò�>Qhf�߯m`�X�@ᬎ_�3���v7����x�A�b�>`W�D�\s�"��1�`���d-���[U�r��%�?�����߻��a�RFC�C<AWA*�KZ���M�丷�=V����Q����5G���� �8�ءPsY�u�ơ��ᣮ�?����!̸�<�Ҧ�:����Ͽ���Y\�O����Q����87��Bt�߂Zk�'�UZ��r?]���/ya�����iz>`uq��M>~:���۾�͙�t�2Z�o�>&`+>ۧ�?qƏŕ���V��ȯ�~m�E�9�bZ�Rj\�X�X�d� ���Z+u#f�,���}m���?�O?�@?)h�0���с��ۧ��çxo�.1��W������~0~p�^�P")b���kz�K�siL����D�pS�ʹC����&�<Y��!h�H�!�����[&.(�d4H�7]�93���uM�֜4v}q��v���>��A!묞��qc��1�ݸwvwY �Y���I���ߵ�[|�D��o��c]�>x��
�0|�A�?_ ,P�>�P�7�9��}ru���wR7��gTڠ�
�o$�Xp�`�?��`�l�ݘX�\]���-)��Hll�sbm}�@���]����x͇�L�z��h@;�:�Ypp_,�U:��}�ֿ!-#�V�5�e9�o��U��J�@k����;��>����u�Ӈq_܋�%���uY�d��z�h��f���2�n�0�u/��u��<��;���xaI%����i�[�����5�X_E����ݸ����Unqn4T 4x��om�w�����xW��ﳛ�xn��.,4b̸����Yu(��`��/ ��<!��e�S7Y*���f��
~���X7�!��p��P�CNFq�������<�+��~�;�5j�����.�Z���d��s���q�O�i��Ï���Ƅs�dSD ��+�8�\��#��?xp�<�bW��S���
Vr����1���ڧ���G���={�|
��R}��1�2 ���Mtm=�q�~�fx�Yh+�6ޫ��Ճ�%���k7K���]D����>���OX�E~
=���T3Y�Ӈ;��O�9��ai���*�ʰ��3N�)��Z�,ԍ¨�,��4: �Җ�<��sR���p6�\E��#A��b]���������|��BȒ� �Ӕ�=c.�֫湐�%�~� ׌�?��k$�t�,�tMo,��#�k��u�͊ ��>���n�wI,�`)OR�"�֕���-�y������:��s0aZ�SRy�M�p��py����^��X���%���T�L��8��t;��C�7yz8��W�		7(<H��R�M�8��ߜ������*TIz�|@���]Ġwf���X��\O��@�� �z��5)�����qAې���F7�A�V�@�Ԫ�ϙH:�s�p�� @iYT�/ д&.,@��o�!�?Pz��cq�B�gհ�+����$��җ(pc�j�
W�m�z�0c���k��~8�p�11�F^8��q���\�64��= qʾ�k_� |A�_*���/	ԢRu������Ft�:����?lA�pae�n�x �6�k�D�K��)���,���P���$Ű6s^1$�q�5q=��+G�WQ����H!�:��Đ�ZM|����5��C?o����/ȕ_�i�2��ᮮ'�r�ZZ�P�LDh:QL�NC�x�M�g�e#ѓX���_|"���<p����qRQ #��C�x&Rr�D��R���7��$o�e}U��j(b��
Y5t�|�	Ҥ�'TP.l�xK1Mn��WC�����2H�����&�0��}-�t�a$�rP�WPfH͛.d���	(����OCң�c
Ѐ6��A�y/u�ZK^>I��2�cr	5�uU��7���/��?�����o������5վ��pM��c"���G���Ec� �[�Ae��#hI�����ڱ?|�=���kk�3���MX5�dcV�h@W��,�/�ڿ�۟���WvrrƊ!|����R.�ğ~��_��ĥ�KőFː'�������3&A#���g'?_�ˆ���d�H�v��δLϰ[v-Qe���OL> 4�c���`��^��ADb}��?,� V��_��?}<f7�(��La�JP���O��CR��Ɵ݁�\�T��o�2��w���?���O$ʠ�c-=��}�ƣ��aot�8�g�C�sl����}���9�/�w_���%����J3	�s��=v��uˊkHk�U������2"�D���W��'�Ӑ�F��X�����N �?���䣓��	�2׉r���c?|�=E��~���^��<��M��x]�\�������f�3����
vl�� ��l��ՉJ�������4�f�dm�Hs%Ng^a�$f�)��7�W/�R��s�y,��6��Ɏ&͸��Pˤ�&�<����G�GR��P*�R^;�יSg1��-�Y�|�y���	�i7�y��I��cAm7��{�{��J�\Ÿ8��8���AL�{��/�����A��C�w� hA���b��ͭ��8�a%q{�ၽ~��
��"��1�D�����y����*Ʒ���X�d�i��ی�x/ juڴ�������O�����~�`�)՞ѱ* W������ښE�*�-�4������\m�~R9�G1�H�k3�/���g���{�����u�������}8d��q��Y�´���-��E��rgo#^�7���*~t}�c��c�1㸆QQ q���޻��={e>�\G����'��zj���zE�������8����؜r�
��%x7KYr��װvO?�I��)�z�gH9�  1�W��2��!G/�Q������q �R���5��k���CK�d;�o�%���L�J��{�S#}~�v
`F��=����ba��B�1�f�+%���O�CK�͙,���a�Y�:+;�AֵKYw�欆�J�t5cV��|�
7+tN��)҇����t�b�1�'�ai���zd�SKC�T�pwiV~s�[9��۔�!�E�F�'\�Жr�ν]:wЇD�y��e�aG
��W��r|8�*�"�S�f�����#xM��ll)IF�@R����N� ���H��CV�k(���"k ����/��P"�^����F�P�e����ƍɃ��:a�@Hʢ˸Hұ."��O��d���0�}R���3t/@hӎH����$r�cT�u͝g޺Z%�T�5/5r�97����`vIz-�4�=�(�� ��y]�:�	�� o?M��š��z0����f'}ȫ�P�x�|b$+;w.r���H�I������c�~���s߸�Q�Ƌ��*�PhR�ڌ�95���K}&xBnH�d!������fo�<m$jgbе3�K���q��y�j����:S�`C~�M�Ҋ����S`�����qSSz?��?	L��/u6�gsP��uO^e�]d�N_�3߾H?5� �S �U*�T<���3�+��z{� ��{3��[̜�$�*�pH?�]p�#9�����7�`}�u�gT<[�l�e�:l�o7'��������3M�q��F�5m�������1�����xh����N��vo'&�%0�^��hd�6ك��T���|�2%���'�s���J�߸1v����&�����y�g5��lз���?�#b����_Q$`'���\�[��r(�0���#�6����g���������b���]�z��g��ύ�f K����}�c�d�[�e����_�ί����궋��T{�г�P{)WS��ͮgvt|m���#Ȝ��ƙ/�m~���3�94��ܝ�;��|�s�i+Z�d��y���ћ֭���fs�l��Acώ�o���_��Z���0�'8�_,��K�		��_���@T���,ݧ�k��<S����������fD��Ø��̵Q��=��L ��Ҫ A��=������@�B%�����2&�����������6�۬$E�����U�����<�B
+g&�1����g��^�^f5&���P	��=����c�ƽ�bŝ��x��>��f�	�,�\/ ��ba�a��*���1j�Es��鞠��Όs��wA���+>�Vv��N"h����ގ�m�D㽡�6�"���#�1��}?�k�  @�v����K�x�n͍- oR[#��E����"^�x$yy�<!�_^�۫�o��G�QSg%��Zŭ̔ZV(B9�C̩�݅0�ݻ� ��#�:�0K�u� �[t�~�����=�\�����i���ɥ.���?fQt�y����YQ�==��f������=��Aį�+m⺌����u}f�x���܆��-���+�i�CX��K�G� ���=��v��(�����1ć�
��^��?��̞=�����?���Y�)����S�W���UDY#���F������?��a\C7���D��Tn)*$a�:4}>��a���:Hd�/J��S��[�2[o\P�k��F��t�Z��H���@�Ҹ[~B>9�\/��5���l��	޺�TS/������1�C��[}�g�yt����|\�Z���t-){\v����(�|��%�p����:'{&��2��ݭ��J(R�G�^�g�~pP3�9�����rz��g,����s�e�$��+�r�^�)��� 2�I�c)0S�;��bY���Eix �x�el��^�Z|����E�����EbMz�P�f��4!�äq�t�����]1�g��X������+�XJ(��H]�+��r�{�+�rKz �T��i:up���y���H� �$<��2����ɬW��$`��;M_� `s����0�ɣ�u�7�f2M<K����y)����0f�W��KVn,x��Aѿ.��I��ݍId�+𽼕���e2N�?�2�t�8t�k.c�HU��_��ߧ�PI�Kx4м2�3��R�%8�,�0�WIh���#<0$ť��AN
���'<�6A�k�dѸ:WE	��<� l���ܦՍ�l�w��܃���p��*n��䮭�k� �f�
�������V�`N��}m!󘐫�lj�\�p��\{}6�?zH�k(qJ	T�D.>���;��8_h&*$x`�j�d��G~�Uּ��@5Qm���+{��4��#�|��m{qA�=�1��Y�������ۯ��������|�B,8� ��ф@@��~+�G���11x�`��:�{�§�"{d�Bg���vS+z z��Q���T�x���`�_ǃ���]5�9n������?�?��O1>�K-y�e����GB�ͽѦm��jA(:}>9��	͡��\*�F��@c�8jH���
��������l���-�����q� ʀ黭mE����7,?����a��?�rǸ��&׷����g�xpfwbr;ޘ�3��	�B
���,��=�Ǻlۥ����
�x^u�R�f�b�	?��xߧ�۳w��������׸�^Z�A��k�ls�{�-aĒi��S�1i/ƴ��{���	'fQ���z>=�����yL�n��yH%�'���$�����KL��C,��r��p3&��	�a}B��L��4 �!��+`�a+4��BL�z=�R�;���������г	�+A/�,YYG�+�<����:y���>xo[�qo�Y~Կ�|���B�8�@��?���fӘ�`�����>|:��o�88 }J�9����Ѐ�|y~bWg�����#�m�R8hX\�-��zi�I%]��OW�nA�c}��Ɉ���h����#  ��,���FN��o������q�N�@L*m� ����uM�!(���B�����>	ZN�8����)���Fcs[2$(��5_$�R�v�bI�t�R��������Ϝ�=�?����Tk�M]�AHt!����v��������м^�"XA>��3x�7ы�еn3>��Mg�/���O�K��Ϟ��l�U��-��q��g������\���L�Ǹ~�?ͽ{v3�.AB��V2���l*8/��?�T��<���u�d�H�V�<�$$��T��4�ؿT���<_%@èQ&�h�>m��>H*�j�B`����и3��՞;�x���yD����\g��wr�����f�{@���|�\9u�
�/����,�G�P�-�9uc�E>IeF[��Y�S�l�N��4@�I�y	���	��֕CHWD���/͔7SlV��]��8L�t0~��O2��}��W��c�~���S�!�RF]�O�P����>��u��JUsM�*�l�I�+���:�ζ��J�<J����I�;�4�K�Gϭ��O��NT=�����E �-��ҥ��V������|P�|�7`�	%���g<������4���'���Q-s�͙D�0� T1S;Z�5��J ����e5�h]��1�b)�WY���o���Ql��҉�ڸ�V^d>Lٲ����۴�٩i���풯\��Wb ���C��)�=��yA"h���^�h�:��~S���Ќ����/���zоJ�:˗vM�!UY�/�%yV���_s6�3���%���5�$�����^ysݹ���*�0�{L`����*��&�_����h���S3�(Ȃ�IS2�B�yq��g� �:� @ϛF�ܡY�'��_O9{���zA�����2�hf����#%���P�܈�Θ��Z{���&��v��o��O�>^�6Ι������S���wd���F��Y+9l�!e|ȨX�K��Q�����2�"[���jՐ�W���	!lGj7� X�A�	P���l�_���#����U�A9�}e�&���ʉ�Q��bʢN*��{�bD�p��4ǝ;ۜ?}.�.ؙwe�i�JF��q�Ac�b
{���칅ae'����=�ކ����3����fAe���?�8���5�&HY� ~ `����������mX�w&�����J�T!em!7�ZɅ��� ����\��b�b����#zՅnA�6�E�c2ws5�p$���S{����A��R,�~������(_K%���KJ�:�x�q�b�~?>����{&�x� 7�{��+;:�ho?ܳ���叾z@�#(i�̑i����x\p���Е+%���O$��� KTjՁ&�<�Rq����iD��b���i��os/�dYZ^�gg��A����!��� &ֿŽ9FR��X?aB-��^�K/XɃtcWu�w�.8����8_����Y$|0g��R݋O̧�v}������U��i��Ex�mD���Kx�܏�4߳d�7��(����Y����RꊝP��TuK���������Z̨^rrA�;�����n����^�'衐�6s�cs��ei�;\g��q�ͤ�?	�2������b��}���b��딳\���	��%�񖥏�rl��'�mv'��<�����)~��k��I`��{������b�c�jc�G���S����ٝ�mmj�q<*�T�@sfxVeR�Ej�84Ōx����/^}��/���wvx|I���:vKq-�`E�{ppD*���eܯ��`0�k��������8-��a��Vϲ%@��]¼������+̷Uԕe.�I>����������Z��_4k�Ar@���ݐ�⠳/K����	�gP#��[��m;}qJq"Y�t�k���1��wϼ1��;�<�邼a��Ŗ+xPY����	��P.�K��Rg$+�u$�����������낿�PI�>U�)��,�~�
N eٕX�U���{��q�A��#���.'Nh�Y�ȁ��c���l̅�bG��D6Tw��U���G��*�vP�-��]JY�O��X����|�� Nj{Y׭$�ލ���MJn����Z�e��j�2�d��;j�>��.���yݔq��4�3G @p�JҰhL�%�6�W4�ݔ�m�ݜ�^NGmP%���o��\?6(�0��Ҡ�ko�W�4�L7��b	y�%���L�J)\f�<6��nZ@� �9&p�����>qБ\�F�yE���'��eG�i8����Q�Xڌ�K��m�5�� 珥 ƽ�b�$An����
�K��o:�|�3X�vޑ��B��5o%c.��PP�Z�&��/C�h/L>��L�]���r�.F���;mH� ��A��[�C�زN��h�s$K�UI����?���쒒��ڣ���d��,$�G@�d^�-�n�QE�vJ.:\��� ��W(���������m���_ۓ���!��u��kf����$����̾��o��yC)��df;&�����#z� Y�:b�$�io(@��77ش	�ڱ���
4-:�Ò�5�}�ĥjE-ż:hb������>��o>QE����Ŷ�h�r��y6t��A��<(�́:@����Lt�*;����.���*T�CG&�1i��n�Ca�L,��2I��a\�.����ή���������'��;���#��Q����S;���b"���0��i��qa1J�=��p��i���F���J�ސG��(��B�7S�Q�ޑq�̮��@�N�{ɵ������qݼ���J��xN�1����S{�8�ӝm���5lo�u7V'�r�|*�'ye���C��" ���!W�/P�0[xy5ejd��C��������&&y�T8��om￾F?�͘���ΈE���Z �	(��`�p��Y*���(�(nI�B4�l	�`uN�5WE0
�=���I�?�y�㉜B�W��b��d\m�X�"��xϽ:���b��`t,,���3��p�Y̐3~b6���������Wo�k���o?��ѩ<�0�J���ϵ�A����P
A�E�ƫ�����6��# ڎ�!����!�0%t ��y<_�́�?L������b�{HH�����ٍ�(����"��=��au%��ܡ�6I�0?�Z��r�y�tI��At��G`Ϲ;;{̭�={��s��ՙ�t� ���>��|']��?��?;�d�s�����ʉ,Jb\��ǫ$�"�{�~=��/c\{�����{�=�QP����6�����.�Ұ��A'������;���y��������7�<�G����9����[��0��*���U��
����o	�@��|�(���Lj�U�Y���?���sy~��sJ��@J�c 99����+!�͂�ԭi��V1#��)?M,�����R��:�0e��Z��<�[�zg�Л#���=Գfzj�
u�[�0aR:/�&O�́Sk�뱑�4Z����h��Bs���O��B�*�s[6��P.OI
 @�+�n���T�j�פ�$������ÂsTv�������߶JZɁu��1�èi%�I51nH�`uV��������A������t�*��  ��IDATi�MtZKU�$ހ��.�q��V�*�܆�!�	 �,n%s�4����ٓ����������vq3��s�x #�v5��f˳�J!�g��m-�b�N]
�c��}���H��S'P�Hv*�����+��jC���Ց����^���y�XA��@x�p������h:�	H��l���3)���e�ܜ���"f��#殖�c�o�$�ϵ����A!�9��2W�jV��wh��q�11��7�(�94�uH�u�P�����&:j������Pq@���ITT1㔧g��u�L�6>|�	�r��2̣�D��
�B��h՛T�$9_��g*b��_�d�����|�{9�2g|��RW�!��e�ZJ�S�Ȩf	#���sAɰuj�����Z��b��J1Qj�0��0��;���,����ЉZ��/Ak��xPm%���J?���zz`_L���ۄNݟN��=ZƁ��d<�=�������5�ݘ���zf���7vr���̦�Y�? ���v�ark�T��{F���>����ϛ�t�3Ҏ��������͜b�{�نY|V��#��Ԛ�TgVJ��߸� �����3}�bۃ�����[{��q|��:������$9��mms,���L�q�!Ї��ٳg�=�O�H�:�?C	V�̮����o�����O�>���"2���q����YLLo-K��
������o����wL��Ppp>��&�PP������(G�@�;&BSP<-�A�����N���Ǐ19��~����n�Ҏ0_�ۋ�� r�3�s�Z�yb`�)�S\�7 F�s�I������v��#�ݳ����$zfJ0�614�~8�^;H���6u�Z��׿�b��d �e%���Xɿ���˳}ۏ�������ݵ?�����)� *A�p1��n9�9�f���(>��{q�oa�͂o�{L��Cݒ"B0������goƅ��x�������}��+����?����P(B��rܰA�`���@����]�6�]�@Ơ�(kkѩ9�	��ɍ��d&xu�ݬ���i�j��)��)'�/�x1���h�y�\M���p��w�a�R�ܰ ��b-^td!.���NSyΰ���l6� N�cr���ƯOP��$��u�gRP���b�6�S1u�s��v6�<�d�6�Mƾ�����{���~[tɘ���<�o/"�x�VPN��?�ê>'��P2;o��4;��ev]�IiG��fNUexўw������P�@k�&p�AK�]��w�X����
���^zJkγ��0��1�8�Ƙ1��������p?�ɺ�l{k�6��Ha��p|�{��i7l<)�ON�"�<��ޝ���G�.�������u��C�	^c ey�e������9(������(���x�g����.��X�6�w��츎�~b���)j����4�9���K����^ޕy|�5�M�7���*�5��{�|8���_yC������f�ˣ���#"�Qsު	���4/(�C5o����AeRZ�̘Ӥ|���a�V�5ϳF�x�\�l6
=�
�`�$�Z�4�ǁ���}8U+�C�����оo='�@�;����z��ڕ_�l��9���/�y�3�D��WF����Y��8l�h�hĐsԩ�Ǯ�\�/B�'%��Dk]�&�@�m��(�Cr��&���uА�s�ִ:�l����x�e2�[U;T���K�֬��~�#u(�.�s�%�mjK�ƸS��/����Vr�lT��4�o�6�j|��$���~�_O�~H�v`��A�L��[G�� ]�d�&�O��)qB����^v_�R�S?; "_��Q�O��λSX���<(ܝVA�����è�R@���+.���-���ϛ%����98m�@����`N�bѷ���$!��`�u`�k��N����������i<qW�s�+�}5A$S��+9�5��b��W��g�?�[��,��\ M�?��=l=h-�P��F�L��`i�}�s���:��D!��M�[^xU���f��2T�W�Сh��)�J򂃔�N`R*�����vW��D�ܛ,���J��zj^��T]RE�t�v�Q6�l#HC� :�u<�yc}2�wK�g�F�n鉓�Y��p+]-���<�a�@�R��4+X�c��b@�1# ��h.�����D_%��_���%Q������ǯ�a��9��IaOW���?�Y�T�a&�u�
�۔X����.��.d���G�<&S���`��#�dj>��Ól}{-&�1��ߨ�!9�������z��^�|c� ���.fP� I08P�p�}�I�������G����r�7���=( F�W������u��ȳ'D��U���y�*,�S��I���F�"�|vv�p���}ppL��[ʒ�^�2���q�&�"-a����Dv���(���7!egg{���[���yU� Sqq�����م�7������E fY�܂{D�LTn�"�Č��g��L�=ܻ��D\����.�g=��	�,��|Z� ����=���ĄLk�h����x�Itj%��:�xX����G��:�����><|,�>����D�y#�)Ae\�q:���:@4��T������u��R5�˹�t�֗�MV(�=��_��G����~V;"�a�c���?� @a$�f]y��|~h$�o0H"�������;��?9��w��'�'�hj�[��3V�}�B/|������׿aG6p&����ON���8���5�F�� ؟�D�����{K>B2�-�lNoU�n]��jv�!���������S����rp�,�xI��K�p̀E���҇���7��A<�l:S��񈿏�pxp�]�}[������m�.��|��/�=8b�3Uw�l���縲{��.bL��<����m�sn��߰`�2"��0'����"��RF�U~q�g��A������v{����v��A��/��y��ǂ�,J����ݮg�Z��8k�d��h�=�pV'_C(r������n���)��� ���$�%�M���\�#[��bC�ob�g���S����U�a/8����x
�`���U�}���c.�+�xn�ͺ�Uß�kׅ������˔���>ϟ��roj<_�RH8h(�T�0xx�u�b�����Rn ��%��\h����u�����y+��o�ߋ/"I�����(ѩV���)�칙��i>F	���7�b_��3�t����N=ol�'Hs�a��#AD�Vq:ӂ���yVr��~蕅�[]y�^��Ww��#xK��C~�@�m*�ɋ� ����}��o��x(=��b%e��Pm���0���t�	!)�B��NzX��ʝ��(V(��A>X L�z��)cFE�AY�9��T�Ҭ��8ϛ:��˖<`��p0ס&��U�\r߻X�א�Ƶ��|�%���Kp:�`��,�|$w�`0& �5@?&lL$j�����ܙ|� �|���M�ZA5����B�vt�o�7�7����|a�<{��"g��Z��cR]-\$F�iK �[���잌��2�0_�����K<ܰ� ���1�=(�
��C��uڗf!��Oz#�Z�{H��m0�TT��]0&�3�����Yu(��巹9��)Y'z�%��U��B�����$H,��m�+c��TG�/B�.�e8jRG*u����p�U�֊����V�e�H,#W,�A�D+(�~�0���3_訠������:+�=����TC�Q�.P
��ö"pufƘ�p@��`�{U����*��/q���{@L& �J{���9������rk�"���F�0t��fbֶ�m;&�P�C�1"��cP�Y�nf�
�J�ut&�7Ό�{���/�2�~�&&Y���`\:�,`~"{`��*�I
� ,aݰ����:�,�Ob�t�ϴ�L��ԤzT��M�J?�I��W7{��0��+*�!����)b� ̲lФ{��TP���I�:����Zy�M��0��crжP@�<˂�=�{�������]f��*���1����5�[Hո� W5EY	P�)&����wg��UP7�1�I����͜�����Ɲm��.\��g�suwhl�)c�$>	����:&�gT<CU��ra/_p�����[�nF�(��\�N�� ҚS�L�$fIb�$�4��aW�{����Z�XJ�j%�Iqa��������`��M$�d�-"0����Ut�P�_PI\��ʁfG�tg�W�
^�Dvsˢ�Ts�3��i.�FG��PE�q�[*6>�����4# ����v|<����&�<S�C|(���I(�h"zkaIX��s�t���
L��}�q+��U`Z�y�э�J	hHO��c0[pT3�KӸ��yac|!�N�� ��6�[?9��o]Ӣ�����`D��x�=ƫ��3����ZcA��1�m��f�7d�\ö��l3�?��!��yY����,�sGn�r�;3Ϧ�� �2\]�F�uaǇg���kۊ��d(�rЭO��A|׊[�!�N��S���R�iP/��0�1�dY��!��&>�ۛ�< ǐΏg p�q�T�(D��x0����Ĭ+���I�c�[<]HN��MCn1��T�]���r`m]d��+��ȭ���m�U̅�̋�!V�D$�4��Y%-�s���;N��sL�l�瑓�H�L����OW�	dI�^�d�4��l�%~���)K�\�t�e�I��;G��-f+/޻��j�����*vTj��H1���$��J\��ѯ5m�AR�K_i&&i+�Y�~�)��@76x��.O�9m�yuLIR^�4�=
_-�)T�Ơ&��Q�|x�=��g[5�`� ��>�1��Ds�hVu��*�����A�6e�^���a�+��83�� )�½��1ZJ�خ�uA��Zp{8���z���]M_��Bb��<��0`1�ښ%�mK�$�t$ȾA@��]8h+DcC�j������H�N�90k�n�_���'�5���͍��W3���J&� ��{���c��C��~�.v�NV�Jd��J7�{G`}�ϲ1Ywo��?����[P&5K���X 3q]���oܳ ϫDiD�ǁ=�@�h$je3W7�l���N��ݴ���'1x�rވM�u<��l��#A��G�?����#����X�JE ��@���hKv�+H��bߐB\4�qd��Pb�N�IT����s�5g�D���-�*%+�/��ˠ�e��!�*ڭ�aв�eE��RCF��*��l�º�����z�;�k���ٹ�a��%ʡi�/�P
�eHv;E�f�h�`*P�ň�5�(n_'�/�s��6�/���L�A�t��)�G�v�������&�'��"�mL���0O�w6,�O�O}��!L�T�C��h�9����g9�P6~KCΝK�j116bKj��!�OD2P�@�������KŊ����;:f��wV�/�v����5��`Q3�-}\j&.��.s�L�D5=$/=��p��"Ƃs���[}Ř�bM��a�10�t^�J�Q�\Q$#��S�Ms�T\ţǇ�	%�3��>4'1��`QP4Śk��Y+��sHؤ�r�����D��!���d���$���s/�02��S�J$��T���|�Nܘ6���ɼ0!	�@�r���t�7hO]����KyI�Ǹ�����w	�850����--��Z/%�:0�-��Z/�]ԞX.:&��z��r��� ���5���iZ��+��gB��r�];셐��DO�B�����%�h����Q����B?�+Ү����;ϙ1�@�U>�O;�Ҧ�:���|�B5�Q��к��.r/f�ݑ7S�{�z��/�1�
��"P�0�:�.s������16�_G�zL 4���ފk�\� b��nn+���3@��#6p4d}��7�qEne�CK�P����&Q�����S�H@�2~�Tk�ڿ�����)�7cnpgs+����D1	J��A��{By���@�a/W�-8��=d�����y.�#P�8�;n�<Eau�爳�L��X���K0F��n�� �cTlU�}8��M>Ko}##�d��]�M�ֻERٲ���T\���=8���{I$-a��^����%Y�O1�����^T�<[��w%�Ϣ��>�%���7d���4�=!��U�7��xHR��S�CZ_�"��?�dA�H��
V�<��.����hW0!�%%ok�����C�k�Wn^���%�[u��k����+�����d����\T%�噼�����j��0����Ab�Z5��GL����"�ҿg<4��C���V?���Õ�m1-\��cYz��jd��� D;�����Yd��9��0p#U��*�U�5I��y���X��=��O��5S�@�t����N&�Cv�d�I1��l�&�\��K��Il�>����g�A���%�I����N���_%��@��<x��9Ej�oP{��k�wR�]3c���'몚��5SQ�2QغL���ke�߄�#7��4�l3���jV�8���S��q�Q����C_X��C"�'��QX�A���,����K�ܼe�_�O0�^��`c{�pP߲Y%��\�SY	�[�%ڟ��i�w���8?ve��+��.u��b�ՒØ���o`��T���`5I^<0
z��@Eb�Å�(9an����V {b�w���}'�o�ב:��i�Vi˃�(k!Y�4Β�[�6F�c�? ���u�^�4� ��9�4[J7S����Nv@�N��HY�I�I�\\k��1yU%:F���A`����YR�h���L�F�k}~|O"E�����# 9�lRPu���̩:���:��k̆|���+���:�y����-:΍�47F' k�3�7̓�2`�x�E�d0�kUװuN�e��@�h�5��[���������M�����R�p߶N��A��~qy�*�� fT���1�Y-�-�(pس�[$3��VEV�ѥ��,Bv����.rYx�3�@L0IC*��i��&ȼ��ӛU}̹@� �A$u�u��br6$um�>����������g�Ao�jڱӊy����ɰ�|��y����e�,���'�E��U�W5��ϸ�-��L��6y��1kM��{�u��� �
�?�j�z9����������w�9L��?A�9}-��\�wv��H�����Bh��	@,k��bF��Pr�j�4�څ� �;w����kgR�r'�����2�K��������V���a��,j�?kʹ��-��>O��d��X��b�d��Z��U�ͽ��L+�m+0##5Y�f��g9�xsY��m8�9({b,�<7�h(�7^\����p'Ɩ��d�]�ȗE��P%Qʄ��r=Ƶa6�_��TJnX�d�TPBG���K�KjL1��n��q|~7��F�g��:c��	�5^j*�5̙�{:� ��A<�p�P)S�|�HEW'�l������H�F�P|�HK�*g�9
���+���/~hLD�J���5^M����q��{q��ژIp�t1�*�����E���"�N6i���{Q0,� rƂݾ�o���K�oy�}A2ϋiR���DuL��k^8+��En�Y�~I]2��f��v�{���������6	�y7~;a�T{?$MmF��~�#P&�n:,�����%��E��9�i^C�z����Z48��\4�@�n��aB�"�'y�ܿ��J��-ڧ���vQ���	-%s5�S����27_�H�ȝ�W[ݣ[�U�eB��k�P=�� ��}��>ѝ2m|������c��4cTV��	,��֜���nW�b� �媘#�X�� ��\�;�/�ΐ�jc%1( � H�Y �Z# hm#�B� �B�sA��h��4�ۦj��Z��a���8���\�@+O2@oP�)x'$oH�DJW��
�8L�j����y�m�I����M����b�U�����K�#���@����`��xh帤B PbV���S�x��k���c��wm��}J�� C��y�a���e�E�D7��^PX��v�ˍ���bm[�:H�;�{�U=��H��	�8G(�%3B�+k�9���59��Q���'����X��gY���o�";�cb�o�31�_T9����MŒd�K�XJN_�с]��v{���߫� _T���2��,Ni�%��խܪ��l�g�ܒ!P��xx|5�;��H��yl���/����"��f�����煊)^
xx�[Q%���+�&�lV��V,)3[�C3x��S�؉�0o 	��p��6p����kg4R������u[�x�E�N�غ:$�3Pl�;~�o�D�[rG=qZ��t���E1��BB7H� ��"������ u����L���{��|�jv�'�� �sU�}��b�*�:�dı��B^Y�۽���ݽc�(�1���ʝ�Mۋ �������,��3N�ړ�{��޼~� A�;u�ԭM
|�h� �%?-e�Q�/�Yls)�E���
�(���vz��X����ew*c���lr/�����O��j�����2v$���B���X!��{�3Ѯ���)icA/�" l�ٖ2���V�w��Nd\%{mOݳ\�1sJ|��l�����������Xup�R';��ɯ}f7�|R.�g���gLD.@"Ck�0Z)Tn	�D[�lA��n���nT�Uq����F�-&�5C�g��
���2~΀Bĺe�Ahr���Z��_j*�f*�@��l�TZA��6�l�����Yxq��E1#@Θ�옾](�Gu{;e�g�V{�ŹA� k �ك1�]K�^���w^g2V��.缆,��Ш�`���} �l�1
J�N��E.�B�g����� �����D!r˒O/p|&<�:��h}�A�^�Wx>�d�S!��H�{.
jC1+��.�C��</~�\�^�W�c����kk;��V>ǚTS�&��	�k���Bݫ43�r DpY��X�,8�i��3�4��e~��ː���U����+�GI��{j��	FL"�%jK�H&5���I����Z}�,�� ����v�L�R(Նf?�� �̵��l������
 ~��M�p�B2X�V��ZR���DBx�Ñ�ߙ>ӢZ�9կ�Y[VA��Ce�W��a���%�����ʠ��_.P�VIK�Ȋ���ɬ��vd8������ƍ`��!��T�-�5�n�Ե�c�T@O�K M�|��`�3 ��� ��
�{ܔ|��V��R�kP;@�dx��L�[�V:��I���q��t�3�I�!�Vv�vi���Y�o����t��v�r<� ��R4-��ڌ�XP����B'_/uQ'jn��p>�V��F�y⻤�/W�P!a�)`��Ey���$@W16M6lms�6v�E�u��[�<x����l�]#�	��
cq��2e �?�����N}�(hF�In�ƖpF��ڨR��0��yІ���Ö�fYq�!R`���d���Eg|���)�>�h�i�7(?����#�b��pJ�����vcb�ww�&�HL�\` 
����+�t�g�QD@<��g=[��ѕ���Ԓ��f�yV�ohH�i(=8iD-O��(�ܺ�[���N����^�G|h� ���&	��>9�e<Dk�h]� a���{
�Wtcu�X�-�7v���f����Ȯ�<�P��o�-����[��Ц��U�ٍ��i��"�y�Gƚ�"ٱ��g����P%�P�_�$���6���7NE2��i}�P++����
�M=)�m�D�`ObN�'	H�:����w[���:7z�I�Ή� �(���d��g���薷�hc׷7����Ҵ��W�y��1��܉_[��TZC^��Py{��3��_��>Sh " (�P g�^�L^��E��"���6����Ө��
�&�UJ�Y:�~�����`i��]���6�^���r��I���Ye���!|�{�՟ښe�������U�E=c׹��w��E�dّ�l�E3�+*��Hպw�K������W/�t*"���n3����#�{� s[h�˿��^���[�g�*�,Pt.�e=�,f��`�`A���}�p:7�-r�$����1���!T�,U>�z7q6�vˊ9�<��!D!��
��v�R�D�bC춷�7�u�A���$�p@�~���Vs���(�Pw��Q��yN:'�P��0F�6-(0���,ߌgB���2F,��Kjn��N�q�����y�B�����MB�����t�8D�����6o�`c�5i�,XB	O19W�F��D�o��B�l��Z�[�* b ���ns�l�.�C��=����rS���Uԭ�+�zzb%�Vz,Q���SV�u���P�X��:x¿ï��腇*6|��hܫ.s�vF��s	�-���HQ:[6Id�FI�ѢM��Jԏ�k�^diƵ��%�lC�Ұ����P�]��~6��t<���.ޤt��lL�a]�R�!�
��¼� �ƌ�o�B:�ld�U�Qƅ�����q��Ls�j_P����|q���V5�<�30ȋ �f���A+Qͅ} $�E�Ճ�<[��*�aT�²pn+��o(����Z��'yUdhI�IOI��b)5)�j�|>񞣅OJY�T4 �o��R�H��B�.�,nl͎6�&2�&?>1��P�$u��50���� ~���C'Obu��2˼Q����t]ū�H���v��Sh��9��2h�b@R�At�Y6t;8E���O^(nH����D5���%v��ͤp�=�c[�t����=�������{�%, `��N����6vl��m�xúb®<����m=��K��댾qLP�+k	r���4��ҁɨ������$z� �(E��Ü��sK��e;^ϑU�Z���!�M�]�B�����
��ώ��i�V2����ß#|�>ω�&�G�mn���6u�l4�|�,E(Q��}��rPۼJ�5��;V���ص�%w��Ʃ����@��Zk�d6�_��鷪❃'O���tN�L��Lf�� �<N��^��~���	|0���#u�Z>O$��(�Hx�]��^2�{�!��:y��!r�4����q��;�޽欒�y�(�"�}#:R�h��zs�D�M�"�#�B�������3ia�>��#Т�Һ�W�̄4��h���,���,(��C�f�
�lv�����9�f�.�_a�b�d�R�T<%|��Y�cĨ���=������?�O?�h���?�O	�1{��110����\]��鉽}u`�?��^�|n�?���*�A`g	6D�ʝxZ+�3(蔩+/5Q	�4��{�K��_������Γ����T<�=��f������|Xi?���� Z=y�����d��4w� �ȋ��T-.�������{��Z�b��UAUsP�������Zv�:��7-��h�J�T���b"w$
9H��,(���H����F�^ЇE�$s��,�OznW7��&��3/hr��;�u��4��9ɠ�=�5B<�Z�SpU˂�WJ�[��y�-��C؉",E�hA0���LU�U�� ��<g��Ѽ�����4AB�EK�f��R�j�y�p1{��g�[ԭ�P�������֜�z${�M� �[�<��h��5`���dX �s9���BL�$�ٔ暖;<[lA5ԮM�t	���AOӖ9#�%jI��L{]y]*8+���`�n>;��������D*�oX�\���<�3��d�����^`O��A������0	l�nY�kK��rUׅ]��Љ�|O��&�]y<��4���z�}��+�j�Q�7���[_Ѵ>yN�g�'��w�OcX��THOp�IE�JP�m�l�����{;�]����9+�H�m��M-<ݠo �Z4I�ܘ��='R��R"dː�8��N���7)�T��A���{asSU��$��;::����{1s�S� �ΖH��TCF94�8(AB9�Ǫ���^��y�����v?3��ѵW��+���G�-yQq����ȑ��(ix�� �b�U�y��b����1��"�-tM�
=��+������ȥ:5�B�y-0���K���1Ԓ���ws}��u	R��mӯ�����5�@���!tUy����+�5����p�ٶ��;`�l�w��s�rϕ:z-��[H�CrA���[I�z��[�B �!�)TQ�'���$�t!W�����48
*�kVN�-��(��3��yl2��W&Jב+'"i�}`9��97�)% �Yl������B�fE�T�6� �2q�IcY��Ƀ��u�ڸ�;��4�b^���~
�$�Q;�J.�	X�y���h��^wI����[��jgg��
����L(np��C;>9��"�X������墭U~��l��h;�\�5.�c*�dN]�T�V���������0&{��B�9xbÞ�w�ۥ|H@,՟;Ju*�	e��U�;Ո���}h=1N��՞dJ�\���z�g��ԥ��Ү��������)
�7]��n��J�� �RB���T�����|m��V\�*�a�v[��X�H��s%����	���;-����~/�Z "~�������f
�{�����>����ƶ=��k����o~xj���k뛢�jGÒb.�_E����{{�歽~��^���>��[ؗ��7�,}=$0�Nk�����5�5uu0!�}m{�%�ٌ�q�&I�>�_���,� Q�����X_�T}��	�Z=˯��</���;���7Е�����P��X�
<9;gk�@8Ո{�g������g�@L`ڀ8��L�
^Kqj�--Q$���m�{27��D7m\:��c�����}/����X :׹��Mڂ���
�,T�N? ���Ǒ��)������ǿ���BF.J"�Q�3)�"�4�4KK�\4]H�K���E��n�Ә��Pޑj��S����A���g5[�KF�
���(q�9����XH�/N���t�9���t2�<0���oEѢ���`ɼP�u�V�5Ƙ_�Z�S�/�9�;g�����Gg�����!�SQxj���� O�,�E6���\��,�u�L $s����*u}���]`}�k +%���TO-4u������6���w���F6\�Ȥɐ��Wb /�o��wNO$�pFW:+�(ҿ�O�1&��>���]�!�2������.�U�U��j��P��7�Ͳj]���ne5���	硲λ\�QIV|��m^����~hM� 97 :�١�&m��|(���2�T�l�h����7�.����c����f����h2�����}:8����xmH*_u�(C=�+������񢥭�i�A�|dɠ�u��R�$=Y�w�J�h��.��2zcC�A�� ���!����/����  ?]]��o�c[�3a��T��Җ/L\#��>o�y%c�AE=WVA��p��Vh��y4�?��\xeC�����ۦo�l�|���Q���f�Xݨ�a��%4��(�Ӣ���
�p�q����9����8��G�x6���f�|6.�a�Ǚ	hc ה�e:���@�B�0(�]Va�t�z��uҺr�̕����\t��PG�ƫA4[��I*��cs�5h?�U�Ԙ���@4R7؇��^��3U�1q͕R��R��pZC�I �UyOP9��͕du�J�I���R)�KX����l���
�&������1�B#tT�j�.��2�^A�����U��lo�xܨ8s@@���BcG�17���.��B?7*���.��\�D�h��(=�L�ݫj��݊�ȹ1��P0��ʾ��V������Y*�b���#}���|��ÿ-Sw�ݕV�Uj\��I�9M��`��I��ř�-\Y�d�sK��~-���z�=+;Qw�Y|�@+UUYl�kW�3O|�^�֞��;�ijn��a��
��0��D*�P%���yփ�v%a E)82)�y��?���c�k��I<<��f� T��:��g2ٝ�{���}��m��V�g���A��\L(���~}�����?���};>:���)X*FR@�sC�EQToYs,��9�΁�KV�G�{̏Z�,unbJ�ThTL�<��r�	[�h-AU�[��T����`�-��}�x��7:Ɣ����/��s՝
"dj8�@�Jz[��`q�ܥ�eJ�����j�j�W\hf=�Ra;�y���?���y�b�9����f]�ʒ�Nz2�O~�dGd'�W�g}Kz�y�)��I�U�H/�*��.��`R8�a�7຃��?���?mo�,I���GD^磌o�`fK���R�_���H!W+ >, � ���ޑGD8]U��#���jVvx���e���nnj���-G���D�}'�j���}䌣�������O�}�ڤ��or�|s%��L&�6��Z���r�)�� ���D*!�٫����=�^�W!c�'���X�I�M�)G��(|E|Ʃ�̔�� ��;��mR|��cv����SfUy���V\k�M
���
��DZ'�a'=c�9>[L��L�����c��V-&R��10>jbZ|�S�����zّ֣�}�I��F�ɌS�s�}�)�֗v����"D�ru�v*�:U�-[��s¡��0�F�9�|��J��k4k�Cg��Y$K{E� ��r����Iݣ� W��X�gP��veC���|�|`2lX$	�]�Y�xR%E�"*n &:���P��ۭ�'��5��O����uc������k�������?��_Xwc����)jԮ �uw}W���t���(� �IG#Nz�v�+�J3��ꢊ��=�9Ja�~E�bM������.��`���t.��Qe�Gު���4U �(�Q���!�Ū�7�*]��ߋb�������L�sv�E'ǽ��ҹD�k������%qёh�X�b(�d�I(�3[3�I�6��{���`D#'mR)9�iNH�s! õ X�C�z}��"�^�>)�$�o�g��ٶN�(T�� �w<?�8S���8wb@ �8�{L�yP#����5�#�z�F3ȸb���g�XO��<�X}N� 0��O�|ql��bXbe�zF�@H�Q������`O��ax�w�(Z�����M
7�m�� ���#]故g�([Y��큨�GJ���[�mn�5��	",��d$Q,�^ߩ�����[�� �I�R�d�7w�D֖���6��'e�P4=d*�E=P��)�NmA��������m�
8j��������S��6�1^��_'=/�����C��)�1��p�!�����������.��æS���d�*��i�%�+�K�F��arvAǤ��"v�x��@֝\ۗ�;/ڴ�Ӝ�+���0�:g�<�!j���h��l� ���zr�Z���׬��s�r=אTƀK'0�?�վK�2�&�{�r�k�ʑ�,�8>�KIQ���v�Yn���l����u�G��+�kkW�vv��Mk��A��do(@�o��������X��A���0 m;x���(�6�Xo�2�B2��`H�u5�w�Ξ�׻�sv�猒j��-�W�z��s�36�Wm0\�T�>�M!�m�-C>��x�'W�c}�טFC���xF;�h�^)#M]7I�oH����X��v�S�wa?`M�I�k�\�ۈ������%0pԆ� |��P6��.�T�XmeVE�Zr�����~����Rͱ�ɞS�m�zH���
��#��Ҫʩem�h;��@`�����R먨Y�VM�e��iM�^�)J�g_SH����0|���G��c؅���[oP���%j+0"�G @꿦����k�zx1�({�HW�`���Q�X�1	�@f=e����P��"pa%(SY�e-�Z�|$��֧~���l��I�RD�ߌ��#���#��c�AP���/VCeE08[�uV������Rd��3Ɇq�8�q�g��ʘUS:����zk�Vev�
̭�A��
��a#f�b$��=:q�����/�P@3�C����,S5@?�|�Zso%�랤����8�uҠ���<��9��?�00�fuk��)�a�0L��"����u�Ϡ��S�;z]LI4S]̤�-��i -�Ĭ�g���~�YNmX���"B�i�!�ȘR�s�|����䲯hR⊱@��0���ۏo�������!8�X���)�ص�� I%o�i�^�,�=�z�j�D�`�%��� ̛�;���w�s�y��h7�]��k����;j#��H�,W����<�%_�eO�����=�U�����&ё�����F�4S��#[���i��r�|b��O�O� �"�:}j�T��D�FO.������(� ��isQ5���x�5x���V&*�<j�N�T�~5���؍2F6�fb�\|U$�]Osa4�$ +sn�zbl"hS�4�`7�PF\�{au�Hg̟��(��"�Y9n�N��="�&9�ꟃ�4��#k;!�MZ^��E�c�������\9kV]��Ƶ=�7}�5L��"M5������ϼ�472o����O�ZCP��l��:6#�]zA^D�:�����ċ:4>�<׹]#a5:f?��g~b[���򷸆�{����ϡ��Cnv>���'�8��g�Η׸����x�dE��Q��3]L	&9?���	��T�QNqi�%ې�ϋ���<��F��g����=y�߶j����;��e�E$}�����Y{�o���~�����/��[l9�߿���������~��?�Ͻ�T��m����i��bM�'��xr/@���٘e�y�fb��#Hm��Ž�|<���E�t}r��O��z,��.���^����[>[��u�P	Fܐ��T\+;(�,r�F���կ����(�X~�?3���g^��S7K��j��g���; �4�1l13���f���t��Mʤ?;�?9���lSd�OT ��	C����\�'u>���"cs��Ge�HIC@XW7� �3�V���0M��O��U����E"���,z
D�����Tm��6�5�a�9�L/}2�O���3 
y�����AQe�E/5�)R� ��o�}B�`�i�<@HTE�F["9��\Ԇ~rY�U�^�d)���̖׈��k�g<���z<��9��0|��Ӥ�4���� �k�,Ւ%e4��1���H�ȜYͼ���Y՞0���<t���E�*�&%�O��=�U�LNݯ�d͵.(/칥8�����3�ƥ��߲"TxHkQ<
�6�n��;���T��`�ZT 8իHV�u��c)X+����v�U&4$��?tkz:ԟ��)8$���
�\�TĬ��BK��'-t!��5׶�����If{E�&��T�8��zj�o/d2��)՝�N�q�3���H��$ղ�N���;͔97�]��{�X[$��T��4�u�فP\"E���hv���SR>�ፙ��B�skq�+�����4��:r�'�uAa{�\����M���6!�h�Q���+��U��v5���T��g2�f��dvG0�gtI�Y3d�1�:� �i��10c��� +�2}��EqN�[lp���5��<��5�pi�u�M̭FuZ�1�ٝK*?�~�=`���x�]��s�E�������HC��	!6R���R�QOHG�)u�MR19h6�ZN�>�K�.u�_�
�9E�&Q��������J������0q.j�\�a�i��Z�E��7���묬ii9�z���������g�/��g���s����Ի_|�=xF��s�x�����>��G��'�{��G[ 
�����]:���vm^��ȎhO�1�!hBT<�(ȀpG����{���Y;��_�zI�6����ho޼�~��@�_��_��~O���(A��5$�s�@��v�1��Ͷ..p��go6�.>\ip�︽��+����#�:K��u������8�,�g�P�z7�'��3�(��
ij�q��k]7#A�d��)��ҁ���݆z��N�$�4^�#w�����!�5���m�~UP�[��T�m̫�v�ⳅ�h��q����
�۪m�)��u�,�� QB#���g^'Ē�QY�[؛���Z)9��q�w'�%�X�f���Př��{Qu�q<1X��g�޵���tcˑ}��%��^{G��A�h�-;SH �%0��x���%~q��}B"0��@3�9�±��d�t����Hy��93��"^'�m'6AU�3a��h�C	R�KU}Rܑ7J��+����ԼA�%�`�(zrƐcL�W�;�T(!b�NN\�^�y ���P�$��D�G�6n��
n/��4y��̬��=d����U�_(��G���h���6ma���/��jG|����Xi��FY�+�Ȋ�\j�۹0;�V%�7��u�R�֊�av��#�B����H~�y��&%�����%OQ���A�0N8��T/֭���&��Q����t�,n�Vl�����vs��hvW�{��˶�=�}�q� Y���B����8� �49�H��W��S�U��)y}2c����C��qs�T{<�&��@ƍs{�> e�-��W�W��l.������q�U�Z��Q��nȱ�O0+�բu���cS�����)���{K�0wF->���E��6���A|�9qi^_(�v7/�����+)u=K~Ur���.dd�,�)&�H�X���zV�+��)s��P�n#c�5vk����'����Sn}��s�Z�e������It�WA1
��aa�$�c�ؙ��k� 
*XD7�%�r�JZ������ĥb�q�������ДWN+J�� 	�!wڬ��<��s���s�e�;�n�_�ܛ}6y���dV$�*��C�����|5�N�[e��k��PNqvςk���g޼�f��G�����V}�O�:�!�� Zf- cƽ|��*w<���+��� ���;m�`SjASk��������i��Q^�0/�\8�f�����]o;W����ӔЙI��P.כ7?؛�o(���YP����]b�߽'�B�Vʽ؃%�!n�+�{a'ڝ��ٴ�����mr�s�e�-������;���������\���@V �z��t:W+�6p�L�Lo��Դߪy��ݩ*��̝�Pn��g���2f"���;]2ۃ����N(�����{�hR)�y�G�K��
�(��#�����̋���A�ѳ9ǅ�*���k�����k��|52�5��ݜ�sP��HF��#��x쏫�������9[bd �{|`�I����Ȗ�iVe\	���$�]�l_1��k�Q~1�^���䇝��H�E��#�j�P���dj6��Y5��u��T�vr�#w�I't,�����
A��T�t1�KE�*k�G5䵠��[�^C۹P�̹ĤB2�;&��aVO��J=)�u.n�� ���T[/1 ��[I�q�&ܣg[�.���f�A�&��[������	�hF�wGe�n�����۬����:&��V�-�bϰ�03I�c޲�
��.H��H5��Z^%3(U"&�{=��5ԩ%"$�ԲcA=���UdwAQ͚��Ԃ���Kz�U�B]׶Ial���1�F+Bf��0f^ Hq���pFCݪ�į8��i&Wуwy�ot��^�R���Fk}�0�٣.�s��$��[v�Ao�)�jy $��,�\���ۭ����}��o�����_�ۇ2a���g�C�i����K���1a�Д��
��5��ip���su���<*!�qk�9 �dH����9���ҰβT�p�;yt��.I�0��|0.l*�ID�i�AQ��5)�I ���2�@ga���;�0�l�|:�gE]�P�	I'�O��U��wG��8'���b��B����N�`+P�1��j�[�Cwò7 \cSX7��!s��8sU��EA@v[Ef��%Zg��p�e ���s���M��u0���
�R�<��dN���A2��A�1�"��~8X��:&�VFv/��y�����_�M8W��̭���M�FeJ8,�䈙��*B���M$\8�*R���V�'殮��]1�-i��E�����sk�}Nc�]���}��t�����>��{EEǓ
ֹ�w��\z�\t��%��:A.�`r*h�"�a� ��<Z�y�V����3rD��Oj��k�yog�ds�h}.���۽�p��G��#g{U��-��g\`v���JV��
$�e�)F�=�ߨpf�?^�\%�۷��B��hZd�j�#GR����n�*��3g5(F�v�S!j��/|�N}�G�iV1�0�����|6�IP<�_��\̿�~j��8o���sj�:���@���k�Ώ��f����x�K�%�MM��;�F}qZzo��z9��N��'�E
Ĥ�kD]��L�Nr�P���<��vc^�|v���qn"b����vl��l�c%��XZdK9�T�h���ՂM
<%�u��fr�)䊗�C��*��e��o������?@�
�A�����Y.d�)��l^�Ns�j�$|p0\3X
(���_ �'J�r.�A�$ Q3y���>��7)�� �d����Վ�j�ǲ��|A=@	��6.PK^�?�S0���p u�s�Qv���5�Y��+�ӓ��Q-��xb�t��j��5��jǞu�mA�YE@�wK��RO�Z0�a<�&�'�%�f�X�a.�� )t��a��/W����ؠ�X�ۼ��M�w��A�i:r��Xx��]^�Ϥ���F�]��L�c)�����ڋ����k����� �D����ɠ��d�ޗwt-Q��$����xYI�5V^��j��K8��]�򵌾-^���I�B	IAR����7�3=�{E���������<Y�௧�2&���R����(��>o����fgϞ=�HYC��
�����&iP�+;CL�W���-���@��/웿�+{��/m�{Ae��;8d��-��ӱL��mn'�ٌ�5��>R8B SD��"��T��a7uɓ��,i\���H$�9�P���(xpEGDA���y����bD���HA��+�h��u��4[N*0�C1�� P/��y��)����q�,ea�p�Y�x��l-s@Ys���1J����37�26+(�ាW�����g@fw�UD�2�rW\��rp�I<��� �A��P�A}�)gEh�'i�}0��W��*p/ ������ۜw?Σ+'���*����Ξ�xn��w���n�ڣY�w�?>z��Я;�
|x�W��f/��S��5���_=|�q�\���9"1yDF�����*]��tϙY�#���lz&N��C`F E��J�\�:�<���̥M�;:8�r]�~�A�kNn3J^��S���e��'�Q1��0�[�lxc���,ݮ��l�v]=c�%6������9���A�M��N��h�o��Z��`�y^|���L���T�t�ζ�"5����c�$��Y����N���!��9�\U<�V���f�,hRqm��\Y�,� ���9,i|�y=��>sVϚ�G�Tg��Ng���-�.����^����ހ�������;	�DNU����p�ϕ2�!�A�t6�"r1�L�%;���s�/2�97p졀 ��W������$:�����)��x0��+��p@��D��3s��h,�gg����F��8>Ɂ���KD)��_��,fX~�os��7��MN'"5�����'"�r��	Uf�D���:?���T{�1ɋ��Nv�J�=D"��z١n
��-�ǘ��xKL��u���u}�S7��Ϊ]�T��]�pe����|���32��;���"�j����^�f�u��>1�����T���H&P?�P�.�����3�m�o������J��@�����+9Zd��6>un���X\��Nc��
�Do��� xD��T �t�8���\�^#ޫ5H�N��������U�%�Ѽ��sA�v�(����i%��9�@��J99��!R��mqm��3L3}N�i�0��������M{_qG��Sd%D��6������6XWW�
��w�z��&��3�e���I��i�s`�Z�V����w��Es,����Yd���2����]l^�(l�M�,�r��� �2�wh�j+�$��Z7����k]� ���򝫝;*�= �O��T��B�)���/�/��/��=�ԟ7^��x�ۺ��b@���#M��_f���=���io�2�o���bxo�������{3ٻ{(��6wW�� D%�mBF�tl��IR�µ�/�z�j
���:��а>)n3����]���dP�]5��L�5��,���ɉj(JQ��`z��J�|�ӊ �&�bKk�c[��~+�q���~f���;@����������S�� �b(�g�}ԥۛ��l�h6�f�Ã;xƨC7l�oh�t�e^���bolDp̑B��?m��I�퐓�.����
@���� ��XΉszz���,C�ۡ��m1l;H*("���'���,�hW���;{��x�����ʘ����y�փfڌ:�W�S�DQ��X�@'��>�� ���z�΁訩�"��٥4�d�s�E-���.G��i�)�����#� kf��)9^ �Y���)1���C�:IR�^R��sP6�t
IxDYy�\���6'*@W�-��Q�1;�_�,8�ľ+ �xm/�������[{��=�{ε��� ��tĴ��~��)TO��^�t��I���hy�z�;�����X���l��/G4~����I������g��.�����vȸ� z�v�#�~H�K��M
�$���$�Xl'�똝
���%��˃��#Ʃ�$���^���½N�#Nu�_̏Z��.��N�����֞C���=���� ��7�6(�� p��:�et*��Om��_>h��+��0�F/��'��mR��j��I�J�Y{������&���\
0-�kQ��;�	G�l�m�B)�}�Z���.W�IfG�{�-��6P�-Ӽ���Z`�2��7;�Q6ux����<P)��m� �u��¼[��KD�pA@q��:;����+� �O^�L�N�a��@�Y���ű_��N��9�$[�^B0S]������j&߸�J���@�s���dO��A��R���Xs��\}V�lr�Y��k�?`Мz&�&�F�k���vp�ՠ�=����g&����wۖ�;�}�̽裩�$��� �M�͠����2��HM56����]I��A�AJї1ڋ}4��a����sxν��g���HQ��[p��� �!��b'��צV�*0��٣�}�wuhl�%���1Ze�NK$E��Kվ$�A���=�bQ����f�c��X�-"rQv+&���}Fi`0�>MN�[���
"L[?2]*ޭ��G�m 0#Ⱥ* �v�4��~�%)��.��(7���˗_��_c�~�}��7���t��G��@���x�=�=V��T���U�I�Rv�#��������~��#RKA�CY��
 {�)&[:��������V�S�)��Fj;��cT�5�s�l`��qH ���r�l��젋i��v�N��U]8x��n�:��g[]�&�ƍ��#lsv>+�R�
�G��&�u$�̟Ԑ8�e��~�H��y� �,��?둛ǆ���]H���0�W��"�{C𨨬꧘��\��ρ��=b��)��AO-��X��q:��,��(�X�'�����P���p86�٫�0�]�{ϟ?g���@��:�;�w�>�7n���ݕϾ|������k������L& ց�5+�#���Lg���e��'V�[8S2�s�M9�-A憔�]��2�;��k��'�$sڐ��C�˱��T�̞�'�C�߲}�zI��7�H��Q��H�ȳR�z̭�U�ĺ�B�E�I��S}?�c�׾���܀v&8d��O'{�?�����=ج��n���<$�a�+ �S+P�+�%�IǺ���._y룯0��z�������@�Oͬ�!ռ�U��:����V<�vꏿw~�t�>���|�O��_k��KT�<����Y�|1t��ĸ}���;Ug6�M���d�a:�JD�W+���l:�׃zh�<�{g..�j���6gWi���Ƃ6Y�z�v�Qͤ�����I_M��뵜��zи�����A��Yu�!o���D�%��,N^�� �)�14S�<��锫�Bn�w���.;{$<[��P�[������;;C��}&�cQ�1{�����Ȭ)J���QOۧ�v7JFd�h��l������P$Y��U[P��Κy�
�;-մE�S�� ���T�{��lQ���݁O9t�	R��>����}LR����'r�X|%(S7���0��H=O�}���Y ��I2%]u�5�z���t�u- ��q�xn;W���.uފ��10���Y�:��|"y�H L�9����ea�u�>�R�i�AM��{�A�����P�`����ծd��_߰����&�� ���y��ށ���~Cj��a����Z���byv��������!u)1/lpJ~?A�sP��ޱa��}`�lq�fՇ:OV�o����|ɧ
��4�v�ZÃ����M�v�0f/�S�T,
,�pN4�D�3/��H����残�y�#
'_iH<t�������7_i�~��}��wd}k�w/*Ț��w��P.|,N�=��gqh��dGr���?�*�
��d?��Vbd�`�z?��c����[>/9f�8���LƉ�~v'���1��N�P�,S6��8�Ң~r.��#A�����C�c���~�s�(TV֞*UvIY��
�o���C,�S�:|���zokY{���nC��g���B��咱O����N��n	�ny_ ��N�Ll�!�(�ON�ڮ
Ⱥ!�rz!����w�1�mMdb`���ܼPO�r��65���qd��=�	~�
hz��%�Ώs� ������Y�o�kzvgϞ�( �e��S��ov��ᮜ��LଞR/�����vwbo�<�����<^�<+cvg��mq�n�7�j��&���>!�6�[��*t�5�FD��NRD�u�	 ��R]���.i%�����\,�X��e\����H���5pf5���0���,���׍+'k�D?�K/�.��Hq� �Ź*nW�
g��h���b��0�5f�Ԟ�� �g�R:�ןz����̾���{�ϟ?^��K�Q=��9W���?y��?����:���r�5ޕ��/~p5�#� �-��/��!,���j�A���0	����
d�]�7�%]���u��;�qOK��H�`^l�5��mԨm<���.4ڮ-�Vd�"���[���.Dp��N��/�Z�3V�7����>�۵^+�ü���U䮚)��� pZ�Y򀲟���3Qcj.P���b�c�w��р	����β��/��@����y�<��^Z �L���^������ ����T�v1�����$k�lk >�i����q`%�z��0��t�RY�1�+�H�p��J@Q�ʺ�������|�0Z.P�Λ��h�c~P�?���Zqt�l�F�~����Ĺp��7[�W���?<׌��խk����H�d+�����td�����_$7�L������c�iw����-Z��m�p�����Z7�q�z/�U�T�����C��d�A�2}����S���U��,��~�8�ގ�DA���^/�J����^�}b�b�Q1nؓq<��a9{}�I"�2�Tx�m��\E���OX��VkR�y��`���vU�usn��ŭƬ��ӼTLT��#Y����S��R��9�II:_Dѣ�}�I���B�H%�T�����ݭ�x��^�,��g�]�))�p�z6�S�:��nʈf�p�+:�`=�X0
���'{z����@t�z�zEK�ѝ��3�Hg��O���>��w�h^p��=�\�<�B��M)II��݊��)d(�P��KzA�!S�%&�2(���*a��� I@6���QF-�MZ���G���	�"Gm4XQ#7�A�R��Mk�е9�{^���]��@W�>�.Ȉ��'�6Di{Ei��<f�v  �,E6�:"0:�Y̓2�jȺc!'
x뫲�MM�X��"�5����F֯�����^]�ٮ� �	L��5�����C&k�-�qs]����u�ke� K`E`{$mT����&)#�u3e��${�fE�������[��67̮�@�8��˹x�j��H<[>�4yF�'I>
Ի�I]l��H�GJ��<��-��e
�[E�ݩ�1�5H���ò�1r�S�٬E<(G�ӂ�d��t�q�S=`vlveΡ���t[�f����ٝ�.θ���uլF��(`>&���,P��]B����g/;��s����>��~�;L��i��Lf?��\ljէo��^��w�����g���/qAG�=�|�
�\f=Z~1 E��A�yE���g"�}X�Yjm��Yi�y]����[�z���#���g�s����\]�H����R�.�Fs�un�α�:2g�� -�������� Z:C�d2���N�L��s�<qo��Fuq�X�<* ��X���j�G"x�4E��k5�,C�g���ڭNm3j�J�#�D
>!�xz�����&�R0]�ޅ,zoi�����}J�}�-���H1R|�M��,���G��܈;�����?��=6hg��9�R���s�z>��;9�a'%��m��5K�P�2.���l�������N��r�ͤ4,@BeK�Yw�@��H'ͣ�k%A1��<�����q��G��3Y~��8Ùo�<�=Y@�:)�ާ��x�2�������0��z�A�t�}5q0�N���e�{wb��<j�����p߇`�@�CL^L�uJ�>?��_3A�gd�YR� C]��;�T��us`&�,u�ӑl�W�Β�)���p$�m_���n'��]�ף*��x���^Dɪ�\�}\�5n�����s̍f����](�������p<GM�����7\4����L^��	���6Q�`��O� L�|Iq)IE<�t���ŉޗc����6�i궶�wv]��wh=n�
�eϡrΡ�k�u�.I�vN?(�= !
*�=C���<xd���7j�R���=�M� �H%.*U�̥.�����w�נ�mxm����kMiW��G�W�E2�7�~�y�Qh��S��H��B)����Q\b������0�JiԚS'�"i�T�[W�S�lX�Ź�g���X:4��%�Vn�ۭ��r��o��1Mec`�o$R�n8��#� ���� \�3�^q9F?o�x�(���,#��^ۦ̡�>S p۝���{�~� ��P�c;PM�ڦa�Q�r�2��	�X�8��6W���$g
����D����܃��W�bad��0��n���� ����h\�w\/�	I�e��:��]@YX���M'��˃��7g����8�����3��5&Fh'�0/�I<�e����)QO����'W]LTvJ4/8J�B#��O���M,M� O����h�IGEҮ|��ͭ}��}�ꅽ|���%��M�G;==���H�e���(g�5�95KǴ\/ a)�G�c4����-��y%�o8;���v�~�q:�B:��������p|n\ �������>14]Z�F~l�����w��lI���5���$�p�6{� 2����
~?���̩�(F�-��)��
VV���0��M�Bj"��mM"Z��m��[�I���;��{<��%)q�g�ӝ�����Ǧp㗝I��-���~���ھ�۵X��˙���qfe����Pq�1l2�����d jѓ���-3`_`��Yg::�1� ���V�[K�0͒�~8��Ԧf&O#kU��Rȓ�agI~�N�E5T��3ީ���M���XEy*T���ݼ����yPxhR���dU^�)hif�?���Ȁhyʧ��=�~Mp���$�:������H_��{���\  �<���x{�������� ,ڎ`pE5����6"�X�`�(��D���X��SW�-���
��܃�pwؗ�R{�P�a���lPڱ�o���=գ�Ⱦ�����>��h��{b�,Ir�X����{�L����P]r���,z��/�p]��r��J�Y}�������vf�o}}���l�O�>�����wq�y�]���P��u�*c��(�����P�~~�^?������,�_hs���E� +J�K�m'�G������I͐�?��؉w�{�b~6%"(W?����Ԕ��{��y�
����0�lo߽!Ȣ������X\�裗�>2�� rv(��q�T �t"(��y�\Z����������=�`.7�e�3U�v�
ߨet���9#]r�A�Qw�DZk,�a׌(m�"�5�8{�P��A���v�Y�qC]_�pٕ]lS�:��j6IWF�D�\l|s�����˃�����ӱ�*I��r�Sg�(/��A��_�$�[{�?=��͵�_5�c���l�Zd�UZ�ZlLtx�P��G�~#{��4�6�;�|f�![��L{IJ�#�?�����y�!�6~���6��2����Cf�'X���������$e�X�"/pVZ|��K��2 dȠm�͂�:��@"u �0
g���]�v��<�_,RF4�S)j�5�e?t�xY�k�F2S�It��T�M	�Y�֪��s�����*	��G� N�ߘE�$����h�g��.�ʎ2��TW�&�u�4���T�̍R��h����ؾ���j}�5"Q�@P8���8ܒ�E5s���!z���pPƓj�@�d�r���&�Z��pJ�Ήt�x�T�H�P�87W����s��/�/_؋[Χ��2�'H�&Q6�*M
�y��J8����]ʿ��|�*��������Ws��y����k��R�)U�Μ�s�1���wlq,���Q�q}�� ��D�x/��?�:S��@��YÙ��`9F9�����u���QZo����q��E�G�NB��6��I�
g=%l9���b�xr�R.A���@6�k�Hp��u������D���yt�Hq-)T�� ad�:�1e/Y(c�z�eI���y�L����=���mI���2'����V��J�������C����_D=S�k��x֞�"k�$?Ϧ�����X ��A���,8Ȥ�N�T�.�6���j�H4��j���`.�8p�R'%C���8���&��s4J��G]4�^s� !��]=Z�z[Y��4��P��~�Ϣ�ʻ�O�zv<ef\;��؛VL�L���=�2�Ȟͮ��uJ=������	,���&��Ӭ�����,���"8�)�����ww��ژ1+�':�IA���0(���Kh�����Ʃ���n~~Ro�Թ�L�{�=s8��G6�ɷ�v�ѯR<I��<�W�-�S\k�X�]�/�@L"�dy���};�g������Ld�<�0�{ �d��� }6��s�!)��[;�8��
`-~7)�ґA�����.l���l�m�?���mKչ�(��o�̃������Nj4@�����u��蟝L�t<��	$�
:Χ���ӁBs4`-�,'�)�H�a彲�f,:o�
�J�À'V��rK9���0Y�2k���H^X�㟘�j�'bS]r��o��B�i;WR2�X�&P����!�YlVK'�,���37�T{��9R�I��h�D�:�4��D�g����Z�4%��S���e�`�IԷ�JoGOE {F�R��ͤ"�'��<���H[I�Z�b�/�����8���=�;FI8&9�q�'���M�irN[{�3��\=J K4�����p<�֩)��Q�t��;G����u*�Њ�aε��.8�̂�{��j�h��^� ��!"�'����% ������16��������h�&�x����\q J���cd��lVRt�������E-��(3V�qW��M��\ֶ1�|�?�6�ݻ�N��Wj�]a�g'��R@��Ũ݁�y���ꋯ^س��I���
�,���}���	�]���^ϒs��BG`g���X�|z� �'�ԇ����RW!����/���k�-�Q�"�F/����ŭ�h�ͩٱ _ ���-0����ߛ?cF�ʒ�Yc�i���Y�]�������<��؎�I��nFPpa���eF�kmЬ�)�_�_<;��(�C6��-k����//>ĳx�<��[��JlL��e;���|>������#>J����S�5��@,�A�v��9ǔ���Y����]_oق�md��z��Z ��!ʅ��!n6;R���@�����y��p�4s���m���}�^��؋��O����=���tHw��`J��N��Y2���S�� -�m@5Cv�M���s式��0k5��JqS,D�p���*���=��0��I��������يf�j�S`��O����fD�SVYI]��θ��88�Uh��G�]�={ml7�C�}�/Q�>��&?���p"�M�k�L��!J2�������V��	n����B:�:��4 �@��)���騨��q�K &�"
��@]���L�X��C`G���\E9{C12�pG�@$|�,�)[�s�eѧ&����Z'�0EP�ӣ_�+�'�3ƗL6_���4։ȯ�2�_�}���@ͳ�
���}��:W;���:ߋ����s���u�os�@�QD¦�\_��+/����
[��?43gc�¾_D��ѱ\���'7l��^���͑��Y}|�k��Qςt7%;1�g��H�JIx��cA��6
pL������������5��\A��XC�ɸb�Gǈ����:qϙy��U���CԜ�`�G9m���Ƈ��F�� ��Fq���?�!�	����>�kU4"��}��R�D�,�c�@�~��O�N��A�g#E�3�R��|�o<�['e%C�Z�t�2����'"/�����ONd�P	V ��>(���;fv`��Vak������&�|�uQ_01�K�)�n�2Z��em����--���1`�h� <~��T��>�Y�&������}VF5@��ٟ���yP��� W�g�@�r�ޚ�ef&��uD�8?��
��ܳq �7�LƮ� ^��ʪܯ����#)�4� 8�ʱ#÷r#���|�t�� jэ����%�di�r�b�D40>2��fʑ@���[�#|��{�ol. +�!7�NQ�L�������k{��$7�1Y��Ǝ(1'*
v(��X������YT�0����N�b�ǆ�X�؀^�5Q��W�R͚��>���+]�� ���g�`~�<��P�6[��!��&g?3������?/��?�v�Np�<�/tq���|�x2�A�Lsˀ-�ݹ2u�A�o�)վRW���
���1z�E�9�=�iWQLz��h�[=�[�~�T#��*���,�q�Y�5�뤆>+ּ�w���@]�}99�r��b<��E�p/U���Ә� L���������W_��/�z��F��}��9��;ޭ��{}{E�%�k��o�������O�\1j�CcV��$����8�?��}��?��޲�N6�?������T�E-�R ��Eʵboڗk},?����D��DU`�U�`�ۭ�6���=�0w��߻g���q��c���z�N?��� :�It�?�3n��'f����Vz3	M^�<K �줋|D0)�-��6�Za�M٠h/ߢ�*��������U������i���1+ssrJ&]o53�,��]����N,�`&Z{v�P��N����f�?b�zur� dB�K�NF�4�v�J��#d6��A�T �O�i�(N��Q�s� � @����)Y�����D��8*3I<AVV������)�U��fe[M",���~�$W�5�1P'�֬H��I�ş�_�{Q��L�T�Ϩ�a���a�Zf�ںvv	_\ئ橧���QȜ���G�TKay��;��^��6AVtO6SI}>��ET`� @��uIh�7J��	�,�g;{���+Fg " C��/��W/��m����@�UK> �j�1ב�j�E$�ȧ�],�}��D�-��ف jg�$ZW�!���Ѿ�T�u�m�|Mԇ'����8U�C���G*��{���B��FM��?�Uq�`w��繱���3<Ls��+��M'���k�W�j��A�u�ޅ<r��E�Cj~c:P7�y�ԛ��JX�� �Z���xZ���=���`AO�=��rH�xq��n�{};+�M#H1���4���MA�YQxr,�xFXe�Pl���̳;�.�A���8z�@�C��i����yO�#l�4ۈ���c�xؒ.8�s]S�n��;�2h�eͯ� eW:����J����9UIm4�r���vh��1R������w6x���ڞ� u����ª��6NR�V҇��H@���8g�B ���^�g�aJgw17f�:e/�U2�ڷ�����B��_��|����灬9��gS9����Ӱ#�Q�G��Q�!R�1k�T�d��,�_3V���m���]����9�;�kI`��|Nf�s�`�'����:I{��H=�JQΏ��B�+�;�3ׄ�PiHtgXD=!��`x�5Խ��m�b�ۙ#�?>�Ѽ3G�3���ψr�f��{q�j�/��Pn�S�{�Q���v�;��_㻿��~�_گ~�]������3�}���ݻ��@g��S� 7;����>�Q�{��o��o��~��O<��ǽ�P�]��w�����^�v�e-˿����/��{����l2�.�o�m~����] w[ U��h�K.?d�ȗ�z�w�����=��������^��gdh�?�U���˽���-l�����'�M���������e'� ����ڑ�H���ys����6�C��:ͣSی���*wN����j/7?��/�Cg}*u�f�T�]���K��%ʑ'�Y��Q&ĕO��T�����*5�&�̠�AW�Z���fQ��8ܗ{eTIG��
懄����s�%_��m��Ġ8w�����,��)�;;ݰ��� ��-����S� 2������Qbhe�Q��k� � M�������A��ԝ��)�Q�9M�F��xw}��"cg��61�"�c
6y��%���s|���\��w��a|Z��0��؀�YpGUs*GLo��M�y�YQi���n��!��F��}�z�7����W�+{��}�ŗ��/�.F�Ʈ�B��k=%�7�ow�F��duѰ|v�1�5�vfq�2�M�fw��Q���7*!yG�ttn0Pׂ�Աpo������b��C�#+]�1a�����e���	��ϣ���Tg���s[x�qG^�'|v�>�X�I�ca��ļ�prC�+�\��jRzXݲ� �]�À�L����7�.`��r��Y�p�Ej��2`t�<�7=I��,L��U-���{8)��XӪ�G.zd��Z�Թ8����,9��3�\i��z��o'U�k�����*�
-�*�$F�x�����T)�S�=8X��́�?�Qr7�s�z�!��� ��j��F�=dv]�=Ib�0|땢�נ���y���_ߍlr�������K������B��On ca�G��+�hd�Y͑���ꧠ���W��@�� a1�GNͼ�kС�J8�5�Tmu�%�o��Z�t�?u�4%J����F�N�g��޳���������xo	��9��U'7�ES�b]�)->��e�iy�K��s�/�.����p���M�|��ɰ�Z�4J�q�٣��|�Rؠ\��嘳�q�su����r��Mu{��e�.1M �������ŏW�g� ��9�B�|���Ξ���_\U�L��՛* ��渳۳�Q�/^�����������׿��}��]���#���D���� 7�H!���n\w��۵�|uk�X������2臛�X��B}fW�����H���s{�%�+p�]�E�"���\;4�g#�$��U��\��Ȼ/v��� �{,`��y�"�їױ���Q�t(�Q���K)�rS�8��F�������������������R���k��&L��);���y��=�r��GY� Y��im���h��� �?ꭦ�U�~���.N�:2)n�gS���ѹӄm���p�}/g�enn��2|
���KqZ��0E�g}�9ᬓ���w4'�h�\M2�Λ^����bJ��Z�W�f��^�J@��C@fAȢ�U �O~}���t���ū�#pI�o�gW�t6��oP�4qSx�^��r�z���7�7���dͮ�ΞP��%CzN̞1�}��u��GA� j'׫�k�*C��~Jr&[��U&` Csu���p���+f�Y�3����-�)iP$�:H�S�b��2��8���4����WT�����+��)�Jl��������
����Y�;lK����QO)���5Ѵ`�^�jT�DH�5���,�*�8y��q��I0�S��tjhy�긅ڞ�sa�$vNg�[�7L���5eYD�yݍ�z(s�)SoDt����d�~Ԗ���s`|R0��:�g����l�.�Y��EH�V���4[��5U`���i��gg�{��i��Z/��ȳ�!N>�y�ܼ���;WGj��'�k�KP�Lb��>�5��e���Q����ñ�}�D��5 �T��Sn$���)�1���<BS>��Nߥ�r����pP�p�ٖ��>�"J�.�yZƋ6%���:G�,�� #;�k.0Z��~��Č�Y��NPio�g�������kܠ��� ��}���`k��ZPԚ*�
c�NQ�����~x��޿��B�l�|⦁G��#5YdÖ�:�3�j���,.���\ȶ��g�?��g-nZ��h�gw�?�k�P:��?Ǯk�'�῀*yiO�O�?6,��O_c�Q��������9�-f�_���MRaƧ�R��\r@)?Wl��P�q�=�j�g~:M4��.w0�D�@(���%/j�� �e|��FG�i�3ٞ]?g-,l��4��n�>6q�R�9���v,�>�(�?h?&�����9ZG�ijwn�Į����~�����_��対-�GO��=v��×/&DՖ���T���%\o�vswm��K��Z1���&����v~��M�z��<��q�:��J1���ޡlH�RO"�{,J`R�YgkԌ�;:�������y= [���5�r��.�=�);���H���Wt��{���~��-{3�6�����D��� �M҇c x��w�u~p��j�&9�)׻�l�����ԾaOH�=p*�rF�|PXu�Ꝟ9z9D�L�~��Ʌ�06��[���*�ȝ|�ȈB͐48��A�`��b����+I�b�P��aG�n3(X*A
紧���H�meڐy�=�)82�x�Jɐ�S�f*p����ˊm�0��+�h�������r��Agl�ʎ˲R�~Ԩ(�&�D�:��m �47P+�~�q,��4�����J���g���Ы�<�sW?��L7)�~��*�K�劌���Y%����a
�)u:yr$l�Q�3�������M�1��3_����,����5�����SWdH�Q��ɒ����<�k*-{��օ�۫���W�7�?��~cϟ�����n�vD���֮�B)�WD�N�¢����	��Pj�E�`���1^��wzO^�)�"��jo쫁�1*�.ì������P�R�N��{ӕt�sr�\*H����72\� .�Q���0�-�Z���O��4/�������y��"���XJU��~�?�4�/1�5�G�)G8��>�����E{��q	$�},9�i�x�����z�����ҩ�?tiQ�Z�.a����"����;��z�t������g�9��٩�M�N�&�Q�-��~1b�+#���i���`�g�+���9V�`Y���$��\��K:r,<�$�5hl�x鿋�K<��#�7���i�x �;��=�i�ӎ���UW�:<����aO۹�?�a�=?�?��2ٛ7o�O��޾}W�w�ė7jv
�?))^��&���Q�>�,������j���q����S�.`_u�SĵDHⳀV4���Y8�m�
����cA�3@�p�ϩwɝ�O������}���������{a��g��.Բ�";�c��˄H��v$8�)Ue3��PrJ��u� R��b�n�{��M�ly���n��2X�c����ŏr���8��E9�3��#{��/Zb�=i����+u�}nv������}����:۫��ށB׳F�Y`�+�ٜ�`(��=������1��A��=��7��I��,?U~�}�t��SpAd�M����=(4C��%:��v���R��t�7���eXSs*ߣ��>G/�� ��ڲ�vMfњ���m�^1<�j�������h?��}m��6>�o�\�IGfi�Ԍ��	��,��}*�(�n�}� ��L��	Dv�أ��\;gG�'ʮv�(��:��A��U�;�e ���My��5� f�Y��8���N��E*݂f�{
�\���B�MU��w<��mpL��Z3�x����tT0�tz<'����,���&�۵�X;�kY�}^�Q�p��@g$�
�]�deC�
�7q���1����ut`V ��+?&�G���+�LI���.:�=o�u�]T�&
~�#+g	��s��z�a�^qK?|z�K�]m�|��ө�!�6�� �	�Oj���=@�=�T��e�6�])�^�����n�u���P[���aoU�⠆���хZ���o鬱�?�����X}����)-6��������ذo��'Fz
Tl�CE�)_8Xw�W�W��ۿ���~�`m����a�ō,��ꛎ��p���t�f���o�B��$���XN5��4�KN>�ը/wdh�N�:3AÈ�j���k����m�iB<� ������חltpI�F�=n���+�kI�l������j&�r�燎	�R�Y���Q�1y�FY��÷؜�㐵��rR/N�ccOmX�_�T���6mbM�|<�� ;U�>��e�����:�E�ʂ��;��S�T�+=��\�>��9؎�Wjns�#��$�э=�ץ>���ȝ�g���;`�J^��N;��&E��?��#��s�yW9ҳXF���P���r�3L���7��������^+�56@���A���P$ן���t�Ĉ$688���7�cqT˱^� ?�xAA+������#�*�v��3}��쒅xIn�9>�K'�Ί��ESu����g�P-�g��
����9�^yu�Î�*��g�k�Tt@�5J|Z_��{;�s�����z�3�^������ų�s���y ����������
	������������Q�
|Ꞝ�}������_�},`Wʱ�{V:n,�*h&�|�[��:�r@� ^΁��599�8��)-$� � ��m~L�b��I��U�����Rr���<� ��2�5�^C�����ݿ?С�}��3��Jc{S��:�<<��	$uk�^[,Q8�ϓ�"{0q@�CHhg��A-��iO{����nP6�~FX��V����p��C�2�T�l=��� n��A�_Pqs�Z���F��7g����ܔ�}��W��~�K�����˿���֮�;܎S���?6�3l�g
� <@�2X3m튼�Dyv���w�^l]��;�dP����H%GS4#E6lʢvC��I�=d�fG�uN�D�#�R���wf�G#��\Y�8kKs3k�� �V�"�8�〦�Z<����"�E��2� ��U��S�����pĳ���y؟)�0n7W[{p@9��R����Px0C&���ve�(�v�8�DߪG�m���� �#�����P;Lv�tK�T)�0�N�y�݊A��U���A���� ���nE?h��$�&��µC��a��ź�\��	J娭����5_�8�_��bq���D`<#dn���9�e�.���n-�_=�dy륰�U���$w�,�����>-_f�o'7�)О&d�o�BD����'&z���EY���_�Ͽ��������|CІѠ����={I̳jEع|�fʽ��Y)�P�g4��������_�Db犍����M�.���)VGƛA��M�+��M&��v�y�0\��ю4lݜr���6�n���Z�8����`��3�nN�S�^��n��Kea��Ũ}�s$Qs�4*��E�ڋ�:_��,>N��}M��d�6�m���/"�u48K�U��4�y*-�ϔ�tA�	,�֨YHrD�� �u�!֟�EZN������&	�L��c��x~`:׺���C�	jy\�3�͟u�WW����N��3ߝ<u����>�����.k��%�V餂|�ug�H h;M
_<#S�t�������桘�t �����ll֐`��5���r�'�߿�����8.�x#Bd�A�@v�.�u�|tA�l�p����r�������ީs�c ���gq���� �ۉ�O?�ݟ~-6s���tN��
e�s.�~=9�]8�^�.�ڌH�����.��1-�*��k`����?���3Q[��%�<�W}�n6��D�lCP��u�s@�B7��e�Zߪ�6"-����<�ӟ�
�U�-�� ~�/������R��c�`c��[\���&ߗbOM��Z;���E���6���ph���ɥ��*[���4hn������WϋSv�u�����<<�������f����Ŏ�H˄s��t$w�\=+�d'�8�e����4G�	�����{>�G�=P;��#d؋�:�e� �ph]swsk����#�r��DӃ�vd�G~�W����Y��[
xlx�1�Gg�ף�EqJo!ұ�f�e���C�� Ϡ������,�FM�q��#З�;�$�qm2���@��;�5bD��(�[ b�Ty����K#�ۡ�)����Dg/2�T�Y`�Z"�m'�Ҕ=f?V�Kd�Ge,��HM��{i/�Xqo���A�{Z�f�Z=�����#p�(��s�q@�H�cyN(�Y��ݲgЗF3�|�f�r�Ӿ��NB(ndPCX��=������^��`
mo:��k�K�IM��L0��L|�i;��M�(��OaL�|���uhtܫ����T�ϵ�}�k}���ҹR/�27����T0���}JN�n���[��h^��27uG�t�i�m�Y��#��>g9�9k����u��)�J��ZFÈ��3R�X����!� ���9�e���8��Pb��t�;6��b���vg_������������b��M��� -����7�����R��x<�{N�s�Q���y�:�QN=o����	��B�Y�i�dB	Y(�Q���V���]e>Q�;;�Ȯ���������a�+`�z�І���}�o۴j�ӬJ�6�am�Ù��T�X�Ԫ��[��f}E\�R�΢��������f�ߗ�u�\?��8ܽ���z�D#��1�������6g��϶��~�S�����8H^LN�`���XK=����:VE4rsZd��p�>�y�>sPV��>d�S8cU���@���[���B���W�ר��f2{��:�4'����
jDa�*���8~���={�L@n�����9.��FC�l��˖�x�Xcp,Nϡ8�FM�ɲ�L0
�!~�32x�����gc{�q����Q��ֿ�f��`O���b��湯˚.����v��[#�]o���-i$!0�sYKH�PמG�j����h����jT��[�%�r̺��n�'�����sI�<��4��~P����uK:h:K���Y�A�(��x���v5���|U�dq=�︖Jwco�e���HjN��j�Z����}0΋�;�郱��q��Vy���cq��]��U��I#�M�}q-Ѥ=�~���o]���
~![��G[��un����Q͕=wV�~�Z�1{��M��%F�5�J{�G���Q�Y|>%R����%���ΝZ�p��{�m�Z������u7sq.@�����oP����Dq�Es2���h?>������Ï�?|i����b>��U�������{�����l���޽?��;��6R�+ ���D I���%d�T�2�	�ծ8��t(!��H;�/l#�ԟ(X���<1k����^�xn/_�����IǹDͬ�Z�4G�5\û�T|�����m�V;�vd ���<��no��w�}]���n��\��~~,�sπ���\`�1�jE�;��GS�'�zdf<���`-���^+#NQ\w$��i����=��X�k��y}�q�<x�\��N�z�i�`���!�M&q��r��Je*�c�F����!��&�&�A�]kx��bl�%F��,��af�cv��lV���wa�n��Q��N�Ε�.�{qJ̞���@�ޘY������V����lT�5�&;P����d�2�q6ܓ� �ʞ V�:�a�L[�:֫��T�]���^��؞d��֫�w��,�A�5i��(�+�+2���=	e�s�ư�?�K�5j�X���p���ZB+��EC�.(׉�������W��&C�;����=]?��@�r����E�}�V����0������#g����l��pĊt������~e���~��R2t5�ب�Pn�I��r���3%Lon`<Vu��ҿ�أb�1Ϭ�b��N���{fdms��p�	�S{�G���
�����Gqe�fkNC�e�#`(���@α��[V�fC���b��8rs����K�o-py���z����l���]��-�[s�d-��dm�}��+s��m-�^\^`S�s-��Ź�����6��k�P&PW�y�ہ�;}�!�!Q�E�X�i�� E�g��F�ђ*��On��<׸u��ǦD=F�͡o��:y��K�~�B��K*�EP��+�1聧�$9�Q���T�`ԑ�C=���%G���E-D�T��"s?������W���_�����ߗc<����FO�ٗ �VRy�\f{Z�g[Ly3){��8�F�)dv�Y�C]��^%CXM�!+"S3�g�=���gܨd��L���8V��|�}� �oW���boE��P.��s`��K���E����J|d�+������
� �����j-Ր�XƇ*H�li	j�iqV}oiw��a���}Y]~|�b`89�0k�.��倉^A��P1�(/Us�.��� jE�ͮʧᴸ@����{�L�ʜ'�������t�������ü�9{���3L�ď4Q�(��{�{�nm�F�E�g��pMX�p�@1;H膣�T#�M���������`?�~m������?�������b����06�
 c��N?�IPO�^V��E��rNԦX�᝚*[}p�S뚍Ag]�aOe��a �[�P џ~��^ ��T��qO��kF�
dT������x(~U\�rG}Ty�+63^������{ُ�������/M����_���ڷ95d�Q�=e�}a'D�2w�5���GN�HT��\��hs�%>=s���r�X(��!��p>4���v�T:��䊌S��vP�]�]�\��M��Ϲ���|ʤH�q����_����ho�3 \�wX�	$�]��͝7�U�h�=�>��ḁ�7L��F�I&;B��I�!*qﶶO
��@^�5�~`�NlX�L����xG}��j�S(4C�y���*�zw�'Քk�3�L7k��Y�� �5`�@�y@���.0\�=ԛ-3[�����@��p���b�M7�y�V)�19K�:�m�0�=b:E�@�X5�s|������ЎeI�=2K@]�4�I��pf�{���bgώ����|�j��f��5�x����n���ͱ,]�Os"����h�Y�υ�	�8�#�~Hm���ݷ��/�����/X��/~��ѡ�!�����x�vwd�k����o��V|3N�5��Y���CD�2,�}�g�{�r�i�JQ#S܉�|;AY�0Ɔ�NPKD��7�'Z�R驃��[�n��0���v�ӯ�d��Ks�~O��=�<��������B!Y����,��p',���p9y�������Ǐ��x���'�|0���W{D��N`r`4��`��+N�)����x�%�g�qy&��Rc��2��)I5|थ��R�~i��:�1hs�k�(~���z�Nhaf�<�S(ޒ��s�ڣz� ����������2��C��AE�G*@͌T�vGQ#���U �lE�T_��#��݈��Z/4ݞ_*+Ң��,%<.قld�@K� ��"��8�ǲiI�L��Z��BK�5z�����n��^X��߻�'@{F������;�;�S�}��2��'w���J���9x�3���U�{����=ٲ7=��d�2-�5�^�-J7Tm��������gœ�]z�̂r6����� q��d5Gɝ���}ft�"�P���0�[D�v�w���~:��oR�r���|�9k�ȓ�t�z~�9f\�`{�̬-����(�?�7�M����b9��?>�iFV��KvǙ���XU���-��G�u���F<��Wvyq%��S�0G�;귿�����������i��������:u=�v�u�u~�G�F��|GPl�
W��F�����ݩa�}�2�� �V.��ޣ�!�oo����}�|mϯ.iS��nmW�����-P��V[��p�|���Hl迡�t9(����T�{vuU�������*��/^�t�V�AﲖME��A�qR�N�nZ�s�C�������BM��蔭$�� �j�1l:�1�pVu���0��6J�ŎT�_#p�Q����>��'��0.�;x,��f� J((a����"ˊZ��!Ӄ��g`	��������AcO�=	�l�'K�i��;���Aj��g�Qs7����Z��zO�R��MJlHR�u� 3,�Y���5Pwp�<�=��� k����ؔ��g�mt�g�A6����x��7U��\�P��
ۋ��Z�t٪P��ߐ�
���s;��YnXS�;x>�<�`M���i?p_>w�j7�3��~d�T�(R�2\Cv}���16�ΪY<�D9��$,��bGL\,d�޼~S97G��1J����������7��?��{����~x��YJ�n�Ӽ8�d�,BΓԔ���.��Nj���s��F�0Kb:�1#F�u���u�9	���9A�n`mWw�����R�9�ZR�x6����}��(�� Y�]vsf��'�Ki�p�\�x-���gw�yk��N|�t���qz8�5��s>��ù�zz��7]"E�o��������+%?������g@����΍lh��+�2��=^�g��գïK��[<ww^_>���v��>�-����?�xn��GO*p��{d���� ����D'*K������asv����CAh����A���n�k5�d��,'��ރ�s�ۓz'!��ƙ�"/��R��,֪���i�*�����A�ޅ6,��ʉS��j�z�]�-c�Ͻ�m=���ٞR<�ԭ� ܥ=�p�O��s\s"��b%/t��d��Pmer�`��4��v��Y65�S�,�%��O2ehJ�u��M�� �͒��c'��e�lyϣ@�= U���A-/�5��	��@a�χV�%@�>�yj��ȭd��}�� Z~GEr����ᱽ_�j��-N=0 E�+p0�&��	�[Z��wms$@)A^�.�h$�gp�t�ՁLއ�Ƞ9�ϔ�5A�'��H�D��N�����1|���}�ͷ������7o����z�3���[���������O�������S��
R. :F֓��f�Ci/����W��sR�:fV�DRR@�g).����D��сiPt|3Ϲ�&f�o*���既2�7#)���E���8�gk���îY�o�P������>~��Od��X��KG�,�s��vsAJ 5�0���D\kfq�s�m
�ݮ�<d�+��<�z�眠E 8׳2E��=���aU���3+��(MݙY=�,ԣ�keoH+^�;xb@x���CĂ`ƜBVǉL��@���A�Y�z� �~vG�m�sƦ��f;G�_Gϖ�CA�,�u�:k�ɚ��:�Ƒ�T 0�oJ��٪�[���t:6�N
~0��c���	�%D}�י]D����S���j3����Ǣ�������轵��^;�y��  �+f��`�J��LV� �!8���j<��r��?��]���\ySh*
 �w:ߤ�Y�ۇ��jT����{���/�,;�m��u���}:8ӹe�b�I.&0�&8��]�d)x���� �{W��W����[���~o����l���o짟>r� P�x��޼���|i/_��/��Ҿ���a�r�(�̔>�oCç�*���z����eI4"�~�	{�U�l��o��� 	}���"���rD꺿�9P��-��z���9�֜w���#�� t��Q@��QV\�r :���u٪�8��k=ɀ����������l�����J����OˉO��<�Π��X��Ǎ%M97`C�Y�)��H�1'�s�䶾����+�ZG��ܤ�D72\�P�1�Z��q�w�C�GT��;9�O�_7b�Y�k0?1#k���� 	�ՠ���Q�f�ExἠG�|���0����vR&�XlV[Q��6�{l�T�q������S-����v{w�:[mE�IɃB����x@���5:�����,x��Q��h��Ï�|iT�_Ԩa��i�%/��E��|�K9��3����lHv�Hm�C����,�Pd�-I~�1�-���b!�����9@D���j�1�E7�9�Q���|���"�����]���"�*~_�w"A=�;�l��y�7�"X1�bv�� �s*�)�l<�t��j�{̒	gm�
���&Ϡ�܌g�: T��!_9h�+��;����`��NS�`�I
 �I?~�c�9<���r_[���a%�ϥ4��c>���^_����G�'#S������B;�qkЄ_�_��/�����W���|��A�u�����������?3h����U���;�o�#� )��`sh�y�X���1^����8�j�	bX����Sh������G�=b|�Fo
/���?3"����?2�fW@<�z�3Ȼ۽�և�O�w�P>�Ķ���,�lǙ k.����3q�z�̱E���j���p/%����H?�);�}J}���8x�G���VRP��U�]%�<H�O C��|PdA��wJ�f��ޡ�H�G3��� |��~���w��Q�~�	�����d���J��X�������`����{�g�V���� �:Nꛉ9�f�E��꽠W��1�^��͜)�~d�I�_�rj�+ PC`���z��O�ㆾ`���̮>lʴq���źt?��S(K{p.�|nh5��d�b��"j��N�#��4�֐@���;��`�$[J��:�� zu��_W�qR�YEO�h��cA+�/��+"�m3es���B�9M��5Vt�z��m��Ee��E����9�!��������?��~U����Q��n7�4D�/_�X��W��w�1����+{�}|�HcQ�\�%@Į#�4v8�'�k�	�����E[�(���5i�p6s_�-p�Y���EO��7�8i������O�u�����O��SЋ�����W�"���8����8��G[�O���{y�N�� �dOx�#uH�ߣv�7���.� Yy�Oƣ�u�.������K��<	XL�`!�ߦR^��r��ζ-����O�i��i�{��C���Ȝ�CZlK���
�)K�"�uB9}�.�P�lŴp>���8k�ϪI@���ng��}�<��1��TX>��L�{�)�O�˵�*�L8��"������o~k����?Vg���k��,d^��=�ڲ�Lj�l�����X��:�1���J�C��c��h �[4*4��`��Y�R��CY,mZ��&��-xB`SwѾ0�o�}���b��G9q}̆8T`=�\�>?(��'��x��ɜ�a�n�Ӊ"Ty�ނ�v�Ǯ�ӡ�E��ھX��Ѳ�Tˌ�!�6*n�d͚��"��R�Y��bL"���f�81Ҳ;��ذ�V�=�< ��W�x�G���.�c��]Wv�in}�Hz �N��Ә_���\bH|�z�PO��jq�S{�����^� i�$���B6��zp�8��!�qcW�^�_~]}�o�����1ϊ���d���������o�S�+��3�*r
GÕך�9m��kI�	�.?aT����ʤ����X��=/�y�3Z�����@'��C6�@W C(d��B�wPAEd�/I b�:gp��N�d?���j����]����|��+�n�N�XJ��lY�L<�	�W�@�&�)����h�i�f?&�Ĩ[F���I��P�jtv{44�ܮ8��:F�á�dA'K^p0��'eU4Ι�OR�Z����{��"�k�Ǳ3�S��������.�DVs��"��X��-^�ٕh�B2�թy��(#4�ܲ>���wbT5��A�j�[A���L���xh�,���HB� � 3e^l�c"��cqtkv�����*�g�G���d�@S؁�q��-S8�7�cFr=.���I���-��/�A#���GL��s��� Y�k����7���ϡ8��B�@�����L2z� �v;��������P�����������?���������?�EQ�y%ŗzc�7��T8Q�ϯ�!��n�1�P�VPm�N>=�D�Ơ��F�fY�"�}7�J���U|���q4���-���z�4/��K�{�9ui���/'�X������=UL޿���㖗��<=�i��)7�!V� vj�G(@����dO���7寓���r�����=6�jAQK��i��`�w�|v@�s�y��k�H>K��������G���9�m޵�D��cĕtC�z�e�D���G������;�c3@a�q��b*�9�@X�xWB�5d~A8hƉ�y�k�ڬٓ�k�D�c�m���g�������'��ǟ�ڰU}_'Mp"k=i, R5�X�I8��\B�;�����a0
r���]��-C_}���u�G68�v�OLq��i�|�n$l$P%g��E'���`��&��B��y��Z��Y�\\���ؐ�����F<�����@V�������y`�_vm�J[�f��=q-���`Ѭ�;h���*�v��X�:���{��{�l`|�M�+����g�/����NM8+p0�,�c'@;�Ջ��F
/���G��9�)�4H�1�җ�,�9>��o�Jn�ʀh���o��ਨ4�,��2�
���ƽ�2v}sm�޿���߲_3��S���8�+[��m�=�	��֢ k�c�[�T���.�[��O�^��'ù��)tys�_��o�ψ&	0�5W��Co�d	���'�pP����D
��O���o��^�z�f���������{eG��YdPrV�R�!%���򍚸�(8��YdZb.�-�z)��'�9vB�/E�R�=T��(�V��JI�q�+�̍ �%�/�$qsV)�B8W�}mZ���Ƴ�s�yH�{&�͠��Mj��J�l�u�} )�}��mAt��a�Z�~ä�Y���������ŶDĀ*w9�M��\���e	�9С/շ�"�d�x{#������)�s[�C�^dGs؂��9�@/�߿X��`m���\3���	,{�� @翡Ĳ��Bا�����YS�K_���s�m�'�٣P�,����Р�G�϶�f�J�!�х��{����?������_������Gn*RT��ё&Ɏd�X\9��n��sN��C�'��z\�����}�pb�w�6��؊��d��,j�l��ɚL�����-������>�� ���Na�_C���s�C��'~A̅��ʏ�����R���gѣLV�^K� ]ԼwƊ5�������,�,?F�� mh�o�&C�G�+�/��Z�R�՝O�,����F��e-� ��[�!/.���'k���p�:�U�LݤIᣚ�&�^J�����8����sXJ7srs�����
���g�Cl�$�A	ޕKDg�hE�Y��3#�(�m��ٲ�=%�,�#�H>S��������B��� |��g�LO�$���ѵ�O�����,��S6-s��/��z�Ρ�O���5;��Px�ާ�A�s�^��j_#]i/^�k��xM��u8�(r�Z��+���{lN	!�24��T�����s�~~�Nt&(��0�-�=A��u-�v1Y=�+KУ]P��5�BC��c�j�H�ݣYS�
{%���
�g�lJ<���'�O *��|:�߃�ce��ꖾ~�"~����Y�q��=�d'�$|,��o`�m�yI��ى"Ų2ǁ��sL؈*ջ�L�����Wo���w������ގ�vu��=3�3ORqی�<��7�Sf�x�
i��zIY��+d�9�<<r�&��)hM]���Ą+��d-�1��@l�-&1��c�x���IA$=� �suEa>������,������'����A��_�\�4���ן� �p��}���@�~X��D��n�'�u���rH��z�Kƽ�`	ssw�����e<01�����o�S�̒�R{���B�6�m)7fe�6����E[��Ū��=���Z� �T��1WP���k:8�"�Adyx����q�A������&�p�h:�����}+ '�-�>�p���(3�L-����0K0*�&E%ĕ����pr{����6�"A1nx>mx�Z[���۩�4����7���m����;uIƱ�Į�� u���*�s�J]Wu��'��Wk;�s]����o+�����׿��~z�	�����ꌨ�i������y�,�DD)rwHhx��㉀[�����H̶�f���2�Z�������2��n�\jW4yc�;�j��g�#t��R<��b�h�6]���>� Z n��8�}Qyy
f��E�Sj�$-���\s\g�B�ܹ5g�<|q,� 
�7���҃q/''YC8�= 螪,j��N��gW�����|wϓ��{%�Y���A�1��r���&@0^�ya��_������y��dI�A��6��>��k>.�jC� �Q���r�E���Yp��Z�Y�.��h���m�)��^gT�d)-AZv,��2WX��0>�l�4����r���mP�rYs��i2�c8�YR،b�$uNo&�4�Y�^�c(�6mNhR�S���@�.�0�G���O��T<{��L������8FDʅG�#=�%��:��x�rR�q����VV@��v�ۼ�O���,Ns.��jΚ~��o����'M[	-06�7`���'���<� �1�4�Z���ee��Q�Zi��i�{�N%�-"#|�Y�Ĝ��Ԕ���թxf��� ?��n�Oʿ�.��p^�DԤ��^�g�TS�{�c3{Ѓ@�����V�eX�U<C��6*�AB�;�A�R�5�F�\���O���?ڧ�C�Ad^V^��؛�,��b�~2���Y������=c�vv,ƽ�i��\tҳ��Oj�Z�
NO.O����]��+KnQ6u�L���=К��Z�Bs
�2�Ϟ?c���>]ӯ�؄�"��C ��� ���6�����[[$*AO���M^�;���B7�Y|s9:(1����Գm=
`!S��aD�(�\�c����=���1[��I��F�	�?z7�p�=�H�}��WH7��4��S�;�Z��>[�~��u���>����= ��9�a_9��XIY�� �T֢,>c�~)��)���qmw +�A�~EYhh�T�F:.2Yc�*ٞ��1���`�x�kqľ���!�� ˴�QIr��V-(�ZJ�%}������6	���c�S�<gO��λU�؁�R�)l�a�>WV͙z����#����k�ư�v�,#��6S�|ń#�����W��W_٫ׯ��[�
�pt�?2"�c�_�z-5���+usd��c �P��Oʤ�|cLRw�y�}�Js\��@��^����-3�oƗz���f����$/�tjNk�P�P?(�4��{�O�����Sa�b/��� ������Z�t����|5/a��`���n,��	 �hrl�m������	����ZKB�+����C�z�{%3�~���Ł��4�~x�ݽ<k���Th8E]F��I+˓���,��;�5*�%�{b޸��s<�Lj������sI��Y�a;��5o�Kl&���wzoF�ˤ���/*g��r�33���b�Q�I<6�;��,�u~�f���FR�2��u�"\T�}��fmԖ��w��!-Ur�!�aA��ܞ�Ơȁ�C�4�g�[4�a����5 #��X��1Gc�j,�k����z�X������S$�DK�����ԃ���b���9��m�$SY� ��ù]o#�<A<��e���50���[`�T��N������ ��������@̇��35�����ˮ��6�(�Ŝ!����$0���L�T�i���^�Ee}���5{T<sJf|Mu5��B�E�#�B�r_?\Ʈ���(�A��÷��Y|���f�x�F�m�-��`gf�9_i�V��Ӱq)v�|�!L0+�w#�뺂��~�����~uEQ-�t@�Sdu >�E�xP�S]��ʈ�v�ȴڬA5Z|FGe��F�g�>�@HЇ�G���v��$x���6@�+� 3l<�\F�it�M�b��Z'X��(�H����*Ⱥ��vV*�Z��ن����j'�������F��zk��҂J��,�2��;y�]Q�դ��0���Vi�6O�</sX����`�]�1��#OG�}�)�P\2>��A˃@��M�la{��xf�|�*A!���6n-��Q ?��G��4{	��I���l�dld��j_Kc�$j�r�Y�*�u��4(��^lVZ�&y�/�:ͳ�Q�Īu� �1ӄy��@����� %aSi{Fe*���8���x	�|�=-�Ɣ��#���"�M�ɟ��K�:���4��̜�h�ٯQ�`�ܘ,�l�=������/��ӥ�ߵ�x����eۣz�9t��<�����:�5/���Ď�PD�.��꙽��;��o����6��Z0/6�Y������_ط�a���{x�����V��Ym���cS�Ml��(��J�#M�b�uX5�����0�gc�ގu��[���~f�1Le��Y��!Db,"��%�0����5/Ԏ�9�ȃ޵����v�]G�Q�}8��e���� WQ��'�O��5���+�'M!Qn��6�"���;���,��֜:�u���x���.��3�i��������52^iu��Ꮱ�U82�z�]v�2Gx�w�o?:�#�Ə��D��|i�g?t���{�A�@��1Kη�{�-|�Ҁ�2ߚ����?|t�y[��wdO���6	���=հ{ks�����2j]�լ��E�3���Zڸ���b�4�*�P�I�`w�s�����p�7�7��n��jc���C���NѺ����ػ���͍��}��K9�@��ʮ�%{�|�DuG�]]\��j��6�x��#��gWԢ�ϭ���7k�[9�Rd>s��n9T�~~1b՚�;�xZ�Ue�w�K&j��Q��ƥ^/���OG��d��/i�j��=�TLd���=	[�͊�b���׆c� ͩ��LMQ -qnO���e|�Ã&�gt|�X
-)s�䙒b�ƕ
�o�j�y�"R[�a��5�&� �n�o�n��9��ug��a�ˤ5k�2'�Lē'5��z��U/A	Q������<h�9�u�������s
.���jT?J�S��6�m@��Y���n3�E33�,��Y��o�O�ѹ�j��P@�s��;��X+�*�͞16��Η�U]�h���"�a��-Fr���[���:�Ú�gk8C������uC����z�&zҼ}vu~YA����ӧ:Ǫf���zuG�r�\@��.l����衔�/�09H�$��|�����>�N��Ug՗y�:�g/�U=������{�T���6���Z�d��XC�u��܇ݾ:�����?W'Ab�t�~K46�~O�Tm��g�_¾ʚ��=�6���}��	>�=�cI�?�v���!���*��{�·�+�	gљ�$9��f��//���3;ߘ]l�s��s�!�^l��D�Q�@�Pi������:��c4D=;�׹*���z��jo.���&8�ޖ��E�!`�N�\9�KUv<��͹�_�؇���m��@*�P��P�ͷ�XR�<c��i{ɹ	��q'e��z}�����L�W��2�.\�z��,���Ʉc���LBؤ���|A&�쌵ih�E���;jA�F����z�%[�����·�J�v�S�u�N;��a����8]x u�bpd��`t@����^���-׋�y0>��>�u=��'�;��#��z]�X���y��[f!���P��N�1x}�mb#dX�O�?�k�Ӿ\>N�����:���^�+k��x�����PJt}g��Wl�=y��F�F5L�9��9�����X<���@�W�%��հ&3`{&!�#���-�#��E��ﭠ��7+~#1�eĎ.�<9a�1u���>B���#����6�&
A�,� �V��z/^<����L��R'��/��ۿ��N�;���G{��-(�*���ƾ��+;�)]l./�����- �
�U��Ŕe�I�n�4O�"�����m�e���hd�h2��;�'��嵧$!4�f�Թ}B���tQY9�ÒMq�.�>����O7�8e��š�V3Ϣ�W����c��-�G�_��XP�J(�D\�=�V��O��,�?��"��\���~����Ex<�/- ��Ч�{�Ǔt������䑥Țv����4�h�5_�o�1�d�u9���|j$%OMʘ�f-Ӛ|>��K����%{���y�蟇���"z��&���#�t�Ge� ֫hX�h�9p\��R�°��~�;E�@^'���V!"��C9-"^�|ɚo���N��E!���
�`���ƚ{/db��k�Ȓ ���PL@�8(�4��B&�T��^9�1���� ��	jIH����ZK[���	T����]� ��q-��ޓ��l��8��!@XJ-+7�D7�;T�@�P&�|��lT��^-j���&s�M�n�5�ò�|k���/��zj�?�gz��2>c�N?��k�O��$�&�s�bs?�ڶ�3�F��9�XwB9��R���p)�@�Lr۔1�<)1�|q<�m=���9A�1}�Y�\�X��� �5D�.@7'�v�%�n
�;.�e�E�ϙ��S����u]C{4�c�D�\Q��9�?�[�{�{��F�Ua�QׁqKu|����D �)5��娝:�,�o��3�\�|�¾x����G���ޖ~qE�[},�B�8�ݑ{�ٶ��/��rEJ�BQ5���L��``�U�����x����VN�M\qm�ф8F����[G�$:�瞊��ǶNTb-��&�v���=; ^sn���W��˫K��ߗ��;�X�T���D?���mNۂ���ǵ~ k��	�:���W�AW %`�s���\?C�£Zu��WQ��BM��zy]�3t��s�_������gy�)����5s��x����ڷ�!��w�@�1��j�Ϋ��IY/� ������ђ�v�͚����=�Ic��&)?���K۟��qQ��j�u�X[k��A� �dW�\q��	��1�a�������0+��}
�{[Ac����*Z�����^{��7����n��v %j��k���Ω�1�\ l�E�s�]����h���y��c2���Tn����v�DA����5�<WWϘD?843��|\������R(-*���ѧ�Ȗ7+_�~��]�Ȕ��es�[S���s�%5�(=�I��xY�R�b)�Y�&����B�L�1�����g:_�����;�����lD�����#���n(D�#�I�I[;v>�R�[��H�%R�z�JI8���k��,w�#�#Y�G>��翴�'y�m�˃�4���g�V��w
��Ɂ��%�i�
g"J�t�S*��yS�����:�^�B��!��X�nEt!^Ծ��4?O���ε\��ٹ\����^V�ܣ����X	����I�O50ߕ��ƫ%��Љ�9����nK|$����&<�� \�@�zZ=x��";�\��k7��N/��.�6K�c-����'���2g��N�m�5�;�$�"��=?��C�Q��l�yP�~V�3ի�-�����^Tg���7��c}���D.���2-��XȻf!1Z7L��uҋ�����ʕ��m���&����G��% 4�����7Q��B�n�s:#l7k������u����:�9��faX�Ȫ�d`�I|�� ��F�?N�6��dZ�퇃�#���횛3k�`A�bl�Y�1F�N�'?�d�!=Z���u4�O�"� J�Q��ݓ#S�A¢�A�@g�6w�?լ ø��C6+Mr�P�2N+�5bK.\@Z+3��9������+<-��Џ�������!�5�$U4��(�p�<�^�<X8bp4�3v�5�C٬����Qv*���^�T�;;��#��?
l�8�Ԓ�κYy]���p��[  <��(#�1��G  A�]���.�9{�0C�~m�=G���K����}i5J�_{�����HY��֘��N����{ `M�_]����/쯾��*0��*߇w������S=h�u�볫ޓ�|��}�Ӱm�!( ¡��:IPp���v��̴�V�k�^�Q��H�$��h�l��]������.1�	�?��\{]����ٳ՗{a���?f�q����#���9)U����'���=� ێ6�}9[#�U�BZ�'�n����/��~�y��Ce@ڛz�[ �-�֬]��?�k
��<{.3յ1p���(�[&n�a_�yroH*�g& ��B�م��5�	�E�&%�5�Q���D�.�m$�|�^��w�g[=��^L� *$����\��ڻ�G�(ʚ@���Y��G��ge�+,�Y�C̵���Pǖ챣�؇1P��޹���{B�h���Q�&�t>a�Y�p?�����<�9p�c�,i�ؚ@5W���=cѪ YY��]r�v���9�*�[���m;k��5{��O�bnL\/��&�ET�����Il�dw���B�^m�F�b�9���=Kb#��e.I�+
w�4��wL7�ݪ�r���7~a��?������?����Pӷ\��޾c�@�if,����D&�w�P��ܜ��Z�p��b���ڨ��V���
'5����Qk�����q=vZ���K�#k��G>A��[�u�x�J�Y�q� .��F����V����p�&��+�=r�mq�,NG�-W�	�T��H��d���UD���, &����!	��v>?�T:��ey���#��/`�T��<�T��HLj���,�	�Z�I�^��\"��_sԞ� T��Ɯ-.��l�� ��UJ:y=���4c�L;�����k�[�͌�g���ѻ�K��s�U\�z(W����F��w��_өB:"X{v���n�a�pqyŦ�ϟ?�#q<������jI�_��	 ����9&W߉:I|�F�z|f %b��D�,j=��82��TR���`�Nq�Z-e5��>y���������������/CУ;f<�uE��A%�(A��QA_�!%�{�8�Z�I*6k���T3h=�ϒl{y ؃jcݠf���p�Q�!.����oKx����t�9N��v�e��_��sh
G9�iul�� �EXV�Lg,�T������	:.�x�Z��<��������gs$��E�)�l�� dp*]�c�S��>GP��{��Q^	��GN�.��V���w��5@�@�R�ke?����͸X[���\s���j;�ď���,J�y"　��q:DQ��>@�D[K�;F�Aɼ������5���� �9�=i�,�zS*5ޣ�����D�ĺ@����s���|m���g����`�����~�/�����h���
$c=��@�8����ǚι� y�>~�ۛ��|�l����R�AwM��m�7�ɔ��oH�h���3۲9K���>��'��������5����7�_�T��YUO��!肌��V�1gmi�QKmh>
	����,��Cf�8(P�{C�j��S^���i��OR<� �1!/�?��֨+�H����E�Ѽș��}�Nަd���lRb�C ]+*dy�j7��E싦���s 8l�?��:ϴ!�y<�7�ذ�(%H�H)�-f�$�������OI�I�G0A��:2W��x�ss��LH~ͼn��������c}���{d
����V�u�efG�6�D��q�I�E0c���� ��W�?���}�r{�xuà��迕\��x�G{=擈�A]�Q�:y��7�p(�Z�E8��>;Ӂ�B�c%c8�ą?v{{d�	��T4�s������}�ݷv�����=0 8���翷�����_}�}�����^�6��gG���QT�^��aH�&�w՗!����7+ �
�_V�:��_Z���R����m�9�@?�<��_UuD�]�JW|��O.�NŮvn/z���5�ѢެE�<`3��r��'�!/��F��W��*č����\�S��F��6�t�Qm���	��a-]��{�1�f�]�P��`q^�#���=�J�y�8�{ŦԠ��s�,�an�U��h)��NP\��	G/ΑBMj��\�Ŋ{.m�e�<8�Nֻ�] a��gݺ��_�j��8U}����`�o=�&�-��ԳA�,ȷSY���+�5��P77wvs����\��#S�mu 6��zY���}�j�h��Ъ	�(S���<����30t$�	�` a�Vc+�@Dw%��P1
�r��8-2�&�Q8l A����M��͚6SS��Oj���V�����O	��~)]��hm=U�B]PH���H9
���6p�ov� +���t<���
���g&���RH�8�m���e2K�<h�$u�O�V��N~K'/4��/�����R���$�y�Y � {"�;�ߠ���Nk�'�b���g~��QٞҔ�J��י�Z29:�*�������u)�-Ŗ�}ų��\�so�L����(Ij4M\鋀��܋�m�Bʰ�����Y��]�kΓ��*�P�}TmS��q�Eɗ+�:fsG�e�W���ñڄ;�T}�r�zqQ���I�����k3ϋ��Y�I~mu̱f&�����.��׹XU�������5��믞��+��^%���W���#�MZ�|̽��(�P�o�-�W��o��,U@7�a��?h��|'
�#�9'm����)ث�\Ȇ��Y9���ʶ+ YoR�@y�;X�n���0��EF&Mk;�
6��6�-�bE��8�l2rh�g�;���\P�a���␶b��"��I�P]&~����\=Ru98Ǽ�]� Hh58�wE�����u�&���`]0��Un�u��x���{��ql_��6���3�4n���ͣ���Α�p�D���83�����U�ײ�CƑ}���i��W��lE�W��zi7K:�GNbV��)�6��IP��a�B��ͮWb~(��j�v�6K@I�6���q�v� �� %����`�=o�l��,�e��D���+d�x��e�m��Yl����9��K[�
��OYUe�,�X��MQ�4�I�N��q`���2�XTH�S����o�P���;{��
����\�XlV�� H@ zb�}`@�����ӵ�w��F�.�- d^zo4�sq���4G]�����}=E:�I>�R�j�9 6�����#�=��ͿHޤD��p���H='�J��������{f�D���H����I��H�.slt^��S�&Bs��Dy�NC 2)<�����Ʈ"�0۝�с�"�2j ����vq���ٖ�d����SO9e��"�P�vB*]���~	j��J��kz����gO�s����<�o��i|C��q�[����-���@ֿ`���1ksgp*T�=�,�OАҼ6����?���ȃ:��$\�P6���a�\�l���݂����qp�*�WY��Q|q�=B��3��eѲD*Vt�g�6u7�����0�(��9-n�fz�G)PI��vS0 �R�f6���9��K��A�-�@�a��c�Ό��t��g��.��z.���no~��W��A}6:����f\���D7�ٝ�\``�D��˪�	���ѝ���L��� ���}�$@����}"���䓚�c����㲏�^��9�$���)������B
  A@�GR����:7��Mp-���֦`���ƭ�Mr���(ͽ�=��1��uG�4O�:���f��%\���~f�A�s�:'�um����Asb�����Gd}��c����_��傿�X��u����/�O��W���!��f��&W�(>��x�B|�=�v{��\TFОF��R/L @����y��DsUg��K֖@ ��2��z�lo�i���/��ky�����z�=N��6^����6Neq>�?�̃�Ky��w�nu*e>S����Rfoi�!�1����?A��W�[�^�Ad�d�̏^�w�]=��΢�:`��:���gw��n�����\s��`��9S]o�Y�����.PCc��'|a� ���<Q�e8��W�>��n//��y�e�^*�(�AV�J�&Js�Ll!�i�� �Xdk�W�GT
�Dv62)	5`o�z^dn��I7���1Q���#�%�/lhqѷ�+X�k`Y�i�ڇ�� [7x�1�+�܅ݐwe��A�=�v=��k�	͐�q���Vvqy�t>W����K�b���Tv�á�Q����G֞�r�h�3��^��A4�]�o�<�Îk��5I�Eqja
�z�?�0ٓ%��A��:��e���B �l����ACq����;��?��]�W�U��rw�� v㆗d�e��]
'+��'(:Y�\�s4�.��AJT�T�k�x=K[T�:9T��A���O�IϮ^�7_g��zΉwq��ΠZ��ɽ�&ߜ��(ѠK�2�A���{g�G�-"���PX�!Sd:'T����F���Gh�}&X�t�-X���6�ٖ���v]N�t�SyH��5ĳ�BwCʓq���.P��P��R�l���	�䘪x?��)U�o(�1{��Q���dA֙g��J��K={��Fa����ԭ��,�Ћ���E��|���i���cH֕��k�������˻�Og&-Ș���5ʉ�+'��](4ŧF���h40˥u���u������'q�������Va�Y���[����C�Ɲ�ZA�h���ݩz��BV=+г�z6V8�y��M��������>|�d/^�u�sn����y����]�������i��X�0{��e@�A�+�beN.<@綈.7����j=z�(+ږTc�<:��1q�e�O�M��j���!���g�P�����V�$�xo� �nKN���ɛ8S��3^F�
�A7�5,��2F���ܹ,9X�9U��{�C�,W 1�5�UA�l٩��LL����2z-���2���h
+�} �x�%�־�1:�B1���2�A�j,U�_��۸Rp�5p\	�v_��A�j�9x �7�3���� ��?�P�����Uw`�!ZКPoq ���۞�����HQt����4TF�������Z� ��-Z^�M�`������D�4�A2�*��6�/�&�߸I8�ǃ��ຎ����H�it������ P�t��Ƽ�j��@3C&
u>�/��="��ٕ��}�Y�F�M�u�B�����. ��pKg�������h����484�}�ϱ�}��Q��%�̌ �j�:!?$�7��<�زq��<�a�>����φ:��Dg���E�3S�uP,����0�Є��t�.�#�3�ڃ�"�2�T7R��PAO��t6����]�%��+�c��ٳ*�j98 �p�]�.d�kz�������H�=�����Pr�ۻ��9$^/����g���� �*L9�
��k���v�|T�*�ss,��-��L� M4��5�P��y��;�̌,��B�����PbN��,�!^3[��
)���]�@�5�P�<�H'�l��JcX\\]����(�<������J�:�q%@ृ1,�^�l;�}n�<�h������OW�nQY@˃}���{j����)���r��8�(��;yv�J���׸������Pt����I��0�#)�r���S=�zg�O�Ĝ`��{k��;���4��<��s`O��nh.���-�Fq�Q����Q� #��U6�FC1��4��
.��R��=K�&�0~j�'�ǁ�1�f/������g����k��FQ�\w���her�
���Yx�a@����;����m��ȂuNd:�u�|��J;�#���5�lڥ&^�F��X֜��'[��Cd� F�����(�~�VA�� E��� � ��Roˋ���9�g�.��E��2:![?2g��,��}�����)Ti�(�M}}W8O�=k�*f�S<L����J{~�u�Nݨ�~�~�K�j�g�kr�܁p��_���R��z��ļ�e/���U|�Kw��BO�������v��o����C ��ͭ^/���u�������#S2w��j����x-O��G6��~�q����D�܏?��O���ngW�#��w�l�Όiv[^���FuR������䥯���h8�G��)6pD���7Lz@�Y;ￃ��L�=�t�F��f��7���7�y����F�{s�HN7
�R�J�Ϻ�č�$k�I�1��y�K�[G� �ad�κ��4.����0���y#������;��O�v" �e�&_�����w�XG���?��˃���m��|N���B}���~MCG�HB���z��jYI?*�t�� 4Q���fG��&��gH	pp������e��qj��z��2x��[pU9х�5�� �t��3�2F�����.��!�a�L���~/����!8��B����E8H���>w���&�Qf �;�#*�\�m`;#�-�d�9y�W��˫��z��޼yC��3
\����P���W��H ���������_�c��O{o�>�d?��#�������?ٿ��_}�P^�g��z����\�}�=2���:�吚����=[�k:�n��g8v=�˗/쫯����w���]D����rz%��<����೚{C��H�+ �p�?W����'���!`�CCY�����~f�-���b*%9��>���j�&<c��L�
���=�6��jG��Pa�`o��׍��� XӔ}�Lj-���)��l3��#8�m&�l�[H��ȔP����+�_P+���q���+�D1� ���z��9w��@@s�f�p�p~V�{˞�CE%K�	���L�<��x$"�Y�Z}����Q2c�{��(���Ȧ���!�=�A�s���
�Ni�XG�dZ���I-L������ګ����tT��������NaT$������ر����j{�-�]-�jN�&i�c�PfP	Q�$I�Z9�ۢ�E����JQW%���$�֔����Kl,�}���2Vo �L	;�Gΐ��Q�tV��AdS����H�4�iP�zj``H����[D�l�&�P`�r���Ԛ/'�8,q��N�C��;P�|/|�O�f��㯡kf��pBh-͖�,�h}�T?sc�Q9Y�cktI��/�u��'��#�3_]׏�-~y^[ ���a�׈��u;��	��s��Y�}�I�E�6�b%�cI��b��y��{�`3m�-�K)�3�}�����r �ҁ�%np�g%[��*>	H�4]���2�y9h� �q�Wr��h���D�g�1m�&�8�h}'s�>?��) _i ���=�lqr��#�`\Oλ�|�-�1�5ϾN^'���fN#͑ɵ�{P���_\����}�e��I�������?����7�����|�Y�}�}u��l3϶&o�����Kr�]��b��6�h��F��ڭ��G�e�ɲYc��da4 �+'6���;�!����(�w�L͇��e��h053��=yt��|8����g����ע�+�|� �����
�2;0�� /j��/���V�VN � �z��W01b�Aּ�M"x�[GgH�Q����K[�Km)� ���yq:1�orZ��TO�쁂����J�h �:,�G��F8=<Vkt}�7�f��dM�E<�T6�/�B��T�N=���#�z�����emκX{�a M�5be*�\�L��Բ]��qd&#�$���q�'�� �)�5�q��cF)o��[���-����gg���{]A��/�P� V�uX�����{
V0X�4'�?�y�~>_�ym���{�����������ꟶզ��b|�Q��z�����tN'��˻g3�=���Q,�;Q8���D����cR�hq�//٣�"�+`��_�¾�@k�/�Ï��O��޾�P�{� +lb8�)̿�Uο$]����O Y��iC��8�=U�g�x���,d�10��ٕ����2%��y�A|+�d1؅� L�P� �g��w�[�&�=�S�� �v2铢�V�v�|�'e�	A
�d��MGѬ!Æ����>8����-�j��΢#�F!
A��l)@����W߸���Ce�r����2�g�hSy���25L.��H%Ff
��6U�;�9N=c��g���UTe�?L˾�l��R��L�o�ɢ9:��:W|��3d����uBNgɱWh�-Q�U�˟b�@�#G=�A�ui?���Y�{Gڰ�Zcg���	��n�hT�mFyِ��]�EG#���y��zӇY��=gp4�=f>PF u�;������^�Fu!����ɥ,'��B�
��J�X��w�����"��t�m���㎟>R��_�F����f'�vֿ��{�&i	\ؽ���^��p��Z��Xx�j�
��|2M�	��/�&5����@'f���{�f9��b��-1O��q���������iM��&�b�(�R�IrB��? �f��&��B��"�:~�Ә���N����&�_�[��N�&�豆�ȭt�/���*��n�8�3PK �6�b�R8;:�`�������9��]�P_N��y-�&RZ�F`����4���@&
[�25�܂yZ�ܨd)�ZL�zp*����=4om�č������~��h�*���zn�tpG=�F3i��@�q����ǆ�k�:��G����L��ƀ�CE�>v����!����ڶ>)��2��MC�1#�]�^��$2/�une�N���KP��D�(>��5/q���m�C�L��"� p�+�b��F���r�O�e~:���3y�yg�#�g�<�ְ9�B��b7��P5l�j �C�bu>�9q����ȴ\�l$��ٳ~�tO��þ�����m�!�u�����E(�YL!i���I�f��f��:��I>���R�10�"V`mF9�s��J�ə-�k��%9��I�m�$.�W�O��1 @���l��=�f8�ޛB�F�x;  ��IDAT�ƚ��>$ZWϞً�/��rC�
�1hq Y?�}K�B/�kV?<�L l�����_��u��l����g;��x���~����w��/��o�~d�o^٫ׯ����;��+�yO`R��`�|O����W��m)�����:����Ƴ
�|����/Y���^�~g�2���3�4Q�@�S�q�:o�� ^�ha6�I�2+!��z�a��T^��D�*��+*���7� ���Ea�!1�s`�8j�P��ʣd/��2э� �����s{�ei-�_�b�h���Y�ew��Xd��p�O3WIA�� ?�skT�����8j��G�g�P�3~��5�8{�Vo�Т�ʐH)<g"� �j	�V�E-�����M^�<(Q���`����km��@�C*��W�r�r ��13�C2g_��ڸ�E�ۃ�q�	��.`'<+��L��T�)U^�C�0
=I ��(������Qv�܉l�`��\�:���RPS���=8ewу��ޥ��-Q�Pe��{=8ELq����Lw6Tr!>=:^�h�E�Ȉ��Z��͎�}S~�|_Ս�Յ>U��1{m��u�i�<�����]ȧ��C��gEc�g�rxƨ�É���l�����&T�5�E����Dq��Y�Úp�i%6%w�cqk�n��`	�����Y�=�F������sL�9͋0��yc6[S;9��	D��dMv]���n���@���E4c�'�� S�M}l�LƊ1�h0��׾��V�QR�9mE��S�L6k!E���EI:_�ThHc@���w��rU����H�	q���4��fE*BY�2���i��*ct�דKB�T�>����.M>\���
G�����MKo%a 7����KD�%���{s�h��[�� �V������嫴{X��1�6�Si�|߼�!D�ߘĜ�ᜇ��`��1kFVk�)��K�Pyl�w�!�3�h"�.�#�-���8� �C�D	�c6$�~L(^�j���/.����{�칽x~�^8���d?��w?}o���Zޡ��V.��r~%��j�N�`lNY��f/�MĆ¿�k�I>�Yu�\-���s�A�x*X�H�gg� h{��U��Y��a4s���l�f����5P�e��iNm혬�
6���w�^J}���rx^�m(G?-�����Y{�k+�B��o�b������W���(r��B���y�Q,s@Gh4��ʲn�(	�䵟ܝ<�+2��{�]��RV���t�\��:�*8���R�<�D�a�Z8HI�����أZ���q��-��СBvu v�����qe���cfvk(��`��[K�̀
)@��`�a�KwFV'��&��Ȁ�W�I�����tV�5�IĘp ��C�jB�5y�ʃmr@���.�0%f>���6k%���}��(��GQx4�;ڊ���:�s[�	�'��Ǖ���������HҖ��N*K�}r�k�ݟ���l���d��pi�./Y����K��o�-��~Q��W��&׈���͵}����V`�����O�?������#���1���;_A�a&H؀:u��>����]��w���6��	�T��廧p���-��4�i������׶�(juuLvP�p�|�Ӹyf�V�nށr[�cbF
�v}��K��	�N��&v�ۮ� J�Wt!�\������Z1�Z*�-!����]���;<�a��L+ob<{��ʥ�3�禂�l���=�0�V�u-������7vq���E�$�q�g��"c�?\��ӲC�f�TX��H�LԹb4�.C���h��/l�r��J�f"�h��0Mw�w&�x�4��[!!(:*�]Q�����Gfޝ\�Cc�0H��t&�J�>�� �)��Am�i�jb�V}��{��;ǲ$pr'�����X��{B橎�|+_���L�������Ǿ�s��q)9��Y���}x�~���NC���A-�@O�[;�O���:���ol�I�oS< �x$j�����ED^ݲ;-���IB�Rmz�E�{(��R��ӞQ�w﫱x���s�ЃN��{&�:A�A�'D3�J_شg�Y0e^�]⍫0���;l���F4:I�ז�
����j�,���ɉ�gx��NT�҃q��8�K��Z8��9(B2�z[�A8(�~IYo a�����T���^~�;d Yo��e���� �ᘽn����(�qݤ?�Q���HW�Q��ۓ�ԃG�mx�4u`��!8n�q8/0r�����$SVZ�S>��~"�E*N��dr�b�K�I} z��������|��l����x}��u9��ce��Ws>��xo\����מ����:���}��k���ϕ���p�����P���^Ohp��9"p��;�"Ә�q��4,�:"f1��v%Z@D�es���%�ë1�`�Z5��G�bwow�7��
l��f���ǯ�3���"���Y"s:�� s
Fv�8�HPq#]?�o�����$��)}Y�#{d]Qv�;���@�ԁ��#N��D	����s�?�ze�)�t���͕��Sv*��j�y��D�|�QЯ*t��|0u:'���<�z1����Ig^d'�0W��qh�B�����y`����Y��+���+Ks�T�l]r�i�Z��4�|K>Fa�$5`�i�<�q6eLE��nLc�%m����I|A
�\�6�5��)�x��3nN.h��w��#�G�}��D0�&�y<��͎�����N㠺#�:��%}���;��ϔFQR(y+ڔ�N�2���(�L��Uʔq@�}��%ʷl ,	h���s�5�F�ww7��?��>��C�k?ػw���~"��}�.�ի��F�T�Î��U�AP�c_�z~Ԇ}��Wv�ݍ���O��_��zxQeqo!�U ���ĵ@f�m\���#����M�ewp,����D�7�l^�ij�y�8��r\�j�`��F>��s���<ˤ_�ƥ^C�W3U)QK5�A��!����U�V*���v�� 8���Y������vql��+�|W��ݞ��7(劣m+ ��x��=��?gO�5�̠1�Ǆ0��Oע�VP
�sy	��g���U��8kfQʤ�v̡���������g����M�)4�ۗ����x�+��3ź��<�~�
]�)��H�����no�I'�"�`�vIa�:i9'خ�Ɖ�*x���/�Y�պգ�~��T�k9]]<����4|�Y�`�V�˿�*w�٬lq&S8.�}��u��@\��<o����n`��n�H1�e� P�5vYǚ
�Y���G�z�cK,W��d?�����F����hǺRl�M�Xd��t՜��{����զ���ܸm��RZ�/$~�&������	�+
�U����g�����@_�x!��d.�x  ��N6�7_����LR�9���7S���s��������Q���R+�7� �N���O�����z�Hj#�aٲ ��q�}��o�����`ij��&(��z1
x�"�*w,
��uMU�	t��)�,mV4	�\.��pWR"(-r�H�RK4B-#����K�*���l�{�5�N�)z/z����*�z��6�Y�j8��)
NF<{���Yo�W��-�P(|>�qN��ï��[K�?:�1}�bUqd���!�*��~pM����#_՝�����M'�1�x�?�ၓ���U�k�0o���ߢ_θ�Q+w�{��l��♦�6�t}��y�-�ҥtb����+���'T1�^�Σ�i�e����ɓ[r���
���on�yh�j� .�կ �� ӷO�I��
��Z�|������i/>�����K$�J�#Q ~�&�d��U��l��N]S��AM
�&zO؏ x��P���ws�"�>�f�e��E륽=�@'"(��1�G���Ή�xAv�0D�n�r�p떔�sN��S��{���:�in���sH�" vi��u�a2P��t�Q_�/K���A�Eԫ�#H�q��U6�8̘x;�`�"���֋���Qk{��ɹ����"Y���{��IimR�
�j팽�F��T�mQ�5i���@/j�*�51#�Eq�+����r3����F�o�3�����#v&����>_����wvt���1�-�92x|�2Ա��֭8v�Go^�5���C���nk>����U�u/�٠Q��6b�A�� G?|���Ѯ���j�`����#�&2h�$��Z���v��P�E���x>?�/��¾x�{�����r8 ��}<�=��8��oo��\��Tv�RI�<�:ms����{Sm6�
�bf�(厘��.�]�r�o 'Կ����١��?�?����"��^��o���~m_T�{eH4��s��]d�������w>��?����������ط�|ao^�g� ���U������ßS�Z�\��7_�����_��S��LUN�j��V ���@��%�_<#�<`�����w���
�޿���'9�H6�;�\��#%�]��n�E���dO�F?T�����m�1'Tk	��t�
d�b��}�m �P1d��R���{�nj��;�'	S�OuOT�h���F˂A`���u�f����v��ye%���>�2 (�?��
�p�H� {����}o�� ��_�Qt��$�&���T4�?U�]� �͛�����&y-�c�����jJ��N��e�B�첻qL��0�(lKG:���3�?�냾�~�����?�u�z���	4����w���?���N�~�(�Z���Ms������E�B���������7ؒ�JA�\���`��v�:�"R���'���>���ҝ�a���R\�6,E��<�u��	�B���c�g�l�a�!�B��q�D����s�$#�;�� ��j�
d�!G�Ɔ����R�ca��(6	��5#N�1U�Ns>�|w�q�h[�#݆Ԁ#Dҟ�]��>r���o����w"*��ei��=	����8#"�'uH&�ݚ�>F2���E��wS��s{�e�҃�>�@��T��Z�u|����v��إ@�v�H���GF�����m������ulC�CrP��ȋ���"� 탊P��/_V������l ��q�7𮲤�U��MA��
�#���(�.�=��̠���A�4�p+�������h&�M7s5x�"�6�<�.��!��{6�r�2T�MҚJ�Wekχ�;��|�z��`��AQ��^�3h!�����328sY-렵=Xlv
0���<p��&����YIawu�{��"�,�Y ��H��${F���P���G�A+ ��Hp�e�OHR����4��)������x{�.I��J�"T��Ҫ��=�����!w�E��J:�ݞ��ܣ��<��oc&:+##����`��Ņ�!��cGNC/,��s
s��*AI�����;�bQ���/5��pv����!(V��l�{ҍJ��=K�f1��5;�-��dR^?��	k��S`e��}7�1j!h�G�w UP���6*�@/04�fK��N ֌�Z]��.�����ѡ�úJ�[A�m��
y���U��OZ��ݭ\�}���@&�}�l-T��3F�YOǣ*r]��(���	(���j!��ZW���N�6[���6Z&pp?_���:9�[_�U^s�h��g�F��ExJ�ڡ�M�^%���㕬6	p���@2A��q%=�L�EK�3��.��J�z�`8�K�� �n(�AY����J �@�{�D^�x"g'�;�A[�l�fЌ�(�~�8��Gr������}������������#�MN��GO���7���Ky��B����4(�K�C��w����ʻ�ٸ�Ϟ��7o��W/���yr�1X?�����Z~~{�|�"�ir�O���7��7��gS�ܨMn7�_<, �%M�����ϣ�hجbz�R.��\�� 
��&	�a΃|����Kf� k����B�}D��E���}�Z
�:��(�[U����c. H������SPo�s�1����%�$G��PUڼ�R�i�AD����� q��~��\�\�ej�t�1�t�s�9>?֠D�H�|6 ��VT:���:<>b�p���|�@�|�f�oo�.��I�=:�'O�Yg���X$���j�=�<,j7�w�&'�-�����Ê0��:��1�>t�7,���������,���^~��or�. ��Ǉ��C9K�q���#A��/�1�I���X\Ͻ0g�6�R��+�{l��f9:�wE����Z	�mV��͇9�9�� ����;�Ne�A�-\�Q��\1�F١ �&٭��j�KSSBq�#Amz6���,�@lɻE�'p8U͉ �������F�Gu���7ٚ"�E2�Fǧ4�'�4��L2�����u-w�&�(�J�q*G��I6�du��o�bgY��݄c�ؘg�4kf���X���)��W��N<�l�hxǇxb J|>�W���A��Al���y�H�7��d��5#������~\�������LW2�9�<��ٝ��T�j�p� a��`(waC@j2V�	t����d�$�P�I�:���R�`�V2��Cr70�0��%Uj�8;��#��9�����a{Y���*jmH�B�ʕ���V4Ny_�cGN�W3�e�[G�E���c4���I캃�-������y��|E]T���G�5���9z��wZ����k���O;{*T��������K��t���V��遝����`����������h�xR0Q�,���N}�Vp!����;�7j��JWQ1!"ٮ�x��4��i�im�5��&�f_��IY
2+�Y�v(�ɹ��!NՉE�|�d���u��_��6�V��S:��9`x�ue$�����d�}��@�� OeZ��[�f�[)6�WJۋa�L�hl�� ���}���妹�mu_�  �: ��f����dCg�)�A�n�^��l�I7����x<��E�;Z.�>��A:��O���cfL�y�}�-(���jAg�Kγ�/�o�Y����[�,��a�@�R���u�=�T���*ݟM��A�B�k��1c,��[��R��	�����cI�6����1!�:9��`n���HV��C�T�~��V�r��ZɄc[GO��":S;^����ũ����F��?���}!g'�A8}�0fpڧ��d��`%�;U5y��J�/�ɋ���U�9;�H��Ir���L����.�<|���'��F	D�'��&x�z��y��4��J�E/���ۻSy�x"�g�\~�H��I�@�ky��<��iވh�z����}H��^��ɑ �֪�Κ��\���"��缧�Z�W���n�����?<0��J=���if*�J�s�T!,dvـ�ь5��F�XO����$,dސX��ł 2��쁲�u����hd,3mb��G��G�� �:�O��Ҹ܉'<�<u�&=0��Mf�9��!H�w{�-��h!+��� ���� y��D����f��a��j� �:Ix�� ��vG���s+�r��'�^iPtc���m��T�	%2	��Wi�:�z��Ŀ��?��_>�I�@c����!�zΆy��i�f�q��cI#�]��˴������`)�2� Yav��f�����c9��kN���kB�7X{�u
�}o��*��9��bΒל�yݙR��,
�v�'
!�8� ;,V�w��57�zz����h`�>����Ui��d�{7l��]IMl�ؖ7A�5Y/���q<!���u���5��icւQ�J��h�E׏a�[q}rl 4Qx��f+(7���RGJmI���=�ls��^��/ۻ���#� ��^C�+��ԃ����L�Y2?�������y��;<���z�;���S��.N���_.cg�V��
�,�cYPfy�l��w�"r�໶b��f}���TVk�3�M4����Yc��{�ʤt��m�7���gtl��A��V�|~�V�i���(�u��k�����֙)����Ll���b�`w����������j�<)�ȇvz��I�r���S�^Q�@������6���q-VGf7�j\�{o�$Z�4;�����,����y6�TA�`�B�!覯Yw��p9�Y�-;�w�3I.QM��22~m�h�>��8֤)��l��X����]F7�xf�^�\h�sG%,��#m���ֶC0ᐨ�{�@�t?���8V�Υ�U�iUL��1�Ϣ�qu��z5��6Q�:��d�4�4��*h�k<�����l�t>h�G���Hq�#4dWh E�R�T`D+���q���wZcQP�F㒢a�ֱ�z�U)I�u��&�-a9O"����|i�M�`����� �f1
��:������~ivGAyk�Q�@�Z�i�'��L�.���q�@�zf�cD�k�$2��a/��/Қ � � �S�*�b�t?f)ʝҏ�M��6 U��f_m�ڵ�$���g��$�_j@U�Hh�e��U�i�����C�e#5AB/d!55\O�8��2�`�r����4�^={"��?/���N���YQ����7�gc=�J������*|�0^&�{����޼"p����1KskZ�p�
S��L�	4�z�H6����Gǧ�$kT���R��[9����q����Nӱ�rtr.g�i|*�}�j�T�T��[M�4�i�m����]k�
�@�4~x�͓�N.��]a���}�'���	38��f�F���ڣ��>ye�ǂ�u���������0c�duJOU �>޿
TA���N�F$�q����X�X#'�y���k�`���� �E|'2ph
M���eN���D&Y*�T����@���AAuJ�z1��fп.�i��t,�g�����"��y�9��o��'��rO�ҕ������]���Abڑ ���M���g�&��9H�4$��@��r-�K"q4%��� |TD�g3���V(�bp�Rfs],��y�PFO{O�ݽn'��������H~n�<t��c`(��L8Ń��d�m�zy�_�Qx6\eA12Xi퐽�s�'^#7=�/85��B���Ǻq"z��]���[0����71���b�Ţ�nZ���&�Xn�P��b6�T'�^�[���y�wg� ��"&$ 9+���e�b3t�0��=�J.�hR���\(kԭL�~���H{t�Nǧ0�}�':�'�:�ʛ���D��]�y�;�[X˓=�Ci���j�I�����020�{_̾� X�O�ә�8|��8�ƾ�(�}�o�g�w��?�2��
��sC�,I'Br�N�7�RD�/��i��8��&I�HNǶb݆�_Sm�j�'f���0٫#:p.��l:���ym���N�L�'V�Մ��`��i7=�F���Z�jG���*�&1�4+��4q��v�M�{�9O]ϋt_D���I��u�ՖB�,h-�Қ��;���Y�)�]�8g��t���?��� !��ƥ2ѝB.�[Rx�m�N��yi�ZՁR];_�����s�Fm��T�E�N��
����4!�#ع��<�B��y��%*r�)���~�7*�Q��)�����.D�N��:}_�кf�t���S���YF�EP�,��A�}0%J�BV�	QI4lc"�c4�Mω����h�G�:8%%�� -����c���C/�Z�� X��|؊��v�ūX��#j;�J�.�"��UkH�Y��,E����mN�`�m�9x�fۨ��:�%�j��i�9���H�Gw��3F;���e�^��=(_�ou���$�v�P�����vJ�ʑ6�e����>Ъs�cf ��1�� .U�~Kg�`lF��)NP��J���w�X�ƪ���њ0��I������X �O�XS^;�j���(D8\,ٵr�"300�2��P*"�X��)�{��:��+?��z��ĩ�x�T�=}$�Ώ�xN84����*",+�"�٧Z��,��5��g�3���ʂn��	�e��<~tA�k}��ʓ���=�7�u !%����� 3Z[%�@7�Yh=.�5vpU�x���6�~����F���w�y pܙh�niJ���5�4���B�Vz_��WFR���"d� �eL�X\�֧�t��̔�_�<�x9;������Sw�ܫLD��� 蛎N�[N��V{�E���0V�4a��Y�����$� +X�`�Ccaf�F����5a[�p0sL0Gj�/e��z��r�6�d�s�J4$�;A������s���g��¢jX,���Oc�A%��d"���7���^�>y�&���	����#��|��?@�	�~��Q�N��cs�8?#Hh۾A&�;�����ȅ�~�:��3J�ć�8�t��G��� �����w�5;q��bԳ Y!��^f�CS�]����Q�E�k��Af���ud��n��M��8N�d;:8����a��x4K��"�=`�,(��d�,Ԩ 5R�t��f�&����e4ĠCV�Yоe%��*:AIM��;���A���'�3Ψns�����b4�U��tm	`�M��J)��c�UI+d���^�z�׆�?3��1�������������r0n�'���% �����/�A�to�y2_�6p<�����_C��a���� ��|��K*P�y0��5O*�w�|�=�\���R�b��(�D�-�!�ƛ����Fl�(���7b^]8!y��2bi緋�)ZV�(���;��+́��xyCաr"����*���0Pl�ҿ��Qmp���[l)�e��k9fĻ*-�kĝm�����iۧ��k���,��S����Fsm
;�8Hr��ET��}@���@�V8�U�;�	��x�Jq�0���
����!f���Y̱N�����G位�Ӧ�Z��n%�G,�`�mQ�U��P���2J�K��i���X!�h@��|�sэ���:�M��,���Jϖ�2�l�FSXtjށ� -A�_�����U����(��4��wG��bvĹzR��fy�7�:�ʝO>�;Jk��6X�>��Q�G���a�h�Y�і�l-h��*�,d� ��vF����
�g��a4��X�K�
�"i����gy��<{t���'TRђ�%씶�[�M�"��@����%ol�|�����(�]�T>�<�+Y-TLa��&c:3�޵J�kFn��Z�-;0��a 8WWr���|��$�9*����ڍ]��qַ�u8c[�%E�Q�lup�j�F5��ҷ��y�8�#k
�F�F��yK3�D�M��:�0ә��5f����V1�����Wlѩ���fF\Ч��}���L�&�m�4@�b������xH+{�����4��,1�[k�����k���A�S5PTF�N�9 lPjL-��D	�h��!.��O� JgsH�ϻm�s<<J~�lL���Ϳ�����#���WZ�m��}���膁�L�_5�b!`�Й�i~ao�~�s���C<~Ӱē�Td��= �!�ջ+OӤ���yM�'�B��B�s�ܷ?#�T:�j��,3��ň�͢��7(x�|�X~������K���Ed���O���r� ۴�/?]���� P8y�"���Tee�7�n��y��T:��2S�ڙ,mt�҃��O�&��qL�d�O�#�>�x���Rq�B�	9ͬ�O�VkB��b���S3XmY�h9]����U��,XL��pv g'�r
	��F���=��i���R3�8���,�eg#n��E�0NF�T�1��րQ0��z�P�7�e��Ԝ��Կ�öL�����$��~�\�f�::ĭכ%�Vq�x&!��N��m0�Z�gR���#J�spX��n����,��̑J��m��8s�E�Y�7p31G�_C��>Z^��ks��ײ��Eo8���ʟ��g���X�2���q �km`��bP�m�����7k�t䝁������hT��hC�H� �Y-��I1bA�s��sp�L�9��@��ze�0�AV�����~�:��UeXlr	�C�Sˡ�R�ket&5���/Ϳm#d�#RB(i�"�����h� +�Ҿ��,4����p��#�z��;;����#D��aٹ��
 \������5���e�}�3Y^��s�&#�)�"?��$�r�K�-�?ݶ���M�4���v�����C9=��۵A|k�P������m�X_1�dc.���u@��V�������E�;J�Pw����=#ś #�_f�������&�(P��`��q�[��[4v�As�h��G�NJ�Ľ�c5G �	dA�%e��V����o��5���!���1�:�ub�6�����s8x�6����9��"��c���{��
1�A/���}i;o�����23�8i-
�I�lTHA�c�!���8j��g,Q�u�I./�>{4��Yegq�-%����0�?���{sQ�l�>��dei�5*b��҂
� ��JN'�`�Œ�N�q�����1KP�uJA��Jk����C%�c3{������&G��� Z��&�B��z�#f�
���]#2P�V�@���;�ڈyo�K���6("v�;
͚�ue���uQP�u�_;���}x0���W��"�x*�����Z�[�=���3pP5Z�^i��cv��Sm��먡�	��X�ʱ9;"U�}>ߑ��yZ,X\�sMS �2LN
ƪ`��� t�5*#�H`�gm�I 2��Q�?��t��|N1��F���a�j��B� ���Y��~Ν���*����&�)`����l��X:�S!�N�>��^Z�@�y����	��d�!kĨ��,|��a%��V�$�i�2�{���c����6�  ��ļ��Q�@��!h��㖽A�L�eR�\�;U�Fz6�B�\�N[�����h�n�
&�O(C��J����Gm�0$�bϦl�}�_�p��^����Y_�g6l��o�j}M
�_��W�/q���r~vl�n�5�7P �Ι+�e8����=�E)�=�������#�2Fw�����/_�n����$����Fs��,W�Z�F��1������Mض�EѠ61�����'�{�*j�53a�-d.�lp;mr�F�X�>[S]���jݐ.�^7Tc!m��Z��!r,lc�ǐ^�`�I����ǀ���k��+ѢPJ����u��"����dF?�R���Y|5�n[>�>�5Dy���s�A�ON{�a��_�wZ�0�p��2����S��_Cq��_�W~ѯ��jQ����}��nޜY���K�R���V��t���SU���Bθ�1|u��B��ju$�ʟu�evwk-�[��u�
��R�p~:nk�KU��Z(Ͷ��S���ri�Y����4u�	��|I��B��u��+����}�I��O��wF��~}~3�Vb_�Dj�����S���g���E�!)�s�i��?K�ӵ��5EB�`�)����$p2���K+�./?Ύ4 -��p�`_"�;A�	7��<�ˍ����!��C�(R��� ��[Z(�j�V:ucCg����G@�i֊�Ҋ��e�l��7�D����5 �{C M��̕F��U�:�Y�
��2_є�(��w[#]o��^�r��H7�D�%�5�ҹ��� ��rwG�bkM^�@���q U]�y|9����������DF�Ql	-a��6��������^"c$�Z׾��l���D{<i�F��L��A���C��Ĳ��A�I�MkN�%#p2������9 T�`��ViǨQAV	Y����9�n㎰�Lwf��4ۙ5�r���Z#��8*���yq�X�A�Q]86�*�JL�~Gz|���6$�і���|�UhDF��@�B3ˠڍ������qd�Q#��j�ܢRJ3��,��j�ڒ��FWwU�۶A�J�U��ݐ��X�k:����^��o�&����=�KϞ=���f6n�
J~�z����o�ؔ�:���*��N��(�����y���l
D9p�V)� >��q���zT� �]:���%�����S�L��C�v����Ը?'�{)wk�	�}Z37��JCH[D�Ĕ����[����.oT������錉���c
Qp��"݋�f�X��	���� ��C99:���c�5���(@Z뺡2�Yr������O���tl�yT�I�ݪT�ku~3g&�	���>g��O�36d�\����g6��2�G�A��b#'��2���*��U��*���/�(\� �nZ�x��2��m�����f �P_��(���(��P�G>MB�S� [;FtB;���v�cj��4�[#�8},�}�6�u,8�5�J��ؠm�^��Iw;<d� ���0�Ga T剹�I�]��j�W�wDӛ���֢$*ҁ6̴��1�Z���pv���L�RԜ�-�yT�cX��P8Ţ�Fi�W�ܤ�I�57%t!_* J�h���;.Z;��JJ������41�͂�#2ZPX��~l�i��B�CUŊ�I������`gi�P=M�XIZKLCo)h�j�&9R�0�-��MK�_^X��zU�,�Q�+Y[)bdFj�X&��e��A3_�����A�fyx���g-���g\Hَi�ѻ"�a<�,�e%Bg��-�ýѨ뻨�!|��>���h����r�6�#m�=����!��0H�.��'�ڍ��O���F��5Os�ȏ#6~���s,���}����Z40����Y�%d�י"6^lB��РFF��l��x+Zͦ$Gb��z�2.�i�n�Zn`i����P��`۔�0��V��>���i��c9N��і|�6<{��Y���ܺf2Pl5���'X-��M�[@hFҺ�,;�Q��� >�O���P���n6V���E��)V&fS��F�ץv�k�@C�:���2������aT:���]��
�`�Y.q���y]8;�7`A�����r�F����<�J���5�,�v�S�8<�)�E���4�[Y�������I�bk �Z��~"ܾ����z�p�iʆ�▋_��.��3h֛�2�n���K|2s�Q�������	6�mM^� 3�"`#hK�w��#_��R1��n����<SĨ���
:�ɦ�
֩s��fCI	�H7n3@����-���VZ�UjE�#h�6��׷M���cx�3PZW�A�2(�&gq�� ۆ��Rڟ� i��$d0��[d�9���8%�?��xʄW�%쬙Y ��̯Ws������k�-Q����LN"��SԎ_$��4��N�(9l8od1?^���\��K�# GdA��5	U�3�P�vY����Eor��Ncb ���`�``Tz&VCG?�aM����~к0��?������XB zT㘈��:(c4��i`����&�#�$Grv����9ە��Kof2_) E���7�����5ޑ��]�Ӵ.৤c%_b�^+�06	TBX7���4��pl�=�|�W:'Rlӽ�p{+���<y~&��Cy�h&��6*����Ϸk����L��u�SL�0��iF''����������n��rzv.߾�	 N���*�S��[m��I��|�����LQ6 �h��'����g���$�;��:���E��k���^���lܗ1У�3&pm�!�x}uEq��W�	0-hN�N(���'�:z4�@��2]�?��Ol{�;M��1|p����4��y��q:~�ϥ�� �X�Z淟����&�߿�݀�ۛ�0��� �BiA|����P�Df�/a'Qό�
����e�6�gVk�ʤ\w�>Z���:���b�L`l��e�e��/�	Z,�i����)Nrt���	`M�ؚ��6_5�dBE�~~���,�$�{����w,�*|���������^���	�NҞ��4 t�}�9��-����Ϧd�,z���� &k�E��R�V	}BY�a^�<]eK�A�=Z�_��4(~��9S��l�� ���	���N4�
0rjt�@�wڟ~�g�_�]����� @������H��9���׽�D�Ɍ����|�v�qd��kC�&�����2ݏ-3W����x�;��#ǈ�B���耊8(�%�*�	�6�����ݐjS\�v:=N�3����	#�0�E1:kp:Z�n!bB�G�*_'	WPJ+�I�F�b\6>���qK%��N��K�"�(8Zl9Ʌ�t���7�5B�E�h��^[��c�Wv7Z>��C��^�;�{����2�Wy>2D����T���>Kj/ۿ-�*��}���w����p���]_do��_k9L3u�/�b�~����Ȁ	&��yf���72"���2�Zcg��J%T��@�0Q�����$@p��󅜢� U�&4��A��f[m|��31�2��$N�t1���J2�S,,�v�0��<L%/�.�͊���1��5�eW��6���Ձ��bfX$v�vY�Z/?���}�JQ���Jm3�n�a8��Q=q�>g��6��mB����� ��琊Y�L�۩�,�k\}먶ə�mYc���N{9Ū� �T���E����gn3PjSi6�d��d�j�A���Ӥ�F��V�
p���6އ}r�m���\nd�LRY�4tڃEkִy
�+�U�v���iJ�a谴&�b8�F<xH�m3��T��hw����\��'L�G=UF�+�ucHkX|�R�&f��\�s��'v���*�ت�U:�c}�^M�
�t&8��n �:��.�~�&b&,�Ϟ'���Ky�|��G2;��o�U��+։�	�X31�eԺ�~]#���
vi���9�z;���d���E��Q�γ#
P^���t޻�Ke���ݖW4��1����Nhܷփ[]�%.\�����pJQa�4�!�\+��=-�\��j� 8j�P�����QJnI~�@#M�t��`���[���Y���k��O?������)%ͧS��ӟ.?˟�����x�~/X���(��7PZN ���u'�	�ӽ�% q!�	8��哜�$�s+�6y��g Mw����׎q��"�>O�#�+ d��$���s?���oTM�":O�����x�'�g����VlH������k�I�lXG�d5i-~�����Y޿{� �B4c<�x"؀L$�!Q��dv4�q�#$:L(ǃ���ŝ\}zϹ��˩��c:���i��H�][;R��>�3��C7W�˲��������c�Z����T��!k��֚D�x�}@V�6�c�LPi^�|�$HRz��#e9��Y���z�@�r�`��TWpj�	ܦ18H�i��Xggg�(�9��4�����g�Wc'�a�P�A��/�7u����m��[��)c����ɕa�n\���]���f��E�w��)�R1p�Dr�M��@�L�&�X��0<4PҶK-�ꤰ@P��_����/| �=�>�o���ڷ�|������@��%8���T-�&u��VVC�@4~ EOȷC�]�v�g7z���i/sk�@����
j����]�ȠacC���J�L!��^%g ��$}g�4;6`��rSi���V���(�< H+��-��Ky�Բ�R�8�:�FR�Ԣ�J�	lr�5'�F�a%z#�k�V�bE��@Kͨ�Cfu$�T̝9�C��� ��>�#�)������{z���r����p��d�~���!�����������K������tRWZ�x�\玑�f\���n�ܘ�0ص�1��Y���p��E������^a��/9���ƾ6*�2߽��A���[�w��.o��S�3xQic�˼�l_�Z�`��=Ź2��/�f�9խ��pP�uW�ch�$��D8�8�	Q�D�>q��\�4C�:XsҹNJ틣�6�-��Wu�A�+�X�P�f���dT��L���1d����)7T�pcY�&�]@�i,�y2�h��
����;�l�X��H���6`��wgT����ȢTg`��$��^RJsގ����8'U�v#�0�e�md�)АP�H��"�\m:�N�]�&;y& f#edu+J?�p�ٝN\��J�{���YZ�e6�2�ZT�Z,<<���Vo�����o<����m׭{�R�.M����VC�=��	�Q�
K�2��)�{*��a��*�rk'S����ް���8��>~����tt�>��$�Ը˫O�e!��s���z��-A�:�x+ @�6t���Yd��m���w�A�(8�8Wԉ"{�^j��'z�^?�k>�w��6T��0�}����{b�N#��]'B�Y�ʬ�׏�Mbt��|�\�n�NL9��r,6*m4��B�>�MŐ��?o����A>|�$��������"j�'��_�_��Or{��z"�{�)C��7�h��|>�.���A~���ȉ*�L�z��u.WkZЌ3���(Kڟ!�9c��������U�=�	Jd{�0�1=����;���t�w������6�Ez��-P���v���Ž|��b�a�&|��g�( ����dG����;b�'T��g	 �M(��m�緤�~�J�jca��k[������马ނ��@��G]�L8]o�5যj���w�h4�F.���镶K������ky����B���D�f��Auަ��$�Sk�H᎚(�V�/P{���UjrG���|�l���Od�z,�d����t�� �q��"n=��?g?:��r�;:E%{b���㿛䀣`nC.�~�V�	��t���QD���v��p�tt�lt�M�Qw�Y,i�0"&�m��0D3���r0��v\�?�9���{���1 �=�2�;�����6��`nI���ne,��z ���ez+�[#Z�ϛuj?�R�^@;�j�i�.��ɐ��;�0c]"�3K�C#�@2P�V��B����8�@���G�����8
`Hǫ��U<��b�v�\em��2ʛ8p�����C�����EXFue-H��;5�/�̻��:A�`� @t;Q1��fd��_�@jS�#��_!o��Q����/j�b�_g���ݠn2�2��~��F����]C�;�! ���8��_<2�⩅����z�kBr��h�4;����x1�^��/G�ՙeƤ�z���\�]�Թ~ E䊑���{1:J��j���Iz���_�"�z&��=rs�!r���w
�	�hٝ��`�Z�����@�^(��U D�����#h{�F������g����:*l�|��ǌ1@� îN�ۨ�B���hBux0!��l�xZ�� Y,���"��#�Ƣ�q����ϲ�pD��^kbǇ��<��pN��B^�b6�t�D�M|c�&���Z,XK�|��X��S%?PI��a�?��0
�ם�Qu�LX�V-�G�ds㴢X r�����x.	�;����a��a� GLv��zێ"	�UeVNk
mr��:�_���.��(BbuY��yt�T�C�"�����`�``���V�:�y禇�z	��ֲ�>k_*o?͹��ɖd��D�M����f{�2e�*g�X�y��^����vN�(P� �"ἡv5h�
�"�r�W �h̊�Æ+|�A�1���:�]�$f�*.l)R)�7@s���1w+�Տj0�w|WŚ��	�Du^݆Z�Bg�
�[�8������:��d��~��d���F�2~B�׶5*?�3�����)]=U3Y��TF�iP ��[*���}�)���ׂΫ���v%�1�f��SR�j���E�������U�?-�i�->��**��Q���&���.}�ͱ����G��`\T
'�˼I��H�h��_ɧ�[�OB��N�����Ǻ���1S_U����T\i)��
TZ)2��(��XD�X���6bIq�ר�L6�!�5I6*�Pʄ����=Vn�~��1`Ϸ�3Ɍ�vk}� (�·=o�\����i�cg����ю�S�=��L8��7X����D� "��p`�̬���e1�����7��f��k5 �k {��cߠ�Zg�Ƞ���-mc��b������[�Z�V�3��Ԗ���6;y��e�7��u��t��3HsSE(J6,�k4+��S�<�dwlrW�P�p4*��M��hu�ĺ-X�W��δ$'O+��`՝5^��
�z���>��]�3k�m�ip�'k�M��}p���4����}pI�A�m0:���"MpM�@�*���y��J���F���
Y��q��'�"�x�P���X��3Y�h4w���v����;� ]0m��N�[7U	c����Ԙ#s�s�.
�g�zJ�6�o������/XĊ�A&�g��z�*a��2�!B��G�zB��'�2jEۮi�)�g�o(�E��P�tK�R/
YX���s���@�׎ͻ/������U�����j	f��?�`�%ټd���H��~:e���>���/�U>���L�Dx2 �!-��4F�)��F�Foa�Bz��H�~W�;��B���\#{�!8�x?8�?����������e�C���P$y�QN�^��(X�]ok�Y���l��l�������@�[���\����ޜ`g��y9�B:ȯ�R����t�ڗnbi�����ŗ��'�5(<G��ON"դm�I���y��,=����	ս b�h�V���� RY�(��'��L�p��J��Z���ц
Q F Ǔ�cn�O?��o^��x<g,�rÇ0SeE��H*�D��FY�ͧ�e~�^HKЁ���FVh�ADA�l����f�9@w\�dbsOߍ@U��� (]�*��C:�{����|��M��Kr�Y��J�lakү"U�Ƥ>R�-h5֗]��4C�J��Xs5t���Z�����Ev�*���"M��p�x�Aoqt~�p5d\86N��b�����6j;;���536��8ŮQǞ�m�_�uZ�ʩ�1~��T��{rAg\���Y��V.S�Ҙ��i�,.W%��I�v�$
Pb F���Z;٫����Ԅc8�p�1� ym�=%�{�h`9�^�*w����]WZ&O�N��uP�KI@�l�$
���5��i�K+)xb`����JH!m����:Q�����!���x�ǁ]G53]�x���� ��~���0C��]c�N�h�6PJ>�6�b�ht�yޘR��%�.�ad�!ʶ�Z���"{����y��������F��N�u�cH��9CѠ߽31�uc��0LJ_�r`�E�gb˃�7�dQ��'�>ٿ5o��ժH�� =lQ].����@	��R���Сe���_�)���.(t��Њ*�U쓦��c�s�p�j֩(�i��X�G��p�j�=��c�[�΍��z�{d��]��T��/hU��m���Z0[�"Ы-Vu=��	p�o�5t������:�7ݻ�$�S��(���]G�ZW4b����Ǌb��>}ͥY�t;��N�W�"��pQa0T��eA�� �cq��bU��	0�	QIvv��jejjr�1�~H�{C�����?��!x�V�D����D��7Y�������H�H_������L����^�]e���_f�T���.r&K�,Jkr����=ք�B##UX*��@E���"��x��.�a�=4���&]��\U;B; ����L�ir�N�X[�M`! Y��292'r|r��$B�������>$�e�r�T׊9®�_0���R�*$���e�Z��ȏ��/�Y�+J5� �^�38�Q�F(Y��(�6A���u������E��y0Qc̳�?){K���9���̂�?oYઌ�����
�Ç:�p��l�׺ƈ��.�Y��24���F�O�9�n�J��=-��K��h:�1�\}t�G��Ǐ�'��̐����Dj�Z���3���t��zv�Шv���Uqj��aѺ��H�^d
��R�o��ʛɪ0K����[��pq�W,(���IQq
�S	�q�hf���V�<�̞�*U�#M�o\Gp,*
a��v%[8T;!��� ��x��C9?9�W/�����:�#(aU��-��V��7�9A �J� >9p�:�G)�ƽ]n�𞠆���[y��<}�B�={*O�=��tftLjH���$ODr?{0�`r����y�Z��"���+������m�wcl��D���u&���,M���O���L6��j���%]�!�9?�)��cRV��v{����\߭�a�rԺ*��l>��%`�@hj�Q�OP�f�"�3LA�bf!t-���N��Vɹ;*;��]���*<��(�:��aE��6��MՕz`��+�S�G��J�q	"�}�S��Z����G*�1�?�Ƹ���5]��m0^|��Z��U�{)���cu� �����Q�A�7���FUt&������P��'�u���Un���� x��_�D��j4��X�ȳ .ТM�U��L��Vm1��ma�L�ej��Q�*Z��ې���t�`23���^=�D�g8��s��W��A�z=�:�	�p`� �[ ������h������� O?�	 ��5̉1|���%�G��g�zO�����	(�4��Xk�lCX��o�5f�ڶ�Ǖ�`�`a�6]g�ST$�pI����nbA��|$\g���HA(�2)p���(��G2Bk�x,���Ԑ�N��F�-G��L�>��X)��L8I���:�lNX���>�+�˟���Cn>_%;��ثw����4<�R=���RaS����"?�9��VF��a�����v&��}��#t��nj	͢5���(L���2Jr˞�*�n� �j�M�CQ��5$�`ɸ_�R�>���Jk0�=�z?%�H�FӋ��ʯd{�a��)�d:��^+���0��ۏȏ�fG�@���*�ER@�iS��?йAŉ��C��	�;���JO�@�d����,���}Sst���
_C��3���||���gV�˦�wq�H�S=�fP�5�	.�l=�"�z`��1|rd�Z��Oe�[�.�i^�7VG�g�9AMe�A3:���2r昣����V��&o8LWr��Q�� 56���˻wW�6=?~���&�� y�j�uZ��4�l��_,t�H�9��n��s���%s��e^�-U�_�ʋ2�J�
�v���w�ϴxV ���f�\qp(�݃2�N���z�E�������X3nϯ�[9G��T����׏aͧ����� =�4<���E�T�f
Џ��D�d���L#\]\<b&��v���L�v}�U3OA��Q�Q�F�?�r�K��Bћ�*����?���x#�a㤅1�}�Qچu���'����Zo,����u�ZCѹn�i�Y�Z3G��5�1��
g;�>��UhK�**�*H8 �o&�NA�0c���|�(�-�����B)Jh��kٮ��@u���flXT�T�OmTd��C�s���y��[y��[y��{9Kvh��UW̠PR�����n������&�UV*�-���]��ݵ��	|�%�u/K���1X� @=Nc��M�V#��B�����ʱqK������=�8�A�}X��ѽ|�z���cm�Ȇl�T|�fV�it�*so8�,⶞C����;��J��X=	��XkF�m��dQtJ��{e͚�ld�$�t s�J��L���@��tڛH3&�6�w]�]c=�h�kĢR��]�� �`�@�``�6���H�j��u�ڥ��p������2����	�Bk:��ܸ���!��G��kY|��(u���|vpH�q �5�M(
�Z�5���ɩ�_Q�32�JN� �(͵0Ik�
}0��>������`�N[4\�Z�Y��-WO�\C`��U 6-P��5A[Q�4s��l��ep�Y�FY���=�Q�E6v�+�4���w�}��Z���� ߥ�gg��Ĵ�xB�Ay�Q�~H�@+�]d� �m?(~0f�4ځ���"��v(-�MP�����3�:z1^P[�|�U/��Q�:-�{��BwA!�dS�A��&b!�0>` ���i,a����5��1�z�bT�5��5��dCi����#����-_'@I_�����/��7��?�k������[�.t�ѵ�Y;��v�.
������y�!R�3�H������5�oo��gq߼��Q[�N~Y���{�����w�3?�7;�ē��Y��a(�á��;���Q�D�:𵤯U����/��G~��4�2P�Q��Z�*���?�(��>H�aB�q�J-��.��}ڸ��?�/?���lnwϢC8G����o�������̂MqT�q� Q�Y�̠���߀~c����K�7|5h�?�3���U���X���}R7Tqa��r�Zl2�"%.�����4W��=(5���G�iT�0��Y+Ů�,~�6�.drwA{)t�T3��#U���]�	 �dM�,��hJ���O�����q�v��ԬC�#Z��Q,��Z-l�m�M;�v�Ekt�UC�7�,B�C^��A�#d��p��!|:@VD���v��j�O���X�9#�3�2��Zp�:0�S��� {�s�! ϳh����Z
�l-�HB����0���g����� ��#�!��W�xvE�B�2�f�@kVXf�̒����N"��++;\�^9�P4�i!���i��ݴ[rϙ�5'������jA�F��j�qf�ڮ�G���j=?o��=��Z���Ͳ�s�]Y�є@,���	
V��.XƪS{ ����-W��f�%DM-��&���+�8B^�XO���5�(��'��Ӻ?�Ӄ�LF��:;9���T�)��2���N�SQ�'2�=Ԏn�Kޯ���\�Tȶ�0�1��ߙ��=�g�_ɷ�� �^���EHJ����;�z*����Vz
��^��O���񟡒 9r���9�r|(����nd���~tE��8o��!�(�`z4UF�$Y�v����|���!��1F%�$h_ԧ!3��0�G����Nhq�l��"&��Q)kKጒ��l�RU&#�b5�����K�SK�8�zN����W�u�uk"M�d[azAʨ�G<�m�
���@�u�q��H�d,���)��߫��z��
l�l���$]��{��VIy(���s��,�8N��l�j�#�Z���%�|��b�}��b���unV�gb�����`a���)1�;��ˇ��BX����Š�@S�����}�'���ya�̥2�x�~_��[���Z��׆Y;�Vi����&ݷ!�<� t[�,dS�NN����A�͵wm�a)H�g�Lj����*���Qt�9.��>�W��ʷ߾�Ǐ��*� �����g��A�cA�ɤ�@1�ߨ��6[j��}�x���1j?4iOV�]��`"�* �2Ȧ�A�� +���6�=�%k�pM�P��H(X;����R;	�;����E�%0+�U:�a{	<to�z���N ���l4�J�ҁMݵ��'Ѕ��ސ�;����֟����Q~��G�a� )S@���.��j����0�.ь�,"k�H�Ek�+�X2A�
cʅЯ�kgk��B
�
;�s�A��*�}M�G�0FkI�����A8$�
����A8���_p�;��v;SGU�-�1R�r����I_\?p |iz�}}������6Odgn���q�MGL��7\����`j�t�����Ç�����"?]����iG4!���w߾�
P!Hv�B��$�xR�r�C<�g||(�Ƣ�&{��_���]6�n����i��۵�,�+�SR�r��QL�r��y�$B��K���|��P܂y��8�56ݑ�P�_�I��a��Ea�M�h6t�&�`^���Ez�O��x�K��F,h�X+��b��Ί	7�Ҳ�̊�:|Q�}��&�,
�`�ǔ5-:Y��0�ꤧ!����F&�rAĶA$�3o����t@�g��F��w��d���b�I_8_��df�~�O����b�n�m1X�Q���y����׾����Q��i�M�z�5,NG��3@Y\�2^E��)��5l��5F�y�"�5��͔�Zx]�[�ahG�Q~w�)LL ka��v�9nûi�?�8�p��7��;�xTɱd�t�;��8��6-Z6�@l��yk���\$��\HKsVt���{Ym��o1�J�ʋg����󉜝ɤ
,,/�gkw��$wr�I�n.e����?J�E������;BB<��:��Y�7;���������/�ȓ�/�L�(�$�壒��"R���XѮ�'�`���ɨ8x�V69r�Ar�K�2��A�u��L���F���9�xNB�/���N�N�ڂ�m}�� �7���=;��Ё�TTh��5�t2_���pj���[:�*'��!���R�4:�9@�Q�:�G��m-���W���T���mЛ�9h:[�5��"Nbr���aB&�5��B}_9��0���-��*pC�f� Ȕ�{FG�-�̕l���5�d%p���*�����Ev��,�������^Ώ���ϭ��/d�j4���D 1��7�-k:��I 0�R��~�*Ӂ=��k�0�b�9>>N��r���	��h���-*�m��B0ə�?نe�2�I��]��ߙ4�f���g�JY2@�Hq[���˪d3���H�_U�C��i�%-�X�J��j�Gt�qI�z�9V�������_��+��qkI%���(�>����[i��b�'il��v��74�N�5M��#KA�'�,d���{eu>��Jd�*��P,��.�-	����g�.P�[�?[�Cb@@�@(a����:*��^<��v�����Q��18�� �<e핢��v��,��-�haR���QZ�| L�҇�N>�]q���?���ȟ��o�S�>&`�+k>M[]�6"� 5�F�S�`��2-��@vN�I XZ;��`�D�i��( ����q�X状yo��[V��\���~.�/A[T2Ը�&Xw?c�!�Κ�h<�ZcGA��	�hF�ʑn[�~M��tsg�M$?Y�Έ��u��{��FGPv@�݂�#��J���?}r��Q�f�Q����gy��=���?~D'�+n�H���$���UH(��.cN��x�*;8��8��GR�������3 �k�<�K�@�/�(42z�P�eMp� k��=���֓���9��PJ�ҺE)�����5�Sht�Ƿ�_���YH�5>kj~8c�J�����)i�G���"[y0K�1�b����|M��0�������,H�x��i����j!���um�����t�ٲ�sNX�J[;�6w���Nc�L	��8�pbhv����,���VD�}�g"r4j�	�h�f�O3�"�'��f�t���7��IΩ�|3p���|u𽬚80������E��.콉5������<]��ʞ�jf�B�c�� �9g���N�YT�'8�&7�=9`ǐɂ��ё�# ��m���i}f3�Ջd8A&Dệ��l�-�Uh�b����p)j�F�kԳY���&��{�jcSH�^Rn�M��?�  �]���j͗��7��L�N�P���ّ<�8��O��:O�>fFr�%�?ɖ��b�XJ�^0�5��bM�J�:R-&F�YA� ��3!��:��l)�	��N/�ￓ����7?���S��3QYR��2P�6wn�Y���h�`;�v�( �L5K[�`�	���L�/��u��<W �F�B>~/�NI*��U(���)Z�D��N�UVEB�Wh!S�z���\�4(�'e)9�� �Q%��L��	`��n��{ �->R��~/P$��um����R!b���F�)�(5��ʭ�q-�&hp_�PeJU_��j�X�u1 �͡U���<�P��j�r�Ny���B䠳�(+�3"��"O��$]`0d^�{x��sۂ�e[Ӊ����N~�����?��ꁴW��|�p)?�����>h�	#�U����>E#=_U���^�d�(ru�a�n��WZ_ ����}�v�Ec��ې��Dag�L[��lǾ����<��Gq���X��o�ބl�Y�M^�fV�&���T�#{	� �������
��6��{/^��ゥ"#�>���;��l�{y)���t�'�
MZY�ZnŨw��XY{�g�iSun!����e�!�O�=��G�� �`Y���o�s9F�)A��e��孓_��^�i.�n�m�a;d��M��O��@�JKnL��L1�Y�#��T�m��$���GѳVF��7@	·w�hi�ˇ��!�_���˟��T�D��N���Z�v��62Xl}�r2#�p����LP�"��UU��Ni$<���y�����X0�H�DY-�=����P��	+{o��'�/���,T;����Qq��	i��(�`�$��S �%L����k˾��;.�t��F��G_��0�J�gʒ{����h�{
K�q��<���)�37���������UYGrz2K�k+?�}+�ӟ���rww'�(&i��Gl��vr~*��|a
b*�j'mT޾�dh4�V� X9�	��Aj(�Yꍴ�{�XEC��a�E��D�0��㳄���M�D\��W�ËeP�M�V��d��y���i�_�ns�����:ƣ^S�P5�E��������A*;r�uD���(� #8�bsFZ���׎+*AG�(k��@�<i�s���N��#E"}d�H�wy/Er�������*a��p¿����$��Q-����4�-��x��O��ZF)u�a���lC���r]��T�j��t<��V� 42e��G�j"��u�QA��h؀��\l�u�EYO��Z��k�r�&M)|gј������|Z�dY�5�xO6�<�!b
�U/8��ۅ{����T'�N� �Z��w�!���a{��͎�?������.����p��Gk+�S�m�%�4_�5U����i�ک]�@]f��L2VX� �`�n�@��"�]��5��3�h��x&繜�ȭRuI=9RlD3h�eF����z���_cU��l#��f����!̑J�����5-C����a��G�jv�0nZc=Ś�� i�
2F�k�XB|TEn$A�r�ݳfvT�R^�M+h��{��g��JDΎ��7���߿���<��g���AХ,����Ý��H}�5F�"�t��;��t$F����^��-�꒶�Iv~�i�*h�'�����?��?ɫo~���s*�-�Kޗ������ߗm�.ʁ�6�u]�����t�øl�!�^F�YDSb9�V��P�i-w ^���j��_#�er�@튁s5f;6���z�5̵��Ls5N��Nc�L�%я�8�4.���jk!.�^7�4skٝ%p5����t���M��ɑب��s���y�#H`' ��8t��/���:�3Pg��'��ڎ�
�5�q��fhM��lI�yQ8�FM�y��WF��ȯ�u��V��xĞ��>z�x;��m�"-�!Qߣ``�5�U�d�
���͟�6yf݇��:�\��`��9�V>�rF����^޿��^�I��o��SJ�E�����a� �4ُ��t�#�+g�"��G�j@ǔV�Q�'��R |N�&���l�l<�9 �!ˬJ�!�Ss�	W�s�Vx�Y�1J l,��>��6,n�F�~"�ߤq�Cq�IZ���J�m�8���<�M:��ۅ|���OW�䤎�NKPj�4��+�]0��h�� D���/f��6�ÀC�V��]c�&��Mҹ�Ҿ����1@[K�H�e����6��dsf�i@��Ny��)z�u�d���J�AǺ}�FĈj���5RM���W����>�'T?���~s~q*�_��;i�P*��-A��?����?ɇ�i��c��,���A�t���PԈ�8\҂�5"2��*�X[�`^�Eg�d���j��a��!ݷR�m���Ϡ'��r~+��,��RV��	p�(���7����>9Ns�ne�>MG5ʂ {���$�7ų`�Ɖ���=��{2k�B��Y)J���1.4�5�0���B�Ae���K�4�Æݱo���WBK�[��;e{���F�GR<������;��1'�^>�i>�ֲ]&w���t�"�� ku���������W��2G#k�d:!Nϖ������\�G�X�t�������.u��C�������?HĿ�y_��r�΅�8{t!�޼�7�|#�1�㷦|��"aJw
�=ͩH��_>�{8�a���c𫿇�7痈�}�ޤ�ϐ�����1��#���=��D$���1
D�:��;��ҟZ����+4�Xj��":#�h�-Z��ĆM�Ա�AdE�,��Z��%�	�ˢ�����oѬ0RDU�<\zV(�?�������p��fD��)UA2�� jA���3��o��IǶZ�рT:��R�2Q�2	C*�1�C�E贁'b�mH璀��i�%�W3��X�S����	y��a�Q��(�!G�@0Չ���}��?�[-�q�o�"�a���t�i�.�[Ϫ������h��\���'��U�d��@���΃I1�0CK��d�7��(\�Y?��,�� P@QP<џu8c֊�f�U.��担�q�)b��!X}�Sa��k0���\�F��vou��#\�y��Z�Zg��R�t�����X#e1:�X�9�y��P�P[M����m��X�yr�/���G��y��Ϟ>��O���`L�Ӈ��mW�����c��YC�z�W-�/س�O�.���C��`��C�{��d3&�����ʫ���w�� O�>g���V7TJ��V�{�ldJ�:��3�v�����Vf�;s.Z:u�@�0Ƴ�.Ο��ݍ��8��d��Hf��b�ϊ٨�Z�C��)x�<c��m`/���
-E8tT~�c(Ҁ�zg�h?����[�]l�n�!�p���磔%͖T���� ���	6?
Fߕ��'�#�G:��i�F�8�,K	�5�C�j�X��h�W��S�-��
�ISݷP0A�u�i1�Nqk��tu�r�A~T@�y�h�h����1#���M�����������  `mO&%?� N�@�%$�a����LJ"!˧29�PIn���e�s"��zZ8�d�A��~��ǰmY�5�/T,�D� ��X.r��`�Q�d��b����t���*���E�[��&Pu)�o�q�߾{/���e�\�<�R�nXGf���&�����B*ַ����C��-�PŎ���|����LιR�G���Rf�ϯ��n����Ff�˩J�#�� ���	�@�'QwV��ـ`���H~��w�O���?��<z|.ը4�FNO��Yu��
&� ���d��O)Բ޲�A�����B<���(P	�偸���:���N�5��A_���5�P��͓wmg>��5!��l�mS?&�%�}-7�?�}�*����rg{�Zש(��c^�7�v#.T���.�0(�������DcZ,�#� ��n�E�����`�i^�������|�!�;8�xJ�L�{Vr5#�P��5t��jBћ��`&�3�|2Piǩ����t��}��G#D��s�w�<��lS�@L�"6��$.&5knV:��f���'�������?Lݪ߾{'?|"]�0�B6���@���;��?�����[9J��@}��W=�R��[3�!���6t2�y�����>�`"���L뫇�G�~dWǋ��\ؼm�5W�>#���,�j���[�V��juX����Em�R�zԌ���S��@�Ql�Gu�V:-���bC��v�ӳ�y���)�Ly���5����l��e2 pf�J��@�����iYj�(�ƫ�=F�c��vE�m�F�mP,�X�I�8q��a?8�1��>#T-��Kc^�%�q`7�Jr�h:ڦDf���<� xp�?�8���?��X�)K�ۜ�y��W��A�$�8O�۩5��Q��<��Go�~�1�x�LY�����fR�!��*��&T���q¬�nIр���ͮ�������z�@y°��k���J��#�<�\���|��>W��wQr�R���QTr��ZA���IJ�)���<��6N|�*��ٽ.�6/Ο @���T��e���ɨ5R�~��+�g|)(RYf"9��
�f�_�޴9�#I5��< $n�P'YE��=��#+����dewg���n^u�F���U��#����2@"32����LMM-t������'����3���s9;>d�-6���F�!k�,��!
��� U����l�u���ZH���(���!�P�7y_8��Ϟ�/���_����3AM%�U�=��n}Ҍ����S
*P8
���RHm�e���T�㍩om�ȼ҆����u$��c�j@�臼�-�ג�#�/34��#Ԙ�V�l6�>��Y�v`C'80�������>�I͋�L�h�CE����(8r���뻅��/�� ����Y�D��V *� =�C'V���GTe���G���a$�s/��r(]6Y��AVm�|�y�^E��t��(�D�ٯ|^#%R@&��n�dD�	]�����f糩�3�p���� �����A�m��┝��k�W��~<0����.mH�P� �EF�QG��8T6uZ�>i�p7��שc��ޞ#0��,�A}�����h�麋Ed�i����ֶ} �u����ւv�̪Y
��"�;ŏ/�/���Hَ�y�N��{��/G�֭fE;���9�f���7��A�b:x=�*K4���b��m��|���a���tG����dY�
`omfj٬�E��aǬWb�KA���	V�����A鉰����l�N���S��?�����;���0��@p���QU}��)�{�@2�����Q>� >�FF2���[��
uV����M�ƣ�4��ep�6ʀhd��Wk����|ˀ���=(�ݼ�����[�"����^���!��1���J���T���Jsfose���������&�w���@��w�#�|�C���@���>�*�T&�v��C_��P�I5`^��'�ul���c`��Ӗ�6����XԹ1�\��������O�R������A�Z��Xl��;���	OÒ7�9�G�*�������__��N��n�º��Huov(GG�r��|���9����]���mM&�ZC[vN�*���a�"IA�S��s��K[���,c3�x��u)�1iT�L��
5�<?�`���(�K���U︻�E�.��5�<P�~C�uQ�;3J����S����LQ^�PxB	����?��([��7,-$��-��T�Y���;UJ�
(J6���*59˛�4�q~$���p�Z��A���ƫm4��ҕ]�f30�jn��[�\E�L�Y� ����Luݠ�YgG</<:(;�6���D�y5&�[ƿrTb+�	F#�\<���6/3��7�灖>�2f��0�s'��4�?�?���WP��o�dC����KF��qxH7���s�8�-���jD��x����	Q�v��+�F��k6�V����,Ⱥ���������VB���0��\t��Q׻f��H[TtU�p�OW�Z'V��i'1��~)0�͉u/ҫ���C9�e��"�֊z��i����*��x�6Am+��}%-�*G�)��z��B�<~$O/�d'=�y����o����XЕ���8q}x�GjQ*~�m��R�����AI�>��n�/�xH��'/(t���K99{��}UO��\b�tƔ���[�s�S-���9P���Yp۾I�iۏ��,���<V̐�������~�8J��b�^���0�ކ�ފ��kɂ���Ek.Ĳ)�� z��	B�c�'P�����4�m�Ytv��Ѽ9�3��Kh% JRt�@N%�;��8~J�&�U���-h��q� ��~RT�2P�E��f�@r�Bm��D��1 Z��%S�8����4��L��"�gb�Sq]Fe�rYr�{^��z�Z8�2C��2�1F4�T��Uᅅ��e�TpAA����t�K�`��*�Φ�e�Ͷ��O���EN��)1�[���X���Ա�>��\-�m\"� ����	�����(�)��auS
�Ϲ�L�C�� 1 ��v"(��kKP}�	2'd�0�Ttܰ�&��z
a�t�o (�X�m� �0HK���z�����yv����**QB����m�^��0bfyD���]mH�m<b��XhK��J�
����g��o^ȿ������y�T�S-�J1�u���9b�A��r�y���Yu!wy��ڕ��<Zd_j�E�i0�������+6^���>���V*�ïZ�m���(!'a Muf_ xHjkQ�VQ�bC�G� ��^��{�·�ZIt��u_W��FIuG�DJre�}�?��Zb�?��|ŹfU����U�����;��v����h[�B��w�]H�7[�_ݑ)V�⬙xгcD�5}d�M��⠨��|z]N���0%���x��m�O�˰W�c�P����p2�T�?����r�䮯n���)\:�T�ʋ��N���Grqq!''�����>���c"Cw��|��JV�G@Jz��b��9�j�)�0�M5Y��4蓱M�����!�#���k76��\oB���XP�!����XX�%��MԆ*�ŵ]�������M�ʨ�����A,$�g�!�p������)`R��N�t.+=Q�Akŷ���h�o���m6�{;c�-��P�B���.;�y�jW7�0��Mu<�JZ�*�hV5;�G��Y���ѷ�y�h6��@T(PZCK�l���r@��"��̷d� �ڨ��fM5{�sjp?�p�2J|#b�TK��P��.t=��-����xV.��T�@�� �E�S��u�\w����nW[��O�k0���sV'�7%;"��t7�W���[��Ւ�#���~|����b�9˺�F�6c�͇A��w�@@3�O�éz���֠�u�q-:�/�]��(�x�J���+p���E���)�z��M�l2����T�1���:nĬf��e�!��Ge}T����XU� H	�������'�œs9=��������CV����C^ח*�9ZCvkw�ʲRLT��lR�����0�O��!�[�8{��/���9�:8��0�	��w!�� ��kc]O�:�uӃ$.��x�8�eGM&�R}��ĕR��\���{������8�7�/e}����-k$o�p���e>�F�Yvn����������!�O=�]�z�&;#��ԕ�h7�t�1�sEn&�tt��"��kl��B��W��(�!�5�����`cQ�-'4�M��+}^���Au��e?&P˓)�����h��l{�`��uZ֚=�`A�bZ�:������u!j0/b��J����'�a�l�
V�������3���*�:!SD{uMdgw��!�0�i4�RS��ޔQM��b��Aa��)�I���׼?p�ݏqa�}�v�o�Ew�PZ��G��ivԬk��P������Q� 5����{�����=�Ή�w���\��9	�,�l�	���*,�&Rt����Rp٩7��˟������ɓ��<��N"���u�������YD�����0+�S�����@s���P~�����˷���^�_<����-Ǖl����6��GG%�֤�ɾi����F��ϴ1u�&�a�Z>^߳_|6�j� ��n�a7�fHQ�S��.{�a����l�R]ۤ�ژy&y�䎾���9�꾯"�U'�k̞p���Xy��E��jP��l3��&I�i?8h5��<�^�p(����GH�k{�v���f���ڱ��]=���z�+�$2 �o�����h��z�+Y���0o�Z���?`�u3��Ɨ{?�I(�^��%Teł0��lYD��i�����V@��2�4A�ZM0�j#?~,/_��g9Ț��Q�g����v'<&��G�y�N�d���0���˭ �w��_�1R=��m*��H*Y�P�@�=k�)[�a�z�ơA�w�hBe���4PV�Oa���O�lo&'ǧr~~�P�/�lmH�HF�3^��d�tZD�+�8����qu� nn��~LX��(�&��aC��������ˠ��
Ơ�L�/��<�!�D�x/�ҶL�^�ր�_)dȠ)z��c��L�E���P�mub��9fp�k-D�,�RTd��f�\J.AzG=l�����^�[�2��炜�J�3�zp��`o��I��!ۧ�}�[���ch8��[�W�>J�O#Xv�������@�E�1�A�Y��/�mXC��*�$t۽;T��ʞ2�p�)#�,dӳq||� �����v��K����ߐ�UBwAд�=�Tؾ�.%+���*:�=~x��րD�����T�Y�.�Ń���Q�kk4?��TT!�"x�vv��p&�����P��NǗO��x=pVن�����������,�#l��f9�b�?� j��	�Ŷ��h橦,x��b�LR2��z�����'/(rqr�$?��5�c	���f*K�&ƾf�dU������`k��#�%�('_WN��ql�ܹո!@�	��>�/��y�n�m���:ͳ	��	Tq���[Cf�L�B��3L�hbh��@�~,�c��j��4۰�$���vs�:�?��~���E�����γӹj�h}�D�kUtFI5���d���
'�EY�*�5j�Cd�5��2�}��,b$��
^P� 0eH�<�:�X�ΥR���(�"�t�����C�M��{~�:s��F{������ֻԥ\��W�ɪ)�~�؃�����D��<����N�]��������`߼���v鞁�^޷I-�Ծa�E�ڂuf�ރ�%P�nn�$���=w��F��� `F�^�X��RFPm6+Y]#k����V�����ۻ�l������pͲ7@��2lM��Z�W��C5�Ji�[�pJ��ё����g����a��;y,� ���*%{��Ʋ��^O�;I_߫׏�wd|��f��9����,�^=οk���ȱ�5#���}<��g�u����U>~6���#�]�v�ًg���������w?��o>���N��A{��n�[Z,b�5F��k��H1�����}�P �eƬ���}dC2&U*���&��oE��pZ��g��轧l/4J{,�`hyHo{��c��W}půh�r%R����}��SK��2�T��?�`M�5�S�8�z3�~e���C�v\Q-}T[�Ej*������L�e�&�u�6��#���T�.0k^WK�/�u�5Q@�(U@�5�q��'�����o|xt �{�%1Q�~�:���g��JkuFu]T7��!3F!4�����M�k ���W�ï`NU'ik���O��^��ő��vg��x�uX�e��)�1r�Z�dh�X�6�0�)�$/�}�_\�i�#9:����x	)����eѮH!B���餡-Go�U���Yvo�,;�@o�x�����k[Һ��>�pw��WlV�Jv��C>F��l���K�oƉ����莩���u�ŭ�e����("��Fn�*�&�cn��W��p�<>	>�Փ�9b<�.�9�X�*��������R;�0V~2�虫�g����_�/}���`ϛ���@C����@�؜!���Q��A������pP)^�l����c�}|�/�k�4Ô
b�V�lYx�:�R�QT���t�+z]����;�>Bz�itVܕj]�tl���ǳH�q�^�Q!�#V������#[9�	��5\��s�������xrr��]=�g����`*�}ί(�:���;]h�e3�E	HJ�E��hm(�	w~�����ѴQGnxp�зd��/g'����39>},��'�j���Z96Eu�h�8URU�Z��Ox=/_��ӕ�f3������D?� 0Ȁq������r���^���ↁl��>�K! ��S�\�6��W�[n8��r5\c0!f4�@
^k��5��F��^3��N#w] �]ݒ�z)�L�ܜ�s�t !���93�M�T��תfCP���G�(�]t�r[�ꨓ�}"1T�i��a�5�����"�U���7v��N�7�[�\����
.�m�F�-9���U��������}/@0Ej�����`i��PsR=�49d�!����}�+�0�۳�]
��Di� ��Stj��C�q�>NȘMoor�|���Aޣ�h2���N����1�f�, x�ʭ���`ᅛN[��L����Y˨�f�=|��%�
�L:8Oo��X\���)Û�+���!p\��N	6�1��v�d�����W���sL��)��̫�P\>=;��/���W/�_t�~\0����H��_��Ї��oY�ϛ���a��5K�9 �O������"y�݄������_ :;;�Y�u%��Xd�-D�e��0u��L��S�f�E�LJ邍52���U�}��|t�JAT-RPC[�h#�J�0�ِ�SClN;�_-]k�-��T6��<��b���}�z@�k��0H���k��1�#��vPS��� ��&
s��@�;�~���7}a$��-��!���(A�;/�|�x2��i��ly`j<�rޠn��}g�0����+2�Uq�5�v�w�(VGG',<���3���%J��mH���(3�>0�	��M(��\'>�s��{Li��4y���Q�Qq����g�  �T0_0Ƞ�&�uY� ��ן�4�����`Q��C�7�ƨQ��`woJ��8�����`W�.����r	teN�����X�K�MeM)��NTi�ֻ�[��N���蔟|X.��)b��������*Nk^jSgt1�Dĳ�T��7@�ńC�S#א��h!8�}ӹ\G$UY�Z\�(�8־� 	��D�E�l,U�F3MDL��_��kg��#n,��m0s>	�S�C���\�П�'s�:V�:)�v��W���W�B(k�|�'o����jVy���Ҙ��M1].VEU��n�Rd�����5��@�5%�F�Ѣ
�!o��u���]䱃vW��}c�R�`r��G�u.S�Tz�B�k&��?���"��8��AF:�A
B_�͑`{���XΡ���Ue4 �W�c2�n��vTzl;'j��JRv
?�W/�˫/�ɗ�.�p��7�������~G6�j��>�錬�Xe'�zH^��&�s�~�Y!�X�M
ꓦ�Km��)Q���������s�8{J*^5ڳq
�X�(T�mA-�R���G}�,a� (Ҙ���P�`�@?u�1W�Pyc}�F;rx�H�/�ʇ�?���[�]��1���zv�Ҍ��Q̸$���N�~L������k�Y1���~�=�9Vt�z�Q�i~�.$�q��s�t�M7r���ۻ�<�<�RYw]iS�eI1�Q3Y�����P��	z��ZRP�"iUW4_�h��_b`A�v���1B����b�7�M� F�"z�N�S���z3���� ا��d�%ܑ5%EQc�A�$ť�\���t�췪B���iv��Is�k����
ŔD,P�g��j����}	��XM��t��4�A쏅:)�>ۭ�ÜkkmsPx�m
��!�	��(�X��u��ohS�Ze}�:��\߭R9;ͮ������з�J�1����L���x��S���f9�Ѧ�nawd�vIM�@����E��0{,;�5��ls�N���W�����Z�="�S�c�Z
�~�V~�=\�_~y��ŜA�lv�$ ������G�r�j�>��u��k�E���ގLr`�Eȼ�A�M�TI-��zq��d�j����K) #�hf(�߫���-��6�^��1� �AlX��*���n�tS�[>��UQ������*ng\�wD5?�S׸H��0��:`�v:�a��m~�k��;e9y-�'��
9h���1�ϻ��6GT8i�G�+#�Pj�d��SDw���{C4��j�Sh� -ʍDYtB(%�Rn*2 �d��
T�$����8��y�����E���q,|�M"h�:�;pT�J[�Έd��ʜ�7ٿ3��$۰��r�I�?S[3� j6%��L�b�XCI��ĩ��x�{]�t'L9���Pk g{9�B����I6�'�%ݟ�$p�̆�N���8ݵ��R�&mZ���Q0�"�+�BM����|�������L�֊6b.�6Y�%QJ�ܠ�q�	%��c��ET�T�1E4����.̾h��a!7T�df4M��\��x+�ِ�TJ>1��ȯ�ɧ��0H�!x/5ۨ(���A�O����E�:̓�\�w��\��s�.�{�=����>qRQڑ�y��p N��d��J@�%� �����i�o��bs�\�� ����KGz&�8b�lvI��yGn������:=�d��O�.�Q���~��������{s��١�3ꐑN�N�7��-5��c9���#�"k(l�_���(5XV#�}+ ����)�
����`Y�ͦ����K`=Wm�:��<:?������W�ʫg����l��cr%w�o���� ��5m��+Н����_OP�r�oq��4Z�Ջ��� �r��.�Yw����#�8���gr~|�w�`�N�QX|��Ak3v�P+��R%Kdk�;�n��v(�s:�S��K�f�h,o��w3���$��>���r;�\C��E�ԧ -b�4�$����y,_�t	874�g��Zv�9���sL�����0����a)��(nE��dG����(���A���D���N��D�bk�����o[��5����j~׼.87����4�P��o���x�r`���9m�^�mtq�b����g�ᓦ�kH1���^Q�̀F��[��hh�r�u���'Oq=]<>�ã}f] �2����4A˛l h� Ѧ��%@��k�j;v�f��(��_��)�90hX/�+�- 0��_,�+m��z%w�5S�Z�9��8dRH*k�ݷȡ�U���	����։;�x_�@�D���>��Z�tf��AeO}�W_��A�S�0`�2�g������;�Q�*�F�4�v�=
���,�z!�ԃ���￑o���\\�|�?j���+��?���{���s��^�T�F��=ր/�1���:�y��Qn���G��?��\�L����<�>����ﳝ��Һ)�J�lLhI�^&X6+��� '*sA}!�"Av�c�&Lh��
�k����<��){��m�3��x�������F�#U�u��:�
h��3F��CT�. 6�N<�꺸)��[��P޷|��SR��=s�t�9@n����At� �@�o���G���7%�Qn�d8��Uvq�>))B�`9MG�,�� VK�1`P�ӑ"Q�U�6<{�$O�/����ӧrzzN�|�2;���XhȎ��0f!�:-U��p����&�4Ca�vz�wl��4���
-�w�÷�O�����U�����q��1Z�@�3����z�/d��z��]��ą.�TY��L���NvF�g{rt�O����=�����
w(ww�h�F�uNSR�f��)��ih, Ⱥ�W�-��M\e����
�@�@0�̣�Q
a�1�-�D)�D\A��xӃ�ib�<�ǚl��.�Qt�-P�QA6mP% �QYD�)�
t�X�D0�#�!Y,��A�*QF�s�Q�n�0�O��q������]cl�*�^�J܌������>��_͏} U�im��8|�~-��c���r�J,������H�Zu6��e��_Kl�;�i^?{�A<�5�Nibk |i]@��72��i���E�A��f�����ڂ�;:C��n�%�)�?���m�%JT=)�ͭ��j�S9M�kVc�b.��K��Y�.(��b �R��VA��ŹU��ҵ�|��Dm���2X�iM��Wϳm�Z�G�.�A�k������ß���g٬��R;�Ԍw�I��Q���?r%���w^C$��|�)�6F�e�7��S�z.(�>:{��ׅT�G�"&*�`�ƙ��ᰪ���뷾�z�}��U��m)s��s�d�_ls�O�������w�� ����0;����l���N�t@]L����,�PH	��p
V��P�N:�lñ��1�Ƙ�����a=�Z1��خe��0�y�QvXSv�
��ڜq8�lI��uPvT�Z�*	�wLA�G���� �aW�uO���4+��ByH] �h" ��EY߭��A��.�wP�d��"S]��#���b��Ȇ�x�vOX�9&-Yd���||���1@Ԥ�Y��8��i7��! ���^����Dsh���w����������A��cruM�w|u��*j�+>�P�����O,m���`��s���:�QQY�����	� @V�8���Z�5�+�k��O�=�6��˗_d[}̌U
�%�9�q0Q���� h�yޏU��!�ɔ6g�Z�qzrB_-)�1�	��"��Z���?˿��?ʏ?��{�C>��9k�R[��R<a�\�b9����r�sC���Cd'�����=��|�n����'�V%��S�5�f�Q>]P��&eL� Q�^���*@M��{�BJJ�@�}���5_�q�]��94��v"�$�������eU9����M�����9�Em������ɖQ�����A�6
����̗�붾Ђ�����I{��1bV�RY\q6��V��J���Mnt�28�#ȑ ��t�:���tvJ��Ⱥ"gp~v�h�J"��
�_}�R�ǿ~%_~�,�� n�c�=��M)jSw�^64`	�V>�)hT����E��r6�Ĵ�c�����cl�ש4-�S�,�jP��_��`��T/�v��q���ܺ����7�ЙMv�����h�#@���u�̟�ir�"J�Q�@��\0 @���Y�)�иC���v�+e6m�`���I��f){@wq�@�w��p7[#��衰��hZ���)]��N�L!_�boQ��N��eB��zC�4F6r�P�ԋ2����2w�jPT?U�!B��Vc@��.���T�@�>��A��*TJ�B�q�� ;�W�_�\~�t�`�6i�/A�yH�7Q�ܰ��fs/�*q@W�m���Ф�JWJ��u(0>��z�ҳ�^�u���N�0:�v� l��-QT���V�-�VG-���*]�$K��46��#Y�QL�ԛYz=��#�U�E���6�P�^c!J�Z��
�Mi7+*�!5��KG���3DCգ}x4�r��A���c��[���ᡜ���TN�ϳl�V�x�Ay�
^�y��WJ��P�#T�:���fʈ�G�mh?%���)�jo,��Q+=��]�3��0��Z�=�qVF����2���-��9b&?���N��=c�s�@�èe֊HzvȪn)gy����3��?|%�~�J.�O�p���4���dq�Mʜ��8��T��ZК&��J��q�JU�ƶe#�Ң׵�`;��֚6]��t��}�?y*{�O��?c�p�U�"�`:Iɤ&S�+�o��.�-�b�S��_&�����l؏N$��,qWA���e{3�O����b����ۤ�����V���;�p�(�h-���U�Ro�>A�ȑ:���t� 4ё�FE�F%߫���촞����y���k�����"�{y���׌��E;���q�c�����(��m� ��ڠ�|�ePn���Y-�ltGewޯ�vvՖ@}�xW�(�R��Zl��Fv&S�*�ڛ/�&�n�G0З��DQq����-<��5��i�7ưa�Dj=�$!z��'�G'r~z������۬H����z�u��;��7��k}�m�<��bT��U^�P٭`��eY�cP�Y�|�5�'�!f9��kؗi��O�>�P%�jrh���׿�6DpP�1�#�2�l*�1`IRʶ�3�3iI$A��t ;�@_Q���p�R�#(�fwL%���]+�s ��L�a��O�/��r|xL�K
V��׷�wxwwM�iԐC�tYr�{`�\��=wr�3�><�9�`������ײ?S�χ$�������䧟�*���'�5P�T��1�*�7������+��
eL��s��� �.DR>��[���s�5�N��TF�[�>�@������Lg�d���`�um�;G
�N�����{R���6�1Ԙ��ӄ1m��H�v�m�jm�%?3�S8��;9��/Z9^R�mVMeV!��K��|T�D�ۻw�n�^�./���]h�co�ز�E���%x%��P�sS��T1�,�&�NEu�H�UdI�GF���`Tᖽ��4�@A�􃃡�=�,~)�:��J�(���r�X��x� �
<�u~1�uf��<{�T^�|)_~��<~t&�e��DTuGU�p�u�E�Ν�H��4N�����nP��J�
�_R���5���I%j��9��y�>���[lNnä�H�	v�Q������^�â����Y��T'ѣ`$C"�)!�����`�(�0B0Fcl�y���� k&G�57��+�QXj�d>�MPV:�- ^�aX**N%O�V*���@7���t ҠR��^Pdk�Q���(�h�z��h5�Rl�k�I�z���CU��@�QfPd��E2�a� ��@��~�1�����6�XXi��V���RG&`S�^��2�·��r��o���b?��$���됦[6��%%SEG6Y�d��RO�u4�K��������l`��B/��:R��)j�:��ҟ�?�T,q4��>��l���AyS�/Huݪ~4�Do]�^
7�Ն�RcCe�X��ݧ,28��v����ĽbV,���2�5 ���uE�7��hIO�`8��O?m
�+{X�|�B�����WK�� �F<w���"�!���6ۙf;���H����o�)�|�L�d���w������������$���F�6G��|߰����5k��j�*&)S�s]2q�ɓö��SJ^C��7xPeC[2������{[_�	������.q\pox-��A+�d������S�]�ʞ������.p�����yR�TՍ��� u�B�ף�/����PG�̠��BE�7�vGr����$�[fG1}��7�a���WNխ����5�d� *��b�}Wp�h��H��@�Jo#���b�nY�T{!�`��c�����M��N*A�lMq�d�S����^�`y��w�f��ѳ��.C�"������.�X��c�V���T�t�T1�	��R�?i�;=����N�S�x뼇� �{&��@BbJ��N�ތ٘N��s�̧	[Y���X���,�1�X�� ��d�֛�f��\q?we�U�vmD� q�XS&�Vt~&g�dBc�c��w�)�����]��h��J`�0Z�LH��?���&j�N�� �Y�m����h5s�h�1Zy��/j�h�
Y�X�:���U�f�"���~�|���L����F=F���V�0Z�T�R�V�����Y�X�~�A�XP�Lԋ���3�A�,_���*om�M���L�fP-�:::"���~>�Z��w��q�p��d�=v��(��[�����{f�p|�,AJRa
�~��'����k��W^{���s�Q��n�5���Pz��Y�M	���,�>@��`�ŧz7����T�j������8?;��O�P��4�Y%:�.��	���;�K"���M��g�����Vk�k'NiC��E���oާi�����#i`��&�I��)��j�J���o�{�'�
�U�t�VV����AUz0�gL��l��O�Y|{t�_�D)���l7�9� �qss��խ��j�ZCՁ2!c�i&V��5�!eOU�PC!G<X�*ڜ�4��:��*��mgA��Pݠ�	4��mkq%��[.4iKs?Ee�+r����ف����yU\���
��)��x`��P��fc��!������(�;�[���I����B2ǌ�&�����ى�;�@�*��p{Y��F'�}A=��6�`N���2/vj[��o���|�s��?��\�ա�]O�W�A%^����91e��B��D�������k9��FCϠ�))\{�,v�;�ܯEC ��Ё���m�������kw�p0��^�ofc<�(}�L�aT�8�L�Q�/�D[El("��G'�O�|����dg$���|ȁ������)\��U�QP'kT���);z�r���9�M�j�5�Y5Wg/��`-�I���uJ3k��f����tg�6�F�
�k���K#���9�����yv��9�K
l�ZY�{�������m����u�{+�O�f���uu���Z�ӆ�2�B���!���>jD���N��rsQ��(coN��*Ik��,�Xb�;㻨�`]�ì�8ݬ2 ��?���(�@@uD��ndBY��m4:��Q3�>�y��2�F�8��fe~Be��F򄴞9T�V
Q����4�{���{�	<G��`�U�Ӧ40w(�])Sp�F%p�bShO�Bh����,ԃe��yF	_P ��]�=ڣd�Gc?���݊�.�#ъS�K<;��9�)+}�a-����j#i ��P@ 
TE�lYkX�1��	�-��K�6���Ď�k:ːfW��v��xĞ�J �f�{�x�^�d{���{��z��H���ɤ��iC� 
��%ڽPaV� p��U���(���gg�����Ԭ�Z��p@MzWT!K�C47^�k��$9?9�_�?��V�o?�������?������k��0��k�����#檫�����cJ��h���Kä�֖�-�n(���yp~|`6��'��5�g,1�'yd6���\���zhYh��3%����n���rŚh^kޛ^8��|��ϡ���[C*�ʯ�W��pL�澿��7kY�� �da ba{��c���\�"8sz�alJ#I��	,*=�l6�"�UQ-��1�^o���V-�5�
�i�,B���I���mb*Ί�7�>&űqH{T.S���%x��a %ɲ}>�ೣe��q�H�E������SK�� ��7(����k�'4s�x|��rr�7���`m���J�Y�d�f��f��ŽRx�g�:6�M�����RrDR����QXb�Ԣ�*13N�tzaD�) �daS�#�7ic׺^p�v%^�.I�.�����Zg���#�Wx=+���"�Q��
�\�A�D�U)��zbk��5x�A�0>4]�J��h�oZ>7�B�l��8\A���#5�H�!���y�=�H��������0��B
�p��=h���O��M�s�d���k�.��W��tP���oG,�sڛ[�Ŭ�H_����"_A���a]��*�,�v�6�݀�b���% n#ҙ[C���f�geuClG�릭�]��]Qx-C��������n�R�ǰ�_ �Иp9{]mx`d��P}�4�h��yrq.�{�B��ۯ�œS�Ͷ`~w%���,޿��5aYv�S	����l��#m�r�WU� ֕N��6�'n��p��v�杔� ���.�kF�>n�Ё�]���έ�<�@�#�3�^��ԭ��<x���z�Pֳ�%�PZU��,��fΨ�e1�o�)`e���ܚ9Р4{jq�|R3h=m:�㿔�v)��R�({�k�=��G�Z)B�*�� mT�����ʂ����o�+�(�H��N�K�j�_�"�b7�3*�,1X���x�1͸�j���y�ѳ��u1SkY�(}	����1_���Q4�{�q4E���aW��Z(mk02ѕ�:� +�|�44X_��k�����;g'��ڤ�q.Z+��:)z}�	Y�����<B��5��h?TXh�2�hw��S��Ũ�A�1u�;zFP�X0ͤ�*�_�������5_���,V���Y-���Jm�i�͍P-���E���/)�其�|?�:���S����~���o���w98�(��J�h��r{G̠�B�|���+y��_���v���YZ���?�1��f+Q�:�/���`Jٯ���o���T���)�3�Vm�#��dK�S�},�C|��S��[�.�pdr1?��8�2�����ފ3�x @�RU_��r}s->~�	��A��˥t�E�]�;=x��0�����+�!�<L�}�l�z�A��**�Q�� ��W¶>�w�8��d�A���E*�)(AV4JOUXU�H���NB�J���(-(�wQ��u��U4[��H�h;:RWGU����hA���.2�U~ɩ?����GC�AD��0ux�u~~-(�>��`v��L�'���Za�O%Ջ�T�q�lci��M��c�X��ѩ\\�����x����c���"�K����Pq�֬�
L��o5,&��96�k��QƬ���)�eL����:X��@~V��� �������Κ�.��C�FP����#���N��F�:/���{6M��˛�;�.u|��>�&b՝�V@�d��(�^���/C�^�2J ��N�^'fpY+fx��`V���Y���z�����3�t��6�X�_w[��� ����g���O[�
zU�:�������3�M���\�&zmc�Q$ȹǘ�w,�0�j\�{ ftP��h��hb�A<֤��6�j5�+�S�W�lv�"�v�-h;S��o>��yS�+��6ж@;cf����#��Nk6:i���y��B���ˏo�<ۂvy+�~y'W����ջ<.��n8ޕ���vF �[�ƫ]R:X��� ީ�}�@��풮!o�R4���X�R�8.<�fwF[1�N���"�� �G{��̄�+�1�E��]�,�sm�� �� ;	O3U}�2D���dk��Ӹa��:Ef�p,��2	%��R ��~&�]R 4Uk���2:b�;�BTB]v�9z &$ԃ�Iק�e��&5��h�����*L���%��syvm��(��8)��z�hA�FU�އ��͹fƅ� 10pD�PU��
:� W'ӄ(̕S �]5��]�A��g��ܜ�ʐ��ذ}~��2�[�j��w���{�gX�"3p��>!?�9E�v�O�	 pA�v���2ޅ��������d�%��'�ڭk�ҽ�2����e�o�	Ϸ1�%�4v�&
<��Og�]A\�Ae���^}�­}�5�#��ʨ����|�q��w�M�q>0	�!yc2��0��=��=�oQ{Vӟ=A6��D�?~$��F~�ҟ��]���&�d��6߇���YLdp  Ӈ��v�G��(���u�u���_(�&��)�K$O�4	�^����7���2M��=BR���Z{����~�S��8��),�y*� �X�`L!����%��)���M��Mw�
� ������r�p/�?���c
Pa>�����;[�}�Ť�=�Y`5(�0����=Yu24R{uD����``LTP�7���q���?š�tS���_��a)�9qƍG%�WW��{�^�!;Q��츬�U�Qx���|�x�����2����! !�i�LL��%�.Ȕ�� �U�읿�I��e�+���GCj`�PΡs���J�6�dfl=�����5$)��OM�`��ˠ�7�h�L~�dw�d��SE����`�&+�{5�[��_L���z���q"x)��e<ųgDU�/Ƒ�Ѓ��Iݴ���AY��*#�d�7Ԑj���M���-x�9(�?7�%zSA�Fl�Xj[��TH�G�ـ�*5,�|�wg�y�]�����2{
yn�Z|m����i�� ޿���xp�6j�Y���OW��BW�\t��m�)��2���i&7~�T���v��D�W�M�)�����D̩5͎-�ˍ�	�8�%�<8+����}���/��=�R�#��-RPT6&/*�Z���X�O驤j�1��?=��� ��fc��m���[Ѐ����l�Y�U�.��3*f֦͐ndc#��6%�.6�ƶ3��-dH%6G��G���!J1�`��Т�6�/v��/.�_�})���+y�4�ky����������f���;"��2Y�6�|�����X�t���;V*�P3�`�6��lV�/�UFVgk� I�PvE�q���F0�!�4��fm�U�{���X�I�qZp��ԮU�"u*TE8�hU�Ђ�.;��(*��W�[&j Ņi�:��&
�p��=����y�(�sP��*�)�=�S���kR#s���^hp'��#:���m���Z���~�v�7��ߩ�gʚD�G&Ů�d4��5�8T�kE@��<z3�X7 T�Qp�Zb����R��Ip8ۛXܵ��I1��V㢵G�w�$�y/+o#�4g�6�ڵ�ǉ]	�ض �Y��`J_�֬���j�x��m(p/���~~����ꨡ�I��ix_�1�G*{��u�6���H���rm2��0�G���� ��"H\��U�
8��(t �����Q���i�v-��o�f_�~#�g%(�:������1��Z�N9�iC�4�m��l�kf�cr��`���Wryy#��޽鈠)S��PVq,��/��/�ɳ'����#���ruy������p��G uA��?����{�Q������{	�1�����^B<+j_6���%s
�h��u�3�<����x��Ko�m�{�AYS{�*+��ie�O�^e�8CD�����s��)(��Fc:0��8�%���l����z-<��YHQ�sq�}azФ̉h����t�
��=Xb�fB^~��߁�-�^ 
?N������ �3ק�ǃt�;�����
�d��9��t,��#����j�/~�o ]#��|-O�\�0E��>|d:�훷Lyà��\�]���.;B�GT�;9D�}��P�T�.I�Ft�~N���;��σhNe�
Gy>�P���0��G}\��J����<Њ}&�7M�ȥ��2�$�q!ݎ�Z�HVZR�*��M����Ni�z zw��L�O�j�Eɡ�2_Ȝ�j��t�8�YQa��a1o&݈��ǜ���3���Z9��}K�`UOe�p�״��.�V �z��-��!�GZ�a� ���>
�gM&�Iq�5|���@��퓼)�>Y�YzWU��T��X���Z��$�P��V?Q�'�V1�b�jj�_5��`�3u �&��v<E����ze���S�r[�:���<���]�Sv>�S�GG�������|<�2x���)H� u_�i�'�)�)��j3N��f��1Q4+lf���~E�4S���;"��_�X+j����}l�)j�FU�K���X�:
�+U���!Eu�1Y�;�޾@c�S���X^�-��B���%����5���}��˧�Ͽ{./�^�4����O�>?޽���[Z�[��)c�6��5��Ɋ� &��T�l��dw�Z����t$�%�b�t[��l�
�}���ʢz�����;�.`�72�����bI�y@�6"(Cn")L�gh���u��#lqR�V��e:U��h�y�KH��/���*g>�*@fW�X��5�@k���u�й��	0���(޵P��Y)H�w�ٕ�0V�B��Ck���Y�:X�:�P�MB$S��zM�'±�����b�s<��6�Lο΋��:$�j�r1�DUQ�2&�%��_�=I���iεR�C�2ڤ�Q�cÌ ~�,ԏb�P	�QS�CL�{�iM2	�Y����#��� �6�~Xn�ܮ�(�������T@���6Q[�De�}��Ii�LHU�b�:��R��sJ��Ң�Z�`�����4J�󇥼~�N���9>h�`���X��xxx"{{��7�*��%N��3�mp�������	����\����=3Y }�OVb:jٗ��8�b���|��sf���(4���i��7o�˟����������Q.��e�"X�Pk����*C[��bF`��3�����<��=�e���%~w��z��jU��t��h˿�7���y��"b���Ԃ����"���@0<�*�.k���y`�M��h�'˭�� ���9�kJȖ�^��r��|���zy��ڞBY��f�aB~;ȲA����
����O��ޛ�f^���������@O�v�M�·^Si����)Vl�����~��
#�j!�{}r�'o^��	TL����s�õg�
+<+���h�wU	��@�O�Y��F��W&����Q�2���>F��ep�r�lA%�z�%��	��BG6jC�h6�g8UI5�L�E'���.�	w�����z����7F���hJSWEݩ8�0��X0 �q�,��eݽ �WG9�Z�iX!@1��y��<wת�膵i���u�{��tTV��٪�Z3n��s�N�T�7���E4�C�kgC��8@��SAN�V^Q����k�qd�R.i���$ee~��D>{�ϣ~ѳ��PJ:m�`M��,�tpp�`�:?�RS� 'h�Y�)�F`���B�T���J	ߒ�{�d7%ま���{Y��Ab�:4�0C���
r$��U,��'���������"mM�%o��A6�nao�N��G[��ʨ����dE`Q�Mg�ɚe׵!�Q�8�u�i��U6��f9h#��rtD<��N��̈�P`-�;jh��~��|��y��\��Jn/����{���F֋;�a@�f�渉����'� ���Rg�$I�#ɍ�(����ۨ$J_�K\E�K����M��f)�5F-�^'��_e��Cd+0Q�gl3�|k�a�p�G#uv�D}O5�F�UY�y۝�Y1��Yf�D�J׻�[���!�̝.��b�mE4J��h5hU@)�F��jo�Oz���y�<d��UAЎC�2��Z��ӡ �u�m�+�Sz�'Zt c�6F�Kb�V�kY��q�34k�a�E�7�̪�G^�E�nNm�d��zq�T�wܻqM�7ɞ=����B��H؞�b.�Ń�AvKmچ�^˼Ů�U!�!p�{������~W���>�0�H�^cM���TEg��"TT���f+E����Sd��P��թ����J� �b���vVI۷P̯ڪQ�	�n�����Ǉ���\<�0�>���&=�fg�w��r�IU�5��	��@�ŵ{?9�ȳ__�2��6�T�&t��Y(cua��'���'/�?�=�,J.�� ���ݥ<~�XN�N�~���Y^g�%0l�½#覀����o��GA|���g�����?�9j�R�(�K�r�� +yǩ���O~�c�48_)����z�4C6.n
�Ok򔙄�tB�n!�Z.]b]ǹ����ZR��Tf��{g$�ϥ�����A�yKMYrq!k�m5ȚdR!�ߦ����B��@[�t�����6��hh�9y�%��We��9�����j�5���F���Z޽�`aGN�Ȟ\�4X'���`��\��ШJ�����s�,�!��L��~��EL[���__�跪O����$_��`����J�؍�e��~AJ��~�mD��8�sYkN�fT�I�S���p�pB���F�4�U��u�bd��O���p��R�2a�����M�m����ژ���.�Rwv�co�hT7��GFJ�[�(!���Z�`���h�8f��{�������௵�G��P�}����k�+:��%r��n뢆�3�}*A2[d�v������Hd`�ʜii�g`��7r4@�(�'}ts�{:uvcۙ!������5��W]��4��|TV��Oz�$����飪>�S~N��P"�-��/�s���F���=�ר*��$�5�ץTPT��x�9���{A!GtAYp��H�0�j��D�Pt��t��Sm�SWל,P筎v��~6Cl0ڂ�)m[aNV��V0�iІ��/3F�9;�|'G�`��W����G'hy-޾����jyG�.Z8��&2k�1��ͤ��h߫F��֠\�}��� GD,-��{�R@cc��Z�,��h`V����@a"���77��ǵ/�ѿ����`���2��C�u���R�am�֗�����A�T�'�<�|k��}ù��gQ��w BY?����ն'��^�iRO��z0eZ��  Sim�$�����@m�v!�&��-[���j�k�1ú��l����;�F�/P��P���% ��&��g�(ثN{|�Y�'b�k"���h>�.��;��fS����h#���l_�C^��b��fmG�?#;��`���|��@k�Jf�UJ��� G�c�v���u�@0�@���M��f<o�`%j?���Z�KE�}� ��*� �d�Eb6�bP��T�?�0�hL"IF�R���r(U��_%;l;�s�>	|(�I��Ù������#9:�ev�6}���h���o��D�O���j���<�u�7+ ��?��(��yyy-g�9`;��f�kE�;F���$�hw����-e�qz~.g�����#�)X'�����?��|��_���VEΠ�iP\�QW���:	�q���}��?/_��|�1(3�k�|�h��`���Z-�����ݲo��u��*�[�x}_c�ϜS�R�ݗ��5�h�F&t�qR(:0mv"��ִAY���w��Yk���E�O�R������.:���!C�|�1�|�l���I%��*�!K�P�AR�&R1�{s>Hkb�ϔ}7�]�����W9��xuI�M�vc�Ǌ � ��&��� �^���e޵�SzN�|�ygz���|���.�|�b�*?�ʇ#����% ���i�T�J�;o_�b��R֕8��� �d1K���3�dd��e�q�t��m��8�1^� ��LC(bΛ;���E��:d�]҄BZ0���ew���l<�2c		���l@2R� �s4�R�j���k̀���\3����%���&E���f�8�D�2��ӻl��E���ۅ��j���;i�i#�)ƲŐ�^u'��R���?�k˩��׽Bf�i���MP�;b0>�1�b#Nu�L��U��@ "�2��:W��p��&����gl����^�B�
n�ń]�Hq��![���F�����`��^|���V��$��U?Ӄ(�6�*�0c��tj3"AU������oI\Ҟ���>g�I:V%ހ\�k^쀃' I6�ύ�@3���}��҃2��:fQu�ƾ@���tn�������ؠ�&�j��P�����l0����۷�p�1_��NN��\g�5�, �Q3�Z�'��5��5.;��=�(2#-B����������\���I�&�/�mUdɏm�ã)�6+��p���=�7G����A�/�'���Ak�^��ؑ�a@��o6ىHZ���JkZ6T�ݰ�
T�`@��T�c��,9wa;�����<�#7 *�	���6�KM��K�J'0j��\�آw��R׵�r����r���@Rz���!X�gĶ�hc*w�TP�؂����z��=�3�uǄ���TD��_�cj���ϑ0�9
�5@�*w��Kt4��<�B�î��l
��f7�*y��'Kc�����{�:��˹
�C����*[Y����ze�u�at�X[����T�ZP�ŌY^�Ph���SQ		���F�S=m���m��S����u������S��g8�����m��@��N$���q�K�n�5�K*R��D��H#Y��F+��i˵�4�`b;�V;�T���6<�7o姟~���/d�?U��sF���U(�7��.�:�6
`u|�������T^��R���|�������1��f���덍O }Z���ҥ�bU%Ъ̆:�!�<�l�Tɛ6���T����EQ�S����̍���T<�ʅֆY�>H����
=x_�Ϫ�>�h�jo�SY�zgS��h-��A�<	ډ�*�*|vm!�8���Hy`�]֦����~��r����/��7ا�q���`e��G[�+1ʈ�� �b�'Q�k��=�z��'Ϟ�����r0�e�����>\���h.�o);�]C���]���T��u��e ����n�k�_+4ƍ\�x-�|AgX�i(\|Q�/jHk59���şQ��ԛ�9���4�S�����~�c��eY��F->�������y�Rz^@�()E/Xa���4�8C�a�;���A6�~���2���.�?m�'&� tq�7���B�yX��Zr"����١�d؛��f���R�i�ȟP���BT�T��cOvTJ�Ž��>�@R���4W3Q�ʇ�]E�0��ƮX#�;�0j�Ӆ�?f��D��իͽ�V�y�Bf�;T���k�� �ǲ{����� v@�Z�n ��/����RB�B%�W#��F��/us���\��������}���<�h%ڡ�y>D~lX`�&�x�(wwT�Ծ'-�~E�|]�������8�X�Y�������-���"UB�D�P|L�K/߉ڜ1T��E�.���D3�I|��*&GȔ5BIy
k�ڳ�!���.l���xf��G���t�`t��auۭ�+�����Ɵ+�R��
k�1�U4�F-#�x85���Z?��0�тp�®@��\Ds�H�1T]�\�X�c�%�5{�*S )���(�b��k˲'�3�D]�U�@k
Q��������ON���yt���v.W���������V�f�5�`D�,Ԥʒ�:�|G��|+�l5�6������l�����j�]K��I��Nw\�G�u��˞J�� �����I��a
DEQ�XJ%N�	��oQ�ʀ�O��_�*��}}��}�4 g��<v/jn��4z�;��۳�\��?@[��Ӂ�7���I�Z-�Z���\7�,6���ꕉ(l��1vJs�#�"���
Q�7�]��Bm�K�|�O`(z �^���9쑠�#[ p��@��j�����A��\/�u��e�z��o��g�����U|�B�h���ihs���i��R(��2B�V�e��x
�0t�U"����Ƃ
�΅W�h� 
���G�%8&
y`/��*`V][s�1_�����wS�Dٕ�Î,�>����~�kK4$^� �����J��"><��Tgң[UD6GM����h��� ��{x���K�̠a/��e^C�B!c*��km�0�G��i��iݍ��Y=h�`���8���֋�:�y�O��`;6*�ס%���Z��{j�geʌ�c ������,{@;F[�܅����2*��'u�wJ���Sf����,])EX���ٰ����s�Z��s�V���ѩ�� ��@�
��+�|�t���Ze�4ܟl�a-�9���ys�J���凷�e�T������W{����+T�k �R�3�?Q��7�5y��]�L���V��)r�����ӁJ�S��&B:����9��mʍ#*�5�vC����ߨ��R�8�;��Eʐ�7R�Y��D��%�R�hLEN$g�c��D�7���WX�gk�
Ui�RZU3��ң;Q#٥A���ifS:{�v�6)�L�������+����O���_�&2�Ytj �V�M��ȿj�������/^����7���R��H���>���C��ǟ���A�* �7�`��&�O�<���Z�=���6g�*u26R����c���P����fK9MC��˷��/��ɸ��ʣa��g�"J�@��%a��*-��lB��5e@��bB�M�,N�R�����`cZ��ƜT�5�r^H۰.ʅ�"F��Q�6\�l"�@V�9�������d�h)cI�:��*h\���!Q*ʑz&�sz������l�
q4S���V��3F`c!#kD� �ꆔw�ڞ�S��d>�0DK
�L���-�gxo��"�Bjs�d@��h�K�߸��G��1�S��-�,�㡀'���s�Mxﴮ�b al�VR#�LJl.���l!_e���vk�|-��`�Zֆ�� ����lnz�f�(�&�$�J}�G�1N�G�t�,&��#������F���:gRh�Zt����:}�����
�1~2rn�>��ɞ�̙S�4 gH��R��`TA%�x�����g������{������_���-���NS�Qa\7$�kx�KX7E�AEg�������*f��ܪ�W����MԈr�y�(:J��"�]�Z@sb�%��D�c� i�U_�b�h��O��o���{_�����c�o���$H*�ˋ�k��aoY�	m"?��B
e��gR�͛=3b���Z7}P/b��Ƞ�N���)��ք�t����Qe��%F	�T]ꎆ�u	qW�f���{y^tJ�4,�2=��m�����dBy=�
{X��|iJ��S��L�C6GP�!�{�eZ�]���9���5a�O�&�����r�R�V�&�	S�^��*<��� _я��z�V��v����+f#�F���Xeu&h)hV2/`|t�C�`b�M����E�?��E��;*�5�Q�����'���S���2�uH�Ba�0�gm��Uڢ"�&�+Tw�a��рm�าl`3Rڡ�Һ��C�X<��V�����#y��	���N�ү됵�짧���z�{�}�HI�#ZZB�(3A�<��w�R���c����z/���+���˼?쫸PrV��^�N�jAv�NF�V;Oq�J3������3���/e�B}�:�q\��ή'4 � +�[1cP h� ���^5H�����?�<����/w�$�R���/{s���b�x�,�+���]��}�UU�vA7�{C_ܕ��5�<Y%�<�ge�2kb�M+�����L��$D� ֚�����>�Jv\�	�E������V��N���X�7��e,l	�h��aP���f�i�J����:���~vf�<y,_��<}�7���T����8/���_�ʻw���#�0�T9`�P6�w_%���˳gO�4�FM	�0d4��=LR���i�_t�fʄ)�k�{�6p�u��/�B8t���l���(|���hCBJa"����tR�^�9CxZ��6z7 m���I۱�,È@��ݝ=��=��������$��E�Y���m�H�]�}���ޗ{���j�J�L���!���23^� 2�͑����d�4 pp0�Oo=��h���̲���S*S�JM,��r��H���`%C�p��z�����_6E�^k^�06F+�A�JF�z7C#���Z++S@��PW��ߨ��06��������p��wJ�Jg�E	�-��n�$��
�䷗�l�^�$�uM��h��a�恀�n��Y����.7Tt�c�����wJtAհ�"9�� ȕ	�������^�^���<������[�F�0���d���p�}Z�D�9���fGk˼�iB������s
���A��F�Y��u9��m;�g�OU���I?m!�f���6��F:e���i�rϴi�����LA.������U��&��)���Ճܤ�o�|�!Ԛ�y�,�e6�����U�4��:X��0n�P�y��av	���`��Ÿ�3;=d�@�	�2�U+Y���C��ބ�z��l٫�Ի�������zK��%&�~m��/w��������x���m&C�k][��	�h�������ۢ�����^rA��Z�R�7���}:�U��Ppߘ����hc|�׈�YF貅
[P�3�O�ô�u��F��!��*�������O���m8+i���]O� � 
� جa��ժ�&?T�0�]B��e��*�	J]��1х��J��1[\��	-��_���������0��{��6�_��b�}���M�6lҵ�^���`���}���0V:8׾:���C� j�*�)���ڳ�YRx�,�,�)0�Z�7]�u5�➪��l����ANHZ�~�U	���9P��	sW��������������l��Q�j�[V�j�����R̗���F�??��|�,B`�{�=C�;�
����dB�@m�&�Z��P�-�-��׾�y+����.�.}�F�&2_Lò=!D�>����h &�E��D����:����}���o9�ko:�?}��\^A�Xe�3U�0�O[�r���v%�����ښ"�W�Z.�����m͒��X�F7K��E�4`�Q<;v[�ߪ��W���Q�:Z�M�n��'�n#m3a�QfE��7#ScC�I��Н���`̔H����C�/�軵
�l�W+��.���B>�{̘����Z�[��-�-W�F�b(,2�fNOOd:Ջ='?��g���o��~x+���y���;>��߼�J �7߾���y���eP��'�p�|%wۭؿ�£+�;t7���g����ox��c���;�x� �T�� �&�prV���6;(4�*>?��qh������ ��Ʈ��� p�t��b����a[ Y����7�t����)�x�r�
�8{S�ц�&�����	䁿*){��y͠����� mc}v�ͬ��'"�
��μr��=yܱ{���!3p���2(P�����KG`��ls����c�D�M�\���V�,�s���>��s+[��Ҭ�ӿ!5�$�%�V�4X]Ov��Cĕ@p5N�<s8��Pd*���#G�+/�ć���['9��/�|��y��=O�(�Y�܀�כ���T�,�P3��U+���XƳ �?�q �{rr"_}���~�l
UNG� �U�}��fm�z���81�e�b&��Ǿ����nG��wj:kJ�8p �Q�	�
�`_uZ�B�j��*�B@����e:���V�wk|��Z�qtp�s^,�L�ړ&���5��T�a�@�&��B�����=A�>���^E�H�,�{�XR װ59|ۓYq�.�H���x4Jg�U��3d��7��:?��\�`٪�{�Wi�8{�����A�Ҟ��<�m�G0	0M�w���uhi����U�Y[�,��2R�A{��n��'6������iV���:DgoX������)�Z~Z��� ����ZA���ÏK��� �06��/Hv��kEfPlӣ��t��H���:dXiEم�FU*���)�=��_�����V�Bg2ծX�Z��.�pL�� ���M�J��tf@b���3�����g��:j#�H��<<$[�$a�{�2��-�&*$7��8�r���{�v���V ѩ�G�7�����������i�`m#1�Yl�_�*����h	/Ӂ;���)m.�U���Ypk����h��ȱC8�g�G���V.������h"�hP]խ��3�߼����y�����D)Z�e4���W5P
o�V����6�9Y��Z��b�``$+o�����Zno���"�n3�&�XB�������n��sp�H�5�ף#��C�ýقU�� ���LB��j���Ez�ƒ��V� )t(#�l�2D�ݽhתyҴ��^-��8��Ny�[��F!9����KLx>Փ����~��{Mh�
��XS�B�)m�$A]��9���}mw��U$�D�8.v�YB��Vז�oz��T�*����RV?t� ����8�A������@ ÍW!�:��S 0��l����������\^m_���I
���y}s�ޢg	��y�Bޤ���d&i�i���ĕ��[֏�[��ˉ
��' PW_�;�-t˿Y4u��_B3M�i��(�ؐ1fV���B��9���iḡ��YQ�W�A%�����5��z��9gLM�ɐj�e��r���m
���f�J�p�ʐ��G��� T��S����Y����ld�#�
Ƕ.�N��쀎ږ ��C�~k�����fzHHP.��X+�EAVC���8��H�����8Z�7t�P���7O�v뽏�� �UAIι���&���I���>�k��V]��A�����cL�h�(���5�	��!W�7�1�� ����l�� �%�K4�}k>ц{p�x_/;|��;1].lPb��oF�R�Д]C.3�A�ۦ�zC�
���4�Ξ'���*�\P�� evE���
���ܛi��2w��ټ#40�#
�u�`	l����<��[���k�P���h��ؤ}2J�2���Y
v#g��==�^����_�������E� >����&ʍ�<`}�|��ʞl#�"��dv�UjP����_����>�h�5Mp�egQ�n��2s���#@R࿺�X�&�����@��@�m۷����/EY��罻��|���_�Եk���ZT�����NA��qH���	��O�i�0;]��*�Ǵ���Ԯr�c�q5���ou��4{M__k�v����^y�� ݫ����ņ ��
V��cB��O��uׇA�X�A5��7)�߶��W��blZe
h��$�՗�XAݦ��
	$X0�r�j���=��.��H�m�P-��]�e��ؖ�?q^{	�����%b����9��oE�jK�c),ɓ�Z'�n-C��܀��։p��(�K+h�����㼳� @º �C09Mq�Ȅ��E���k6ߗE�_ϓ����g���/ .���r���r0@�ȩy�����NkU� �]2��~���ː� X�j�U���4��k\لu�@���I�h�5�qo� �L^�<c���Q�*�@�����1{h�����i�6�Rv�W�ZV��	d=P@����- �=\�ǎ\]ߧx4���C�/���|�����U
s�*f��4����|����*(ۗ�M�� ��0�N��r~q#>|���X˩�C�s��`�A�E;�b�Ĝ�C�D����k�]ͤ��R�s0��`�v?5v����Ox�+������񖅴�k��v�ǀ�ۼ�e.Ddw�ћMs`C���{	��*��Y�
Q��;6,��K�w4�S^Uf2�W���u�r#X��4�\��g'����y�/"�>JV�_x�Yb�:k%30��V���)�Y���,�#HH�կ��ϨC��Y��`��Xh���U�a��^���������߿P9EP<[�����~F��JVQ�RKe}ː���T0*��^��E�áS���u2Py��P����0[���4tm8ǤvT���yz�X�]��a�CP;���| L��ɡ�[����2A� jr����[4���G�{L��R�����K`��e���%A���0h̒SnC)!��%`�<]�J�)�%e����717���+Z��-��IS�$+�=(��A��M�
��@uO �j��ú5`u��fz��������K�$�f��eo3�bM�5�����q��P���`�~�!���5P�%�<{�1[����4��.����"�n��cӓy�6�}��)>Q��+�X@D���q�+f�1� ��`��&�95��f���{��뮰$H[tU�n+VtT�Vj(e��:*�`������T�*�j5+0�],0�{�i�����Lx<;}&o^}%�NNe<?f�5�,�KS�*��b��h8�`�S�`c@+N{�Yڳ�^�^|��?|'�/�Y�ޤ`�44�c�Bи������$�H���܊e�_T�X+��A����7*����$ �+'��{�/�jje�M)��g�52D�z洶`C~�`�|�������Q)Ю�T"�b�����ׁ��5֨�# t��0hm���������c� T�m-e
����G��{4!hR�6j��r�p���>���s�H�@G2��8f5-�;
B��rMB:z:��W6�9CtѦg�$���0зym��t�k��:pY{~5���4;�3C2=�Y�����ĝL����}(��j����]�
����sh��� ������Ǿ��"A"��H~�a%�//h�'�	�e����V��ҡ:5�F&�~���о�:�=F%��se�d��b�Ab(|�D�Y�׵��k/��қ���Ɔ(����Ÿ�j�w��ye��PZ�W@���EJc(C����jA�g�\q-0�*]���p����N�{���
�)ݚ��@Xcc�H�,\���:����cBR�~����	�.d���lq�y�KX��z��` H�ֵ�Mfr|�,ž2F���GJ�$	�0޳4d�x�����8���1e�6�bc��#�2@E`�l]��/ڣ��`��R����]��Ly"���kN��f�v���ȉ[�<�l�����v�	�ĜX�\J�.�>��=��sN������1m<�"AAV.��;�ג�"���.2�l����]Qm�0g;�  ��IDAT֬�q���gY��B��	QB�폠�+�������� @�E�)z��@��ဩz�0/�a���?�ի�����|���ΝhH�x�Fp�z��W�Ě�"�*� �|}Y1����t�7#�Z�=,���2��	�0��z�˨��(�ޱ���5N^��L������s�Fxf��	V��p�YU:�2�T@�,qS�����V*!��=��$����h��M���7���ȟ��A�L@f�.����* ¦�%8�)�Y6[�0�����/l�{�K�k"�2B�:���>�-��ł�E2��;{ܲ���+(��3 wiU�Dg	��ʻ���=*g\��Gv�n�� }G),�d�����9`�!˼��u�[�N2��,r�Zс��P�J���-*LzX�۝��S�z[&����li}��d�kf��X����=z�r�;ZE���(�Wa`��`A7�y�t�GX�r��.�H�h����CPP5{[ƣJf�����R�6a��l:��g����7	`����q`�2��{;��ŵ�����ll9�% Ҡ�j����s'��p����8o���|>�$��eA�fu�Wv$y^!O�=I�j�����v�������ԖU�U
f6�{���1Ir�kŜ,T�W���?�ס���R���t�r�g��\�@����J���	� ���8���6�P�Q��چ��H��#�J�G6��
{��X��[��F��v��Q�S/ei2���2�����PV�_E#��
?������|M����V��
e�}|
�Y����f�Y9 �p�Bڦ��
U���*ɶV��"Q��hR/��
+��87�-D����&�(�a�(���m��^r���-�%�\�U���.to���+�}�$_�TqM+�w���	�L�����J^�|-�7�i]h�@���g�����V�����Gc����R�sCl��|N���>t@5�A��I����*[1�l���N�EYB��}:�W� �EѺ��.Jოծk�Z/5�7:��9��u7U$�b������z�`w=�6j?'��r����R��,�N��Y�TM�RD�^�A�ko4�鞂5�`�,֜Av�����F&�%�~�W�C�
;�?��Cdy��>9>�ׯ^����k��MO�����Ϝ͸�lP��3sy�~��e�$D�����7���]�
x��S��Ws�Y��� .��Ο]qY�k80+��J���~أ;�-�-��}��,��QC�����mKѰcwQ:p�j�W��,�I���N\G��%���ز�-J����v~-���_��e�o.En�.��W8m&�*��F]�k�,6�Ã�P]jQ�?9�j�G# ��ff�ZY���x�G��� 7;�:�{��xj�� �{�w;�E��rY4��~��,$�Z�+�dUV�2�Zz��T�ʏ[��i����퍜_\0��7�]f,�9g�&@�oI�j�{�n��4
�	���cP�N�oUa���.��Q�k�U���#*��-xj�k~��=����@�x6<�emg:4��q8!�)�=�\aC��7�ږ����te� ���o�6�%o����W��_���9���.�1��5X`5kC@�Ȫ�Ȓ=��,��x�����:��@x���_Ԃ�
R]�h>� �&��@r�#�f�M6Ё�Y�����-��|wܻ���g@
*���{��4�m��6����I���d�6���������s(H�h3���D#��?E<Զ������%}-9幇!�dÂe�|�w��b��E0 �]'P�BU�cH�C�x:���T�Gr|8g2���H���k���W��8�*&�	i|�3��Ym�{!�h����Q
�L���a�s)��S����D.�9?|/�?�"7��L`b�>�5�2ЛS�wl��X`�gO�����������Wӡ� U�,4aa�M�=�*�kx'���<^�OU���]�wa�Qf!�� �ҵ�����+�"ڨ��u��ZU3�N�3�����#M��}B"ɃxS�|xXe9wo���{�
EU�
=�H%?bg��8�Eq�2�Ҙ�"�*bQ�+VJ�U3AR`�&���a��V�%��\��N6��o��	\�8~T $�u��(� NOA���4����Z��U;T:!�bb�Ym�}�Z1���68 �3Z%��W^�_�U�k�u���
�E���B��zݰ
�0"�v,�i߼y��h
�߽�Y>~�H��|~ /��������A����?���& -�혁:$���8���-���p�ڡ���P��T[��K�����=�o��BQx/�oYo[@�� ��mNP��S
)�c��ĝ��4��Y ��h7�-�5����c��1.m%��1���kO�I��Ym�Qy���_)ް���ّ�~��3O�����t��O��O�Q�n��|i��o��-?;�G�z�c�J����\a��h�[�G�_�<�k���0zߗ&T�E�Nh.G�j����T���K��=s��쒃�1)-�A���e�V����~C�l�S�:*��6
��$�8��>s��{S���^�S��:����N�-�|����b!��'�P�e��փB��y�<(5I.�Sz�����g�{�|"��!�*V��XX)Ua�@��T��т#x*s6��j`
ٿ;U)���P/Vz��J�">lq�d���:�r#��������5�o^����XG��99`��w� ��U�\��a���Rڒ6�nH�Z.+��,���K���������X�uo6
^
�`M0��݇	�qf�c֙m�R���,T�F��,��5�BUPe���k:s8V4ImE�T��`ǥ��U��ϫ�A�����L"(Md6[�d2O����<t�������q�	�+RY�AKP� }Oe�U5λ���������&j�3�ȵ�ȝ��Xy"���j�ٛf�9q�vIU2��E�* ��틠��
��9���n�0�G��l�U
�tfJS��{m@I�@𧊃��G�C_�D�_�z�c!�UX���=ӡݏh"9�`@�fc뢱�s��*��Ф���������a
n�YD���B%vI�`m�n��e�����d��1��j��3�3�"�����@��4q�����w�@}�%fs$G�7*e>ۣ0���$�z��u
^1K~z�,��q��8>�*b��I��je�"���3R�p 4[[�\�*�qpx*��\	��ȧ�L��4��A�>��4�4Ʋ��^^�x�>��^��l@Þ�;�N�7N{z���L���d�IELSs9����꞊U����df���=ˇ{�->��ûD�"�w7|�� im��Ҁ���=����ڒ
�rؔ�t�5��A7�U�^�*)�<�L�=�S�?S*��l@i��֨5��D¥)��I��zP�-�&d�-�#�'H_֨M�M�OQ�H(�5�?�:۔5+f��P��@���`���2��F��Q�*ad��ײ��9�T�,٬�>�4�_AE���Lz7��̊q�Oa/a�1�d�GI?	`�����9�7��>U�7#�3X"�͠��z��-��Go^Ŋz�1V�8�]���tA�v||*/^�b|�
����\YgYmVlF����m����� G��z��zpi���GKEn"�/m��-��a"�Q/���t.���}li{T��[E��~�
z�c�!��|q���CZO{2�
)t�>+p9?��=wUT��t6 �Ҩ�0�i�U���f}��7��_�*����Q�W���R����H��O�h���eO��e���t���d�Uڰ�����b�7��.�m�i?%@xŤ����ޒ�O.�s��ً%/��-aO�{�!�?�"�M�wE��{�I~�c����ˌ�(|/�N��\9��m�͐�&DB��+Pl,F��#A����o-��Zb`/��0������O�J���g��������;�%��M�����e7������^%f��8!z/��4Ry$�ʌ"�v�Pq�0��/�Q{�_V4�B��M���N(���s�`�,\�0#�A?A��sH�kE�=aE�	���~��?v����K�_{翳��}��_eX;�_2��Vy�������K)�e��>\Q�5d��` J�ʂ�fv�?�X7ɰc�ht�_�le#*ZY��P��k��ͨu��e'H٨���l�Pp�i�A�&���)[�M��V6T�%]p���4��e8
Z��e�l�XrR���}fc1�o�j��P�L0d���l�Ӭr���W0���kk͠�:v�jX^r�$��au�2v̩)=����� (߾b�.PVc c���2�.� � >�)x���/���rPa��\���q�V� r��Q�(u��tF���4�����&��ݥ�����LԂAs0EH{u�spPK��d��3ߜk(ee�i���t��|��IΟ��I(GGG��CՒ�o��l�(ݔ�F1��������%�U�?�z�� ��~ѐ��G��^�B��0���*K�	�����&8���ԬG��E��TD�BD�^8�APrP%���퍊��1g]&.���@zĉ�*l=�R=2�=Ҵ�4)�}��-*J��������=����e����ǻ���|��J�f*{똝&�4��u]�ؼ��
��聋��������c�����ʃyVWǄ�Z�,9��7r��\\�S�ll@�A���+Y%�uɵ�I#�a<��Mm��m�m1�t�ly���&4�88�	D�:��봘�S�d���|�`ŃtX��F�{�W�`����`2���2����xoC0��dW��?�bbLBޒr���1��&�{���� OnkK� 4!��׶a��*�H��13'Kq*.�n$xK�
����,:g�m6:�ͨ���v�U��`��L �����6ʪ�!@+���}1{&��]j�.� ��M�]�'���|(��cO`��(��|��� ]+��^�����/im]��	!�F��IW��`�* ��8�{�L���f���XX�*H�#. x~��h״0?H�o}� ^������ W��$�V%�?~<O@�LF'2O�6�=��{{�ɲ[
�l�$Ě®'�a��M�f$~A�/ӵ<H ��ׯ��������k��%S�'d���/���_H��6�ۖ:D��a����;����Xń���ɼMǋ���lУ���fت�%<I�I����z���б_��y�A�=���7C/h�kbw�dn��-���������E�Pn�V��D������G"	�A�ҽV��#W��w���n�@_W@����N��X(t�׻d��7��-�d�z��>舽���^>H{�n��:�>��իB�*��\�4��P�{�^� l��na�η�6EI�s���Q�2T^�>�0���L6����y6	pdo��a?%���=h���K�ǵ���bѨ�-3�6��t�΋h8�F�&yk�N}�7�ݱ���#Wiu_�mH��ap]��֣M���e1u�6���D���-EP:��qԀ!0���v���"9�v%7)�A_�����p�臊C�U�`C�EL�M�f�#���זr��ʎy
U2U&dVah�L��'�D5ۦ5<ܛucC!���I���0Zsh$��Iy�J׮�,�,�(�x�g 0̣3fէ)�@@ւ��/2���/7r�eqK�EE�h�Fl���A��*�L�P+-@+LV�p@Sٵ*}Wr*�ӟ�23	0�e����L�Vnu~��MR~�]��R�句\}:wV��6W�B��	�KdjA�SZ����Өj1\���o������ýH@k3����`̬3�*T�B�-L�BJ�I���`��5����h�Ii5j��y�Οg��\c�цX�>�A��QYq�u�a0��W�T�[��Bkj��-#��M6�ϋ�gr����. |�hv��a�}VX��7tW
EhU�kJP
P�J��*e�4Ke�� �D�%�g�!O���0�n��Y�
�e�#Q����p(��R��˫�����Kyqv��۰��e���'�d$�J:g��N��W�@��WP)J��' *]�לO�p0M�3]_T�'��� ��k�@����b'�e�A���I |
{ M���
�-�82�鉷��� m��<]�Iz�Jc���=�>���6��o8�F{.!����P%N�M�U:��}s+6�Ͳ�*���SP��T@Dձ��o?����~�ϟ~�%�X�~�A��=� $�RB9�6��V�Wi��cP��H�K��'�"������n($:������|#�'�rz�jl�\��y]�d'�
�k4{�u�y�H�ao@�c��c��e���q%��{�$�-U1�=��t̓j$K�AIv
[>�2 Iأ� �d$�����K�؀� ٛ�Q�~�H8��]J;G�!����EB
3 �k��འ�"�IX�X�ZXЯ�sJ�%CVD٦�&;0��l��%k䐸4_��[��Ƚ4���*�N�v��S�4��t}߾�A�xz,�_�fe�eQ�Gǌ� �|�#��������!�@x���S�x/��{y��[�I�s%�t��qf��S��A1�n�q��L��S����R�Ih�ЙK���9Q�U�*.T�����
�i3�8p��r�k6�kOD����� P�ɷm�'�!��~�pW�O?�����e�?��ᔬ``�2��Qؓ�=�6�p�1��
W�H�_�y���]���r:ɳ��<{V��*��bD[���������Abr�l�Hl(dq!�V�^��<��/�~C�O��1��t-���RnR�%;L�� Y��Ze��4W�g��F{#��]V���'ep�ǧQ�?�	�^����_��Iiɿ��u�#b�mZ�(��-�2|Hk�V���Y�ՆVb $Tur���:=����1�h��,�A(*cu�-�1��.a�d��||��%�\?�!xT�p��x�^roc��}��
�w$~i������0�¥������_�������?~�`I��7�,��jfJ��E�ߡ�kc��td'���l�?� �.>����q�˴����XLg�?X��ב��U&��Y
.8�G�Y��w�m/��fV��V��8#�[����(kߥ$��l�7A?�J~�e�<t����E���z��Eŵn),o ph�F��6-b��!@�U�br�-����q Sz�6g�97p�+m�GZ(�l-%��C��J��Pb%�o�܂�1�l�.S� _�0�ʎ�wX앿��m�y1�+p���cc^�������\{�q�!�k,^��g�T&	�Ι�L�2{?��7a�G��$�~��U�b��ok�Yt.�,�_�k�*�1�
�:�����a���fJPv�m�[�z��::��R�'���*��=�{�t��RZ���};:jp����&�ܴ=Ye����T:2�Bo�^��J|G�F��"��xú	`X���T����6���UG��M:�OGQXu��S�]�����aݏ5d����*9�)e��Y
�_�|��3�<VVk�OK�P��M���Nf�����>�sp�	ހ��l�0]��]��gޤ d���@�/���ad{]�ȡ���>���$�v���r�I��	�`�����'�|��]�ac���)L���lff�~M#v��7�+���W��?f����9����������(�0�ǌ9��lT���m)��aPY7���Z��t;�U�8	g� ��JE��r��o~�/)�{#�����><P�1$u�Z���g��``w����� �߱f��'	8���Ꮃ��?�����������胎��@���*�|N���V��{�����F�H�l5������S)~eA$�0zy�*�00c[ߞHf�]�:�}8�$j'�}mMm�w5�<.��Ym/�U?�UӠ����D��^I���8�-i�j7)�$���_�˿��������R���#�G��K��vA�s��&S{/��������O��V<����AmV�j��]�U��8&���)�mG�V���Rp��D�~�6z2͚"�6��xRp�ԾdO4�@`��\W���@y�K�z��Y>2b;%v��A��B�	����0!��j461a-��RY؇������%�J��<����{	D��-�艅VRa�� ������D�Ξ�x�0}�(K�y�����}NZ$ip!S��O�]ؙ�IK�8p��'U��b��{�S/�?�ζ�w���h�\����r͡���*$7���T�9��A���F��󴾗L(ʹf����<ж�R�Wɠ���*����<�K���z.^$�bw�]}���Pޯ?_���I�쫒���C��7�=VQ�|�7h��;.��+W�Ħ�A��-����}���ۿ�����g6y��PNFs�zk�ڟ/����3� �p|<��l�3����
��6� =�����w�C+[�0w./����+�e�?ǏA��:}u*Q/ �	�1g�-����{d�6�-�z�L���jY�5�z�� ��\��Cz��%���J��o��˰��(=fÀ��
X�1�V 6��A�S�?FQ�+$)���.�͈A ֆS�bm^i)�X&	`c�"��?8H |Az�`4c���TάfCuA���歩r[�"a�����X�,>d���v��p��n_�}�߬]��I��mg�.�x�mp��i^k���c�YA� 1����WJ#{բ	.�����]#R�hjtj������Kh<q��q�z�֝C�n��H^�EV8��տN�A�U���oe�� 5���r�$�Q���N	P1��(寓��d�1l�m��c���q�-`sz�R�t~Ma".��D�xx�/Y��x G�xr ϟ�����W߰���D&��0�m���F�(�},zB&�j�G�{�u�Ԋ5�᫝���3~�3+#̟�bb+�ŕ
 `���@�F���T������1��o�N؎(R�Ԛ��L`C�a�ڈI7�eɫ�4�,C�;��f�CKKL���}��m�����j@E�cT�����W �ߥ �/�˻�Lp��1�8���c�R�P����k$����ث��l4���JI[��.���b.�Gg����r���<���$�8�a���%^p_X�Ya�ɑ�.X���`*�qm�!�Cq������(��~��	�nH1L7H�u�-�>��hP�]U*G�� ��!#��*� ����!���C����HCl�%8���%_�_kY��Yb�Kӷ)�si@�Q��u���MW}����ױ1e�s�TPaca�Vb�*lJ~Q������*Ʀ���){� ��Q*��ϰ�W�&$�I}T	{�~j{_$�M��	y�{�=�T�qu|�]*�2�kR���]�>Ԧ��,A?璕���V5S��k�,��J5�d�Q闔B��s��>��?��W	���^����j�2�q����E/ȔTа�d��p m��KPR�FA;����=�8�:]�;Y/ӽ��&�S\Rʳ�C���[M�r��D.��:�#ꩨl�Fr���Y���)��'�Yx}oo�ryy���zC��m]�@����v�퓆��������ig�o�c<T��� ��0N˦g����T.���[mB_G���'U�Vj�@�!����N��t?�9;WjD��w��=�ޏ�z~=S`=nȉ�.����+�@+���_��?��_/�j��c�&���ǿ���ӌm��?��4a��Vp:���g���f��X��jpԯ�.�Ç���O?�O�h2��/T�`������}�Y�oE�A����A�M�}�/R������h�+� �/��9���@<�k��ع�;�Wp�`=�,]�i�fi㡛Ѕ�����X��Y�Ԯ%�t`��ʃ\��^S݇�vF���S�[�d)�i�9�����j�������H�bQb�����X��*�Zo�oVJ�b�*����+�dܐ����J?p�A5����X���=�3�<�`*\� �N��!j�=gw�t���ؽ��n���;{�h;�U��Eڝ����p�s�Vm+4�g�g�:b��U�ld<�؏�F#zr���f������~L��@^a� ˨]�.g�$��Rnu�E���D��)j�"(�K�5ٺ}R� '��82�=p���b ���zq th���5u��d��}��tol�(F�2�=F����HΎ���������R��ͷ�����2P-Q\��̀?��)�F���X���	o���SR�����0Ԛ��2�X���P�&�K&	���p5�\]��@r!���Y�u�:�o�`���E
�&	�u|C�{#����]LhFzs���zɷ�	]������J;j�F��s�9�k�x�V������~��\~�(�ɀ!��������t�(�T�K�5nAoӵ��3\=wP����q
 �J �w��7�c%soz��U�p��nJq�EM�y �ō���C��NfU峖�l���A:�}
]��S`��U��յ� ��Gk�/����`OA�~��WRݴ��(���U�B�'pX�lz� �+r��U�ւc͸�����B�=�nt�>:P��V�k����!VU��!A3�}�m��2+H�Q�t�	�;�CV����9�i��� Y�_�}/�B�\��=;��/_�UR�"m*���7N@�2ݏK��:���e��90��4�s
�~R	�f�JmL��1����SAi�6O��/u��'�����A �ʩX�l�(;�V{���6Ғq�zPAF|�x���` �t0�)7A��|sQ�5B��`�D��[���'y��'�|~/�aA�+�Az���D������r{��:@V �Ƌ^�)��� �ku�h�7�Ky��|��O)�=O�y��{ѕ\���mǘ�Σ����=���7�k�����l�DK(�Ʃ��~"�~ʍW�TY�e5���j��sYP���
PׄoE�|f�������e)�;d�	]����]�2'g�ة�w_�����Q�%W�������3��c��o�j�-��s����td�je��ق�f�VNK�W�M ��Zs6@k
y

�)���۰�����-'8�X������[ըzv��1���XI1�܄6�{7$#}���������C�!�-�n��f�#4S&y������,�ڂ�b,ՓF#�afM�5[i�t���2Y}�9��vZ��T"��l�AW�p�5�Q�8L�_��ɝ[�M�� ӿI��Z����]FV�oT��t��ѐ���xdC]���T�.�����!�A�����rzrJ�%m�VJ!zCpȮm76��ե>�s���x��e�������ri��p�?����n;�����閃��`���(�;Z���g� j��[KF��3�YĨ�=�-��Err��^�>��̓�rz��J�SsE�K�f�bW�$�?-�G�����=��+xU*�4�����b���Bu�6'RY��8�Xz��A_�#"C�}��;�:�6F{u��w���r�ɞ���p��@֡|������o����l��C�5o���y��S�
��i�+{
8��������`�I45GS'����F2Dб7��؀O
<�KP[�$��(���*��7�����S�c�E��dts�^� @�Z��?,O8,�9|v�
�'����@da��\�����N�{�hs0�*_b��������������w�)�X	��G������Gx=�2M��O����J5m��ȴ�G�����7��W��I`�ҵVIUE�룆��^<6���C06�X��+�6r��0+�X��	��9M 3�.�����?�5��Z�m���1T�0���B��A{-'P�j̈́=P�Rh��t��#���SD�����l��ܿ���P�u)vw�*�^j
��M��8(g\*U���Ҿ"�b��w�qFSqE5c��*DuZ۵&oZS�-=	���~�Lg��������V^�z��� *"��Yz2���y/^��w�ϺQ��׭�����������O�?�`n�8-r�j�d��������!�!v�/^39i�����%y������E�����}m�� ��Z����{2M��{D��]˕�(��RtC���BL"Qi�(�5`=�}�	0��yys/o�}����N�����4^��T��ʳ�D��Sy��9��ARIm�J�PP�GU��	g���������O��Y����߾K��صp�O��؏P�x�K�,���c�^�c�G���}Q?���Ś�ﷺ�cf�t�#'lۀ�&uߵ��J]�d����*��:W�5���>z����Ѝ�w�+�L��k����
��B�3]앟'YBI�Ȕ_;�u�Sp��JV����'nA���}p��U�`�$�CZ�ZZV�T� ����C������邃qQ�Z�6jض�d
j��h��OĂKΥ�5��I�(37[��4�����黶�k���9�����c��s%.a��-��Y?5��Q���˰Ri�RE�y[6�Q�X�
�n,f����g*����s��H�gR��j��?>�~8��3�.�J5��L�3���^T�3���ppP/�/0�.B:[�(�D�CC���Yr8/^Qn2��� ������}��P�Z=��BP{D�k�9�Ei���[S����
���;��˵��{XvV_��Ֆׇd �F!Ň�X��k�U;1@����[��k�2V=���=��돾��fRȣ��r~/'����%�5cYXC�m�v�[XJS[s�������)`��(Vr�J��@?��z���!W|,{��l�_
VF��i
��:T���Wa@�����v�ũJ~��Z������uȰJ��51� l,fAtc$���#9����p.�ΞɛW����iO�Su��j ��
?��(q��?[�ޟ����3τ+}NT�EH���j4a�	�A�����x����l��U���m�[�niY=���2��[������[9:~��h#�܃:�H���ҿ��E@[�J��������+Y��;�|:�c�lfd����F>~x+���.����\|x�
�|1eЉ�^�����
� pqoӞ��Ao���n�|��[(a���\$`�;����������J�w�&
��ws��4�b��hvN�"Ƨ�}e=(���NTM�����e����� x)𠯣�f'l!�� j��ud���D�|@{��.y�[��T� q�؃~v帶S���C��I���zT�HQ	`*�%��V���B Z�*Y�|u�jSQ��2I��S=4�Ǿ��P�8=y&_%�q�˫K�x���_
p�hS����/���� ~���C���O>�/	hm�*0���w�'넒ԥW7K��bUʈ���,I�,.T�}@l���H:'���?��H�����$�'��C4�y�:�P�e`@6@�֥�1p]�M��``�&<@�j�	(���dDv����������B{�t�v�	!��P1*􂏦��Y���O����)>]��}9~~ �H��	�&K5%���j�6n�tMn�-C.���ڥ��>\˻w���� �/�Q~yNp�Ĵ��3���v�[i�8�	k��F���濳M0���NV���z�se[����ŷ*��ű�ν}��Ei����<9[�5>�v��fg�P�t��c{�&��$��x��?��|2͠��&h�O�+'�������IVݝ�+ ��0<���WY�6}b /*-�� �Q
n���T�'J3n6���Ѽ�AdhQ�.�@.>_r�o� ��"1�[����+�i��s�]�}�f�8����s�_�N��o�c���r�:�c�z_ȑF�*r�+h IC���g�{�LY���$C!�%���Κ��aS�q�H�Q�ޓ��XƸ'	`A
V�j�.<��I�f��LVUN����~�!�`�퐒笖�֣�ѡ�u��*W��Q��}V�J�b4����Gx_�{T*+��v�@7��ӱ�YrL'	`�f1�|�QZ#�@5.�HW+��"�*�(Ϲ,�=�B3)XW��Sb�tO�v���p<y�x0]݌��� ��z�0%g�}3��8	%��8�����F��(�*K�/����ht��-��RBh��޾��E4~���q�.Lj����׿:��d���8��"^1,��X�1{%_��vC۽�Ww��_G]�u7��{$yN�$=����ņ$*�o;��2A����f�c�����\��)Y�ȼxpz��v͘�e�F���?ޟ`=;ܗӣCʴO'sV�����^�%�4��A������[/�l���
}y�ݺ����]��~ǿ'�3�d:?��������gR-�d�l��#���kr��?ո���W���!�)�wuIH���t�>�i R�N����@U�ڋYZY�S&�m)�ly}O��Њ�yZ��/k��]��Ͽ�۷����9���o�mN�{1�;��zf�>�� �k0T��41�4o��Ì'{9ړ�遜���o����z��,Nv�KO�v�D����i���_v�s�r��t߃�&� f�QG�O��p�����Iߡ���.i�F�1�j��l�A��L�m�,7��(�*x��7��P�;Q�/JJ���h�Z8�t���`X!P�u\ZϱQ��B+WRԶ���h���K�L�0f1}��������=I��$Q%���H ���Y�~��>�6���G���� �9==�������'0����P�U�YAZ��6r�~���2�R'��G��k��
�8�{*>�O��@�
F�1i�ib��.�B�ˀ�Q0Pa-��}�	��mЇ��Vz�զMǁ~�U
Γ=��=3��R���ώ�RL�S:�[
Ec`D��ݯ)���u�M�?)��@��Ճ����'��~����|����Ͽ�����\
<]� F�<:.�s����=��u^ob:�%�I���w�����|��O���gY����@��y����t�۾}�w�Ξ����׶�a����A�I&����Pş�.Ac5������u��`��q>�K�������mvz�+�O�>[*�UR|;Vl}$A�;�X �@�.H��J�����T��cw����t�_�������G�������1)���� BEV�*b�X���/TaP*č���j�����K�K�qz��D�F��R�Z+3�L��v��@B|vF��S���_aI��v�?�n����?/.[�zA�xN�巟���9�JjV(e�f#�� 5Adk�-%7C;�� �k=�M��&pU��m��Ш@���~^Ja��Z0#x�U�ʿ�X�ZЩ��>Z��$��,lL(�B2��e&y�	?%�[5����BY�p����,9(�$��ԁ ˅@ �r����͙C��ǐz/!�ZZoX`eP)������x.|�߀ hhe�(�q@,���77i;��]������=)9L�)<H��~Z���m��\�=h ]!3WE}yڻ�{�Ýɥ�E�k�[�iD��|�0�K��]������D�=[��a�
�W���sn�*�{Rt�0]����7Z���j�J ~��<�<��#�/�5��)YdѢۀ�K��1J��|�n��-���[��!�<Nu���j���ud���syyz$���p�*[at&�XػF��/�(�Z�$ǝ�{,�r�~'C�7�����/X:��b��d�^��y��/�/)�͊lP X�`A�a&;�}�V4�&��2լdu_�5�6�Y�� ˣ��2�7��z��2`΂bŽe=�:1e� $�М�`�g��� ����Ƿ������b���H�У6Q{�����>3ۇ=�*dU�ꋸ.@�N�{�0�/�^��AC���5��;�6��#�^������P@����3�aL�Mc�)�YD�R&�HA�Y�:�u����չ /�*�1�	މZIB��|R��`L*$|�U
��ݠ�aطӔ���SQu;�)��v�\��~4���`���Q�;�A�m4�'�R1��rU��sذN��m	T��Pz��W�{.Xό�͵䪹��ZnU�d�y>֛I�h�8G���zOK�Z=W� U!X�u��1m'>� �b����s�����j����^��ׂV�)��2(���m6'����:Q@����1��	t�~�VhH�@�s��A5Ik @𿨒����<���s���8=��ްZU[�&D����"� �hj󹎍I�wu���_~�?�i���fi��J�^�U��}��A�9�P��Pf�bZ��R?ܭ���A�?]ʟ��CX���?�,矯��`U�����,ԮH=���?��Ԏ�~�z���;�e�D �}�U�����ь��q��Ե�ͪsߕ�M��ɞ�+�N���9�l3Ű��b��bp3��&����M����[�OW��Ų�v�B�s��
;��\g��,4��_�`��~������D(�+/��r�ņ�ֵ5�+寵���df�i���<P}����W��%����J`��8w�v��_;��nB���'���d��JY��øN��1UG5#�'�^�_�f��8-i���X��e`
�t���&�9S�<Iߡ������4Q�EC��~Sgi�r�ԀƤ��.P�� ą����+Z��5}�5�7�;�@�i&���cۋS8V�ڡ��5|-�HZ�a��9��l��b%>��UBB�q�pO��#��Cn��� �e�,Ѽ��~6M��o��(W��WB=��	a���t�-v�����9���N�A7?�&(�� �_E�4�GU�d����7@��� ��FAQ����@U�ϭ�����w���~Myl��7�4��"�N�!ڞu��M��	F���;�i��m&E�ϋ�gV�����R�P@7}��x�B����?�SP�TO����~�M�����>�Q���sõD��R��+���!��`
F��d>$'.�����/ |rD��3}4~��/t,�f��Pz�l��U0'���}a��{X���Φ�z,�~[Za؛ͩt�M����&�K����N�O�/�)��X�ڢS3-Xh�Ry��X��g�a`.��ᖠ!�d�7�,��8��~8od���ٕe�xgcv�ӹ�0��{�g�-�_���ӧwrq�.�|�lփ�A��p���R�%���eh����
�����K�&��Pi�G�r|�R^�|#/_#�g�\�L�\E70
#S4�����|��}������h�����F��#���$3�;� �Yy/�.��5R�T�o �A�9�0��1s�`1��nRЅj���)H6�iL:<�2%@�=N�-,+��JTI�|sXy�� T���Y���9���ƀ�Is��1T�+�'��F���',q�*�
AնW\�`��b���QR�L�<���N��QHZ#F�<*f�j���X����ʀz�hɲ��:�Q �(ɚF/|D�@���쯆G�S�����Re�>��@�8X!Cx��t:{ ����#P�����  D5U+�|��\���G�v1��ysR1�����J���	��X�dC�t�c�ǈI��}��9pK���3O�b@� Y���#�H#<9>$�f2�iG �uuq#�?��w�?����/o���g&���1,�o�i{�Yܿ�3�O}��G���^����邽�U��u�~+���8ɫ�1�5�+�J�M3�8��N�������Ul66o�U&Π�VQeP�������9.u� {�b���}����.�g��3&�DM���,��G�1�_�sbF$>�q�a��m���:�<�ӌ,N�E�PU�0��7H����b��������ù|x�I�_P��6V��)������F����ZUЖ�����SF�E�@3gȢ	���ɫ�v�M�׳�bw^;��J]���,��p�@�I�f[��ָО-8d�(�?PC�LdQi�	�t �Tr��&����b�\���@g�r}nYz�o�,��9hsK�f������`A�����f�2몢4@��Z�A^r��ڄy�lЋEǳẀcAu�A�S�a���JW4�ͩM��)89�W��^9�A�3s=�����O�]f�m�����Zw�t6Y�j[mi��B��Y�`*M�aѡ�t=9��> =sy�=�a���)���c����A�`�
c;&�KT��� +��Sߺ~5�F.ca�n�hA�� z��� ,-��������OroV�vj�X���C�`k>_0�ޞ%g��PD���l6�;����줲��NȀ�]������:[��F�b�d6��E�*�b>���t�)���,z}�~P��.����gc|7�lˎ�qj\����_�׬8�g3��/��TуA��z�Oy��j�Y�*�	���<x7�!y`o`�I�Ri*����e�d=���q�l�m�識/8[y��]Ї�ւ��O��6�����J�VJ1����|��V.�>��-�`��v�w��)��fU�����}j;���Ri�M��+A��'r�⍜��J���J���O'�>ib�@��(��k��Y$��N���������������5� �A:&%��$�����M���r�oK�'?�hr����FC���	�����t������ނ���ox��#�Ɛv6������������E�wؘ�bi�u�F$�����Z�,�0)|�B4�U��� ��N+���Xl�\O"�FAG"����	vӋ�h}Y���es?�ɇϳ�S�1$���4��� �>~���ӭp�jKJ7�+����FOyUY�F��aI%�\5�Z����9�-Ibq]k�m�Hd�U������~
�:�8��Q��-�Mﻘ����4}?�
�& u�?���?���.q�+��٢0� �T�S ) �Nܦc��L I�Yeu�^��(>]��|/ٚ���ny���5�.�[�,=�`p3Ķ.ϯȺH�s����ҽ�,��/&�A-DE�Y��ݳ�����'�̼~Q�ݷ�� �Ȓ�I��������6[��X��{�����n�6�X�_��,QѼ��\3Q���*�2���4��b�ٮ~%��֎#��z��?�2�zߞ�Ľ�z�}�2����U0��Yq��JG��YGF1i�p�O�r�l��t˺���
QÓT�q�(�"�"E��Md���<,p\��`$��	�xv&����%��r�����A���&��4٢�\�(jQ������*Όb(۠��6�R���&NϤө���!g���'�qаy�epk�¼%��B&�6
룂1*d���g+��Ӵ����5���M�-,�Y��
�t��^W��6JW� !.l9�Eg�Tp0l�*E���<�t��d��e�x��Ϡ����[q:9��}
h6�8&�S8�t�[L�H�/r�eA�U[y�JR{	�%� ����" C�e*��/$���9�ͷ��NqSb�n��q����l�kr�G��K65��ɰ�\��JV����񘊴.��׼��|�5�{kCYYA/�Ii�+Ŗ 3� �עVTK����Ӆ��&�B�9_�}A��w�=i��t��@�RWzo��z��F�(���u�a=���ߠ���jF*�)��e��i?�}�ai�� #=�B��\����4}��Y�������A��vk�M�*�Qgm������AwT@�J��"֭�ڨa��R��j�r��hɾ����hi���4!bw�)OU�{{A�h���I�-Dt�[.u�o��z�j�kqh�@N7
��r�Jc��왪K�D�`@�B^�	�3*Ek4)s�4�2�~N�)���߱g#�����;iC'~z�L�@��(�vtVSi��QEkBS�$O�	�!2�ʓ_�C���$��hK��*��=O{k1�!���o���9���xC2]�����jdٮ(| �8D���Fi%u�l �gL���Ve,+7*�r}��#�������L'�U@�1ib��43ٚS��}�N�pI�yT�/�ZO���e���+��M
�ʴ���c^��c>��;n�{6��ё�u��U�,;��9S�W���d��ᡜ��ZN�^���Iڟ�x�dC��H�tCF����o�"xr��ݟ���x�7X���c�/�;U������%��k���?���?K}w'3�l�g�k�,lM�ӥ�ٸ��Y%���ߨ߆HR�6t��OI�c���4sPD�̊��-��[6K ������!z�\`Zl1\��`�l��艺1��q��X�
@�E�_��:��T}�˴��:I 2JG����f)?��N���򜉇��9�N��p�����Z�)J�A�m�9�����|q!���"����*��a7��� 8|�*��6���-�[WT(�x�Z  �ɏm=z���RO$�8��O����*EL�����ۑJ��V���R��8V:��=O>k��gs�ZF��>��o"��^�N���-��친�8��g	t�od0½����>���L�7��^�t9+ʿd��}�=b���@s�<[���A�[ �)�I��6�����t}�B@��V@�.���^f	`A��g ��;�m-��X�߈�0����Z���
݌�������sm)�Ё&b<�p@oR��&��h�0��AT1�&���i|��iD��F�w�/~
|_��	`��*g�-����z	�	MÌEA���V4l@��8�x���%6����̪�=�&N�T��@i���X�?�N�5��Bu>h��+�*�V�k۵�v�{���=�[^Ϭ�����V�gsE|�yc�`3��:+=ц�%3.��\�����0�Ji<>�P��ÃCy��%��l�=E�d��T�}�-�,�JF��^5i�ƕQv�*�����}�
�݄���~
[�v�^b���GK��,��d�եg��|N�FF �M��L��О��3�i`$���α�Ʉ�ɴ!���4
N�:�N���s/J]�\V�O����əF�$Y�X�P!HN��DVz�M�P	�2�)���^1YQ�]E��T����C��)��c�j�j��/���pZ��$Bu��䊨��̺�w�����ѽ�e���R���啛B�Xl�)6[� p��NA	ƢQ#i��>���zں5٬K!P��j��H���S��h�<����eU�����z�vβ�)��~Ŏ+��B��}���Gl�yьn��T�.Db�|��l�8�y*[θR�������o�-��Od����1f�W�3M�d�Ю���;<��c*PEŚ+z)2B��e�|hU��6ʂ ;] � ���0�{���TqB�	�j�kN�C hJ;)L� ��A����]�_�o?���^�������A[�U����H]���]Y���.Tu����+���`߅I�[ޭJ�AR	5ە��*(��)�aBJ{4�JїZ���@�dol��ϖ��oqCۂ֪߯X
�@�4���a��{Gq(���Q��ud啶�T��d6���>��'�V���Nҿ��P���x(m0>�3���� �_-u��2@�yv�_X��پlO�>���6��&G��TF�����d���M����(�6�V������ES��FE�V4��+��D��#�{������S�P�힋n���ഩ+*�%��{;A����� ������D`��
�P��d������qV���???O�O�7����[�Ι��x@�-3ܹ�hq�M-���&g����#�Ͷ$I�,1Q5�5<�\j�3��S��?��e��Ӑ�i �*���f��{EDU=2���C:����آ*"W���)���&�[%J����,ǢD��O��*[af��D�|P�R �u��~yy!�^]���F6�u�����=�>��������_�1ǘ~5�h�he��z��1Ȓ�b�z/!i�������zʶ�x�v hK�Ge��c�͟����y?��KMb�^�m�WP�dW���dT>����X*���!��I��*\�q�'7=�Mg>AM
$���-���&6��!�}J%a5����߳����d�S5D��8��^��&�n�6ۜ�76������W8У\�Uܜ�-;�!Kߖ�j�W��$�wZ�����mz�_�bΆx
��A�79�3h@��ar�?Ǽ������7��]��ľ+��o�p���W���y�9�~A	��Q���Pcr�H͎z�,���Jq	�o����뽬+�㱝�����H�a��˪b:<�TҙWb��7�;7H��F�a�̑7�q�W������f�n��v���t|VG����d�\��x�53���CE��-�;�`�)�3p�G�mP��DP�ɫ�Fm��vT��BB�X���Z@����Q��y =p����Z�����Q�MO��J:�;�U1���T0�zț����U�qɯs(��ʃ�����٥�ځU�q�`���p`����JR"���o#�"�I�h �絹�ǆ\$�g�J]0�ج"�)3�a*k��4�C��}�ˑ�n�����)L�)y�����T]�ޛ�5`�e=� X��A�0#�����p�&(���y�=���X*�3�(�S���|}�>7�9��E�vCg�DK��w�^�E��Z�g����m��.8�b�\q趈�,���PA���=��M���5Y�oy���Q*��$�`�-�b�	��0����.4�z�iȢvw�]�ȯo`&)钠MZ�fr�^0�C���$�c<��S?�v���1+M*ۑ���C�`Yk�j�`a�Hw���d�-5Û4(��M�nP�ẗ
(��E�����*�ik5 ����n^��r���u~^��2���E�jm��H��	"��﷠h������T��db/8ǋ�U����ë��t�!/�=�P���������&�T8��"���yD�|-J��,5h*��79�ю�I���E��5�d.(���f�ʨ�.B� ?�B�Bx�h�ݦ�u���۴Oe��FJ���`��y�+Uz�$eg�E)T�	��؁����m|��7�*�-��S����5&�}��v�W�+���:��!���ڋf���+6@|�k����#����H$R�pA���q#�����:�%�M��qY��.�HM�o�� �ȱ#�&>��$~}/�w�}���l̀V��r0us�Ƀ
}�.�ő֋�+�6Y��'MN���v���L������ړΩ�hE��'�m���r/�uK���J�������3V7fI�W}m���z�i�ū�W,��d(�m}�m$���h�p:L�Ʃ���%�L��hxe�P��꡹(�~P鋵,BTuo�x/�K����S�=��[I�����?3�n%����Sk�-h�����+5*���'�d#����#���� �O�����3^�@�� %AlR��1��F���o�w�~���;��ˌ�*����$�6 �P~2Cb��dsJ�&8�/`�Gj}Rj~־�nv���B�BHvQ=K�ޤ�֩|ST�Nف��p�{ c{�2r(�:1�9�B`^3�s�lV��
P�����SiE��(;(:o��2#���],A?�&��d�4�@6�D�x���P2HFmF���bA	�0R�N{"�86��E�<e��嬑��<�@���s�b�s߁�
Y�	�6�������,H��R�a����X�!z�Y8�&��w�����M�`��3��=�C�^��A	z��g�`A��{�jT��gcp�k��d���5d�:�$���J+(�]潘��ի����L)2����dʅ������?���,@k.�o_��f�<c���z���.��\PR3�z���և9_�4���<���G��^{��Du,�t}	B�Hg}�^1�7�oj��(7��%{�KͿ�(D��&��;�$�?'�|r��l�M8B�8�ʅ\^md��p��`;�����Rr�D��ߧ��:��#<���]v�9�s�Y>s y�*VƟ�D���K2�NM�oδ�S���Q2��DN�*�nfs�Xf��A�K�Ä�Co��d�Y���c������{��b��Cfw\��}�/��J� q˪���W6�Xj�-�f
��P6"*�?Xu�l��+��M*��_���dXn�!"�l�RP�6�����ˣس�+��+����8"��D�I2H|�|'C�3�8h��[4q����(.�y�7��:*�#�_3�����p]{�V)L��T[`U6g�a�w��
�����'���T�~��߱��嶣�kM,�fsL�i{�US]�U���Kʎ��㏼רJ�I�)���r`3�TA椃uq�777���h�S��:�R>5I�
��zp*�Z�p���
���DKi>��o"�
b(,�n �ױ?Z"|0��'R0�\K�!��#Y:�{���F��.��-��k�	bi`�v�X�?gʐ���Zb�A��#��hY���T��Ӟ����J���4'��F�_M�^1��xKE�\L]ϡO��FT�����8C�c�3�X���39f���E��/>�G%��]��w��^}cs/ƀ�9�Q�܀s�TWQ�*��0�DJ�W�_��}�qlNL���P��M�C�5����6U�
�,6k���@ֹ�tP��s����Yׂ����T~^Ѱ_����y5��� ����?w�d�f:_ٗO�>ɿ���?���\]ް��㘃m�� �z�z&o޼��n��|������rcl6�l\�PZF�������]��P^㬧I��_h�`}-�k/*�,�TntHm�Ԇ�W� ,����t��gj ���#�)�U�o���qK��jN�=G�cy&�}$,#Ј�Pf_��8�r���'��X���8�`��
��1���L~���$`�㻊��1��ٰ�$
�f�yn�qP�:�����ϵt̪�тp?a������N>g�����?���2�zp�A��^P�y�ힳ��{TG=� 눾�
�4c��&E�*]������	)(wͤ2�(��K��&E?c߉@������o�o�;�bZp�k� 7�!�w Վ�m��w��=���O����R�d�F1�b�ր
�;7غֽ��5�/>���bg���m	�7X�Hr���U�N_��$c�OЬ�Ri<��PMP�'��nr�n(�9�Ǉ������{R�R��h�&!�,�l4?����ɲq��)��M�W����n{�<j�/_�z٬{Y�a�r�0�H���A�f���T�� ����_�$Oh�@����-���
`��GXDϗz�ۖEr���悲�KR����R{}f[>��8��yi�E)Y�0	�l&��h�J��u�g���u����L6&l�l6��b=�qC>$zF6�X���08S��z�:�N���x����e�� &�t���-�J��g������ׇs�07���wtfӞ�f�1�
������z�k�?�Q��4�I�1��X�]�q!W�ײ���*#fc�+���&�ofk�H ��[�}=���\�����B'�ule>�z�z<$���v�4�Q+AL����`T�@=3P� ��b���_�[ƏӤ͗��� m���BQB��LT�UM����?��\������Ĥ���ф 4Q����@_��i�j�q&���w��3���+]�ҽK>ĂP�fH�!tFRl�Op"���x�i���7�s� ��牂S�^��w��`	J*EN*h�X����O��０�,d�5S
p��Dbu2`+X�`�eLbA~�1�m�C�C��I�à�nM�+c���#��=�a�3�ii4`:Yo�&j�6��̟�Õ˚ʚ�i�"u,`�y�k�h�W���ܞ�%��`PUZ�%��U�v_�_[�ă�P@��c�D7���
��wt�g�;�q^�ۮ��.��P�Z(ǡj���IM2Į�U|��YL5�,�B�Vξ���M�ǭ^���TBo����/f���#��̙��)��Pe�L��L�ȋ���}�)��W�{��`�ݳ�����8G���7�jbV�S���&:�싳y����W��h��./׬PH�����+��n1 
�Ɔ��*�E�É�����р�����i�v!i�G)�hno�l�SP�Hd�3�!�o5���H@�Bp�)�C6�b��3����:�7�[�'���=F��u�B3�H�pԡ��o��)U��F�TDU>�f���]ҡBG��`U4
[��7�$�S��e:hXŬɁќ�,�t{9�KNt"8�7n����=>�X�`��D�7�
6wX=f�����@j*�q��Ay�����#�@� B��<X����(^����b�������D�� :� (���ā��_`���S|2*e�Y0�������k�x�3U�|6l���㣊o�7&S�IJW����Py�~n��?m,Nc���{���Z�1+&�q�^'T�,Bо�c�с,(�'\��r��u��`bTD��ghL�����(����@����T�[[4 ǐ4��S�{�����Mf08���]_.)v�Dvb:P=m���e�Vړ=6&��zQ_���W�m����W�[Rq~ʫZhՂ21��k �53*�-):���2H�EU��L�A�;�z���ʤO��UrH�� N@+���	:U��7U����1���5�%z��>��*��m��C��Y~o7٨	�8��W�V���~@8�3��i��| �h�
��r���? [�����Ff�%SGL��&�J
����YN���#�"��_���f�Խ:i��>k0F�xA���V�COR����DeZʨG�j�q%��p.$�ɑ6l֩�]����C��%*�áýUm�:G�頷��}x�Tʽ�N��<�[qф�bj���.��Ĺ8!��d(�X�����)��Q������w�c��@��/�o�
���f�>�k�.d� j믿��V��$ih��)���'߫NgK9�L�AHR�E� t{$:ݳ��+SN��5x��	��6`Ť�F�6�QE���ڛ?po�Ã�*[+B2
>ǉ5��r��{(��kx1���8���AN��(�T�""b�0�%t`��lإF���n�O��<?Z��&�chX�\�!Qnb��6��D?�-�V�
�Ǣ%8��%�Rm|� �w>�^�����(0bU���Z��JnM�m�Yks����$�f�p`��eq�U^V��V�j�^5Rg�*x�'[t���^E���֓՜c9��C�(��?+r+����E���9x_��"C0�9���fd޿� �������e&�����|��N7�t:E�B�3�F�Tf�f�M��y6�Γ���d�I��S��U��%�,�\B����q.���Y��;|OX@�?����x���͆~��*��Dc�OJ�5|-(�e*I���cO0 ǳݢ��@z�
��O~By��\2��3V�d�@P�gT�t��`s�d�����̢�zv<y�0�%������ �ǘ\?X�'���JÞ��0�3�	�����3	�yll��,�`��^�&&>nwS�͎��ᙕ*���8&�'��-�30{� +���0h5k�>8uk������t3*���R�=[^Mm�FY(�f�XP$&��4X��r�#��g %���.�[2g����1�.�.;��@�_�@aT�+Y��@���.ٿ�΢ѽ$�9�yt
޳9��l�b`��L�ה�b��⦲�Bd�ʳhϮ�d:��頠x<�0i�E6���VF��$��v�簉w�mh((��O�ꉂ=ˤ:J���8�5s��
�A�V4���{�T0��Cts}AZ�Ųg5��֋����x��R<�H%%ʹq^��I����$R{�R�*vR~�a���]A�S�"	0�YPP�B������(Z��+�[���
�b���=��t��f��bH>>g���y*2��5ك
8��Ѵ<�7gd�����-iX�p�lÐ��h��T &�㊵�da�>-��J����l����,zY�Jf4��c<qvFi@��X��M��f�&��]g�$j�	�C�e�Y�����������$a�!xyYйl*��Q<g�\S2�	L�l�qO��5��b@ B��% P�ZB�<�[8�|?����C��cp5����M�!`>��ug���O��h�<�:p���h�p,�ڪ�8�Ψ�L��x����	yV�R��c��\Y,n�q$yM#؇pů��Z�1�K(��5�H ���"A!�
�(mR���)8{r�Yd�pW;<Y�_����xD}����^'���hgO�$G�-��h��/���kGL`Ȫ�B�БO�cM�jv4 6�y�_�ɛ�E�{k�����,A��y��Xi�>�#���w���L2����P�㸊Xm���(M�����]i�	�SY�/�נ�X�d�.^D�UXH�ޓ�1(�
6� ����#oin1��.�}��	v��k/�x��bj�FjOV�L.�qN�s?YDX���>�i~�m֜
���R�����#�x=�`��qdo�B�L���1����+���\,u(?m�Y�v���yD�vu^5�:3�@/���L�N����1��ϐN�h�D� R�)Nn�iy��@Y�h����(C�)øGp�����d�;N	⁞J��LNϲ;B����[nh�WYHeE��w�D	�'�Ƞ*���c~2;�>��Ƀ��T
�6��⃬��B6�r���~Xs�6bT0�N�=&��Cu�I����rx�w:�Z��N4 �i�`B�0��IQ+�]w��?"�9���r>DY2�x�4/{�P�:�5F64AȕӁZmB#4�9 ��F�O�����$�����,�90:�.�:��gYLp��H�u���,���!w�W ��L!��dp������:V�T�]����@(�B
(�k�{G���6͎�������^J�?�H��|���ᳱ^b}�ޮ�5� k�������6�gPj��?d��c��֬h�'���*�d��	^����m����j�O_Z��I�	g��2K�2���y^k�M�7�V���`�Q�[�&&xt*e�ь\�j����0ɞP�6|���`ߩ���^�Q�3[p�����>T{�TQ�-���UX���
*�I�cC�
?%g��dV���3��͗�sq�_��{�<�:.�Xr����Tu�v6���;Sze_F�!�3T0�����G���:���@�Z�[����E����`��]�ɂHV�3��j�f����ӹ�0Ȋ�@'�30rǊM��B�p��<C�-�AavU�݂��Ω9���}�<�O:6�4L�w"�����%�"=|�?9Ȇ�H��;�ro��.<�iV��4��Q=��<q^�M:*��u"}``4��$����~����z��.��S���._/QpM�s�cd��QV����*���V�q�EG�j��XjK|6�Ԅ��k�-�Bs	k���Z�ҋTyyT
+S�rׂ�=��#��R�������9'��3`J�b���&��N�%�c��q��&�xw��Q��'�-4���j���,��8�h� �[B{	�u��������P 2V����,�ăҍ�ƞ8�1B����_����s{�^��`����c�QYf5��7\-���p �Ǻ����k����֗���,A��q~���Qz��u���W���U�����/mw��$��GѤۨ�BF݌%^�"X�88�7�M���oo1���_C~tV�r1�"b!%"���؎$u_����J��ؠ�z�=��+��C�������"�c�}��iRO���w��o��G���k_�k���nZ�^��|9oҫ��E�g�ސ) �M��{�EO�;ΦA�|sq��T�V�+��]Srs�L/���Ī4�����$����2�u8_M���~E����e����?�IΙ-�G<{�Y�P�h%˃ә�m5Ki�������67�r����۞@k�;�q_�r��0Z͢qD�,��y��2���0�����if���Ώ�*����r����*�7����I�_�T�` ��
!���^7;om;���&׬3PQ;��jw�N{OC*���6�g�Ĭ���{�X� k
���#�;rN��3�Ԙc1���3!=�?9�}G�c�yh��c�wz��i:�7��<�f�x�F��W�ꟓ+cN:X\j
[��O���b�ζ��␃�#�/�tÈ�_Xō�c��G�~,�f�OM��w�����;�)U�E�䃎OR�T����u�J����7������%�"��EE�ޯ�p��l�&0bv� �mo��)"hf(4�9?5
�2�1M��`�8>n6���Lz�o�O���˫~��#U�B�z��*u�,�r���k�B%s�ؓv�	�)��]�ɒH�'Ѵx�����4����տ�����Qҋd-`2�'�i7�t�_j��H�Q�.��{���������	s��x!M,�S�<�`�h#����}�5�]� h�fZ�Y2���s��ő�ȇ��x��:�0��qG�!*����@n؍�=<�<�;�xQ��[����r�Ϗ������QU�x{�:�@p
I��[�^҆+rxiu���be�W]���<ٝb�[{��ao)�����+}�L�{�m�z����n	
h��0��0����B0���	���)}|�LAxdU�������AR�(4A�BOF7fƂ�ҋ�e�E��"I�~gլ`�g�o�ʹ*�$����|����i�]��� ������3�]cBqv軷�1��X	�	}Y����B��T����8M,��)��n�S���,M���#�ǉA5:�;�b�4�F�@��D죵�O�~M)�����8�0��)U���_;�)`�<�?���[ΟO���E�p`8�//���k>�!�s���d����b>+[�Eϋr��Z�ޢ?�>䔪����x�M|�7��{�g�OX_%�w8�
M%K?٪�5Y��5z��ڵW%��O�d�G2��X*sj��jW@���IMvF�Ok��PFn�ؓ��5���i�ఉ�۟�@i@�
u�����9�q���e��{�ݖ9��|�@Z�q�� h~���dnM6��9��p5����޼��i�u53_24vA�+p�ҹ�I�Zil�y�� �����������Wr}}��:�%(j���y#.��4��V��}�R��#R�!1��Z�rp(��?'W� �[pju�|%�{<�NM��CmA�����͎-8/W�8�C��L��Jv YT\�N6�	w�׹*@����Q9�Ԛ�!�O)�� W��с�C�f�rv��&��#�uT`��@ը4u� G������=?�������w�h����.�����|�ӧ�O�emI:�Wұ����c|B�����3��IC�� 5�=�v�a<ڰI�o"���|� *
b|:!��4e��G[*��L�����W�`s-B�j�=�#����m�:iUh,���`I��T���G�`y���������Pα� �N��4yr��2����@b��:���+*����.������$�h���^���BA6[�@�C�4��lO69�����A 8j&�I\����[���Ѳ���5���ߓ�{�[��d�j� [3���k=Q����L�2������EH��:�%�a���H���cN_y��;.'X9����@��.�u�%�F����v�� ��,.֬��H�ge�mU聀�!���������#���j$�0b,ax(Ujq�h�bU�K*�0�Y}Z)d��6� ���>����q<�	�ٰ�64)�V�/��"�;��0�]|l�}���nAV���뉽ٻ��U���=��?��=#�[��w�1�
m��r;7���倽�G���@O&Q��l�	F�q� z9��^.d�8���=|T�;㬳6��I7|�Xhj.�ѱg|d���>]�~=��6�
�P+��l8���5;����De�sA���-.�-#����/��2� ��~�����ǵ��W��A�5���}�V~���X]��s�>>|�YY	�(�ީ�`t���m��������6�:�@_j�o� {�ɚk�o��q��`!	�`�}�����Cec�@����#*Y Yo���1��M
"�g��CL��U�_����Q�O{�ag�9~٢�|�{�0�(~l�>N5ε�O*�'E�g�3��T������!'V�{K4��� @𿘔���v$�h�nǲ���B���L�}v�#6V �V(��9��WČ]Pz<�&�y�ZIv�rNZ�G�������6�&-lA��s?ٮq���z�yi��zY[?��zrn��#%��5�j�k$x���B}�U�}r ����$��Eo�7k싂�~t��:{e�F��lD/3P��\� l�[yx��]KǓ�����;�5����c?��G�\ [#�o�f�zu%�}�Z��U6�=� Nj�K�))�U�"�g��)m�����H��69&F�F��B7<D'lSX�� d�N���Le٪����N)\�mg6���+�&�=��$�R�����᠉��\t�pr�y���ZR$BF�4"x[�R:m��f�q�E�s��Y�B �-�� �D����A8�өc�3��<mQA�2 �K�Y8�K�b6S8v6�5��&d�O��u���:��H����t
T���v��%��*�e��iy�F�a����os0�5I�IA{>@�u�|�=l�T�;�(�������`g�lt~F��g��m�|m׬ �5�ӡO:��V����Z��޾hI7��|Z���&)��Ա�t����/G�s��ՠ�\iK��qo�$]��iu`���#vXBiTu`w�蘡�D��S�E^pW�;i�*�;y�N��j�^��kΉ�9+
�y.�KJeg�1 �ɒ�`��ޤ�=�8R�N��s��)c$j��7���lS�k~>�S�)T�p�s����$io�x1h�ְ�+��Tg�@��F����mD��S��c_�}|����j.?]d��ު�]�=�����J� �z�����#�s�0�[H
f�IGR%�-�,��y�(�q`���M����vw�7��[��cg,���-L�7 ���|]��WFAź��X�1�d����6+�\����U�O�l�<<n9kh��cu�a3�+�(��˵�kd��~�y�A�@s|oI�_Z�*NM��W%m�Ǥ
�*���#��k��mǎ3�Р����1��gH�?�9oU0�5���2�����o���w�D\c֥�{�l����M|�%��3�=I���ª�}�K����@˃���%O�� �+��pϑ���G�K��w'�� ���!V�8� �ͼW��G[	��6� N}��WQ��@�}>ϼy�[�{���Y�j~�~�KR7�&1ָ~�%'M(%�*��6ZG� ��e �?XR��u�wf`H5z�4v"����8*hR������8I�� �XG����߳�������ӏ*܂�F�0��Ϸ�3�&����s�su���u��+������/�?����_ɾz�d��P	�lMF[Sp��(�	=_J'	*��4��l�`���T핽DA�X��knu��*�s9N'��;����SA�æfB<m��e�v̾mJu���a/�O��}>�����}�?s�=������7^�U[�LLӑ�7�|����dQٵ�ܾ`��:t޺��A���*Y�]R������/�B���llC��r���հ��Q��Ԋ�X�&�)�J�H*~x�c�bh��3�<ҧ����s�t������3�dg�ò� ��.U?)(�9�G�B1%��]�Xؙ|��D/��0N�<��&�8�5�p�Wɩ��(Y����� *>�����rD�=R�h���|G$ﲽ�@��ĹkH�")t�k!I_�92��E��ţ�vI�lh>�ێ�m֞sB}��x����j��D����O쳡��a��2�2>�u'���'�г0�~�$�1�����,R='qqz�-T~B��eo�8�&��_�����3���k����=Yx&�fMF�:I��T�
��v�G���1o���EN{�`A�$�!]��B�,R�	�ފ�
 �#�Z� o���׫2"z�*k^!v�&=���� �PF�����)X?O�7M@�*��n�Z��=�����A������4�m�����J�E�~dĘ�V6���2�aV<�yed�<7�U,�rZ���}�U�T�X�!�q�%%�R�[��f�k�4:ZBQ{b*:��A�)��P�t��������XϢe)��jrA�Ο�.�B��`Ԃf���r[��LgV�m���@��
�&�\�M������������43="��QS��g��������k�|�y��N�4��m^׷w��p�`C�=s�J��&Tx��Sŋ�;U�7o�� �pA09�u�K84�a(xb����8���._8��,��*d��Ӊ+@���P�2N��.I��>Bs�����f}Ij~�����*4�=�V�)�@q�%MpZ��T<\�E�����*c�%g�<���=P��4|�QPZ��y-�ׯ�bs��Յ,Ke8��&2��A+�rڝ����"��1�<[�I���ٳ:�L�i�X��� ������O�8" �� Z}���$�e���ǿF�r�q�����WK~?l�`B.L]rd���Ѿ��z׌⍴h�Ռ����>�����j&�M�IL�J�}I(T,&��*�G�^�:Z�`��"���LOy������'��J1�Ty5�3��Z�H�ϩ�}q�t���T�}K&-�*�wQ�o&�ٟ90��:둴�U-Ŕ���6����ߪ�.����˼�)%���C���c���n���/��7��G�� ��no�.��â�f\=��U��m'O�97Jy���O�>:��@G-�'^{�A��S��h��n'�p;�x�a�L��/ܩu���ӏV�HT����F���.hU X<�Im.?��98`q������f�$�O���M)ߚ��j����:��^g��e���{�PY��ɭs(oK�!�I*~,��U�I�k�^P�RgI%�z�[n�C�'�V�<i׊��J }~~_/^S�3էxl�?�����'5�-UA�X��*Yv7=�ў:ę�#v:�~�XrEu��"Ds��Klb{�*�e����7�>*���Y��ĺH��+���/�sC0�N'&cQBu�p�������3���I��t���B^�����rq��7�����R���}[],R����c��>�ՅRZ(�˜��T�_d@��I�����{5qc�;jT�wc& ,iI��=7T�m(�aT/.��X�I�'x]��:UO�F*�t}�&;�ʜ�l��^sPz��$�5Q�C�W�w���+CwS��VP���P�G4��0���!�z���EF�������@�=V�����E��26DfЕ���������?|j7*d)v1hU�&�Z/��IìA�d�m�JC����
�u�#�Gj{ߘBᇻ+Z���#X9��9� &�X���9�0Ne���U8Z�Ո�@�ȓ2�@�T�_�j��G��b/���Bq�X�T:����]��5��~�
~(�=��:�8 ��c�?�*߼��~��ʦ�)/r`�5�L2z"r�������}7�8wg�f�]a�?*�gfQ��� $�yϭA%��93��lyD �}�	�d����e���q���A���QR�NF�����I��u�&ς��)���{����~��-����ߕ`�����V�W`���3��l(T���K	��������@@o��Г�Z�dsy�A�M[��ba�+�TF�Yv\lM#oa8�� ʜ�8*6g���u���dR/P���_nn���Y^��I{<��&n�����j!�n����!x��PP�P�dS����+a�1*"1�����p�U�z���5�Ae�̗�%�&�Kv�칤ڻ�L���%8\�Á�8X�>kRjg�p϶���:��~�I}�ɛh��	��B��˒8�����>Ap�����M�uO�hN���eLR��&U/��-��������׼�l?އd%���c4��G��hFq�W����E�7�:�֋L��ؙ����<nj��������RQ>����`��,G���k?�d� �����n��0�pd
>�xd�OJ1d���-RL6d�I�b��}ը.��,�(�jN��9�"+��ϣ˲�Q����W��z8n~Z%��yT�S(u��a���'�y�gz
>M�Z��&��j:���N����z_� ��B�$\9Έ��zQ��=�Iʶ s�R��V����J�.�
��	�Pbn7��$��z+��5���v�QT�fL�J�8о+Y���ٓ�ڟ�d5��s8�����e�Y6��n��vQuC�ų̈́�� �U����ࠊ_l�5*6'>�yP����Sф����������9(�+-O4T~�-n��S�6�d�ZN�������ۍ5W^͛_��Bf~��O�6�h�U���A�����o `�sd�z����&��bF�nPi.�2�Zf�u���TLp�{��M(G5��rs��@���'�}C~��Ľ�|���l�>���8��_#�Q2�,�B�f	)�����2pQz����� � �q؏z�d�?b��\R2 �F��)O��M��o6;���rp��2��;c�Ưg�vyZEK�2�K��+�=�L_iZ[0���JX�LU7M~M����F<o�ɍ�m�h=1�S<�� w�fL�Y��6t��ۅ��z��K�&x�U��9�k;�3pR( �5�s��r�6���W��m�D�����K�C*<���nG<�C�.����
�T�/5���A�Y�eH���iEC�K��dp�?_B�/t0�E��!�r5l�ۋNV�N���|�{#�*E���Oh=���:�KU(������.����ы�ٝ�ُ5���z�����n���5i�G���j_��X� 6BQn��+�{C1���>��}rP}��
��|�.R@�؈C�M��� ��t�����<)ר�Ά�s ���U0!�M��k� �����~+O��y}�>�s�Uwr8<�k�g@���m˯E�*t�|.���/�f����ۅ�M�^!���E�����������H�&�c��1��8DzcJ��\��"�)*H˪��g�佂���E�7�l�OQ��X������$gہ�w"��T�i�P����E-̢��(��h���'*Uv[�n`9�,�� ʀ�!�X��#I�O����_��_�`
`u0����5&S|~��~��c�<C<�B~��I{�N���v$�C_�xP��B9����HE#�E8C��S��R��XKg��zڧ�V�U�=V'�r����L�Dd����@͚/�&~�U������g����Ϩ�m�?c^q���U��`��S]�M�t#�i@��.@cB�%XZ����T�Sy�I,<
L D�?�S?k}���`�N+A�G��X-��O��R���TrM#�ړN��+5�����`U񉺟�V��e�}��k����y⫂��P�^�r���y������
���sF�����R�����X�`I�y����A���7�������E���SvE�b�l**T�v��W�6���h��"���ؠ��PB�{!J�u�|�t+�ӟ�b5g/2Z���<��yE�}gЯi��-���X��]͵|�^]���%�҇e�1�Ϡ`Zӈk���1��c0�Smv/Q�d���r�A]�vj��#��g��_^ds�s�s.�b�~��j]��!T&SJ���Yi^��1����ff���ʢ�l��f��Eu�Á�N�,iB��)ڿ��\���l�&�g6W�E66�#�0l���..��A+Z��fSD��P�Lfo8��
��w���D2�}���b�Rdm)���4�1���;ڭ�Ԛ�T���IM�d��,L�A�*��0+��t��D�cZ��/YV�
5�v0��*�������M㕯�m�R),���-j��A,��4b�M�~#7�/3����J�U*o��6fϋ:P4�ZT�� r��<S���X�� �C�Ԫ��ho�+�'w�e���SԤ��9��f}^��Կ�1gE�-�%H�;��ii�����$7���%��  ���b���&�d�b #4I��"��a{����	bU[�{�{V�\J�yڏ5�=U���DZ�Am�`H�C� T�<B�f��Mvi`cepuyy!�7�2x�AU�nު�{�����9:�M!��x�-�m`wp�j��� +ԥڬ�`��[�&���C�?�9�,u�˫A6�[�z~-�O��Z�@k{�����̾ �B���g��딁�[�g�@ڇ4ZA��U�j#��7�
�����
��*H\�y9>�N7K���
T����	�%0�����٘}�q@�-�yy}D����dqM�;4��>B�s, ���H8u�R�:P��c�loa`���=�������T1ԇK�j�D4���]��b�?�����fu�_��߲�����Ͽ��˛�u��J�2_PLU(������'�����<���l��m�6�j�AI��Q�֎��=���
�zG�WFe�^J�L�Q�yTN�՞��VE/������fn�b!ى��fBUY/�U)*�Q�������]���1��ӧ;��׿�/�U>�~f�Y�6�n�>A5���i����k����-g)���H*�Z"*�H ar�g��`�՚����߫MJ�*c� 0����c� �?����2=�����	�f��&
��ZN�N-�1yJ�r�.��0k.�[�\9 �/����*��3x����]-��XZS�T�:��`dߨkkd2uƱQBQ�G���&���Y5(AI��� �'��V�:S!�Ȓَ�ɝ�L�P���i����A2FCɔ#1�{e&
;(_M�P!�T຺���~x+?|�J6�/������,��L�U�����/}��k�I���ܮ]!�5�t7��!>!uOyّ���QK������V�O�"�#<;� ���F�kPY]�͆9c��?(*]�J�3ke+4S:��x��[-�{ÊI���w�������H4���P��P��HG��_B�ѕfE�H8�����Gc1�JB��LoG&�@�xa	<d`Ú�4����	�gPON��:����
�*6�XIE�0�|�I�V�`%�3HA|�9�w����jR�O�
0K�m1gΏ�~)�fFc�5��+1�E�����5��1��[q���xz%5���ؚ�L�3��=O#յ]�0�N�vQ
gݥgM�A�k0�&�]2:�OW�"J��OP'�����oP�f�P��m�B9\*�qH�L���9^��og�PU�L��쬥�Iz+;�F�6КV�l� Q��
�L�����{L�A������gy��A>����d��9JJM��ڣ7����SJ�A}q��=|$�G�ώ���B��fz��X]��W�C#�
DP���������2�@��T)\s�X��x��-/.��~/7\]e`�����X�\A�a�Su�y%�Ug�GuF7&�M�bsy�>�o��%�^y��R�f��gރ���Z�QTes��sYe �*ۚ�|-�e�� >��q����<�N���Ŏ=�P<����b�c���H�Ԓ
�����_}�/�Ɨ@�׼XV^F;�9�@��\gm����O����9� �pus���l��)R!T����:`��F��̲OETt�Q�� �j�����{7�{�ƻ�o��G��֜��{B��[�JK�����(��d�s�{���_��?�7�������?������o��H���?��������Rmຼ�����A$�{����X,�@�
Y�$�i��O�N��N�2h<1���h#f4�7�8��e�禯f���(�Eb�'��72(DV2p%��G����6�����u����Ї�����Ó|��I��KY�d���6�I�5�jb������.iV{��[Jf�x���T'��+�=Dj.�b/m�el(��z�EY��\����W��5)N�r���  Cu����06�/�T��v��=��SE9&��'��]/�;�8ʹ���҂�Z�/��?�`B*n�=�c����6���O��JJ�6kRj/�d��K���mU���Ś	�c�-[(y����Y�%�PE�z�u�$�e~��kХW�:;Y=�����Y�O�v�>�\7����.<�a�XA� [Rl ������(�;ZņX�IY��4�VR�j�O��k�o/����bA����ԑA���w���i.�?)g���{Vm$�XC/oh�H:���R� Y�a+��XI	�T��$ER�d����ہ��y�V-�j�~
J�@&Q���/�G.����@U�qLf@u�GH��t�&���+ )�d K�eJ��9S��i'y�^��/��b�F���Mz��M��a�7�փ�3��:�
R�
#2�%%��u60��XI����)�].�����J���R���o�!s[hu�ߨ/��U�(Љ�V���wN���p�U��Ԕ�)�K�������n]�g[ i�>�k�ۘ�����;���Q�u����#=�չa��	Z���=���C��ӧOr{{���iw���z�L%�^��r�<�ׁ�1�l,��p�:�W�Cl����B.�y�v:����i�������#E>}|'����"P$�1 ����{�|�����H�R�
Hl#Ղ�w��r�*%M`A��m9��9��_	U0�Zc�K��yGܪ^��7�r��;����e�u�m؜��*�k�/,����Ai8�݈��Nщu�O2�5��Y�k(~�/�*]7|]-z%��(~�qvT�-󵬖ײ�_�|���#��I��0.�u�/9+)��-i?��>������}|��k�*F=���i��#�
2@�&�LȡG�������$�7�k��X�ģ����1��m~�#f&�L�p�^6��͆ؚ,a�A�фA:�Ai'��U���S�S	�Hv�)�ʘI�]�>�y��6Ù0b��l�޽'��o�`�Wҁ�?���\pf�J~��'
��W���Ϝ����8wQ�P�Q�KS���ZI��b!yk�5 �j��O��R���|9s	fO���k����R�V��BnPڻ�5��cCfG�];�{�~8e���7ky��F�l#�uɟ����3�����C�1�s���z��G��vH�&��1�.�^%���Gk|hLRAK~N�U9٠a�a����������|Tq!�H��T�XWPs.���j�Q��Km�P�#2���Y���i-�yS=#Iy|��km���--.�V���F�q�T�ؙ�h���0���&�� UO��Ks�=|v��^(u��z�ĕ����d��,}�rC���� ��iO����1*F����k�{s��)�z�)i<5��b��$I%�O,��l>43F���\���|��#��>��<�
)�<gc:g�/w�<YS3�m��N��&�ܦ�[�<l�V_��W��׶��N���u~#e�s�1;QmJEp ��#��S��u��4O�!��@)��b�Ҝ����Zv�*���:-Y����0 ����W�����h�S*p���\��%U�p a��Ň
����`ٴ@��r9��v!��S��+W0���� xh$��t5��N4"�c>^�ϴ���*,����avI��2�'XG��)�2m"P���<6�d%@Ue>�H_��4��F�-��l����@�eɢѾ&1���Wߢ0�ѝ�����9^Uh�W��`���d)�.����fcHM��sL� �_�*�P�R�x�h��5�
���@r���^�
eU�v�dJl�PA�7��<�
U���d��>΁�=չ���U9��g��cs���a���6���{(�b�@;R�ss�e�7�~,T�U(cNp�s��>���nw��|�@�,�8���mA��u������>�֮	)-��:��p5M[;�fK��@u$hJ�g��x��$��ZpT�����|@����\��^��A�^����F��W9���o�^�Y�);z��(�5Bz]���j���`���KWy^�����H���j���{'�q��1��DK9m�@����s� �sY}Xf@=���L�k���O��5g����z�~�F��<Z�%/@y��+q��{ž��B���_�8H��N~���ޒ�f�M�`����6/�;�����\���7�Q�ϣ%_�C�0������`�,Va����@M����b���J��[_�����mWL�;����I>潌c���#+Z�����߽{����;D�s}}���L~ƾ�>TB�G���28����V죉`�X�Fdy��JA��	i`����q�@k;�4)&z]�Lj�WO{Ԫ��H�l$�י��@�,�gf���wѮ�]]*��ʀ����\p�D��oP�;�r���~ѓ�9a��c�}�:�C�[��9�H�ux�`{�$����R_��#cW˂��oA�����1����KN[� l���s���k�������6��7f�xP]}��;����E�g>�z|�Otfjp���U��l���*�"eߪ����P_)��_/d�D�'����_J�'���h��Q<���r鼏���ݨU��ϴE�Za���Ó|�}����%��U�U\�~Jip���,���1-٩ �ɻI�S��5]�d���Cu�E5N���$�|��̰A�$Á�g��as-di&��h�?��ҥJ�>��h���p~�X ���������u����M���D�0㌍a����F�}6zM�g�W���@
�5�T��)��?�q{zz����l�/I�]a>���Î�j����|0����z!���z�Vˎ�Ȟ��(�~x��P�2�$t�h���\��\�����#Yf�W�5A~�?�)���!oT1:��6�)E�3rm�nP$C����D�7扠��`�,�k�K��dph��@��P#8��kZ��ؚr��v%N}}rݦ��Tث�g�"6�UA�{���2�����5��]({�A)`砫��qS��(3}}Ǹ�L��ˠ��M���=Bl`�Ji�O���)M,a���H���6�jҿ{<�	���%�T��p��=��&�,�h����±Y��כ� ��Λ��,�^d�5����%���ϋU�^�#�r�^d{A� ��wj� .��w�Y>��+%�W���s������+�0��]9_�_"�����%V�j�٧k�Z�y��e�J�����e�cN����X]����o�u0_��!��K�:q��ҝ��:$k�w_ J9��!G�4pU����/��<fhc�󫘤����!�8H��ݕ/�QQ2X��8�5�9�zp��=�$��6����~w⌿�˽�2��w2����*��A�J�~�}�+��0��]L�:���[۟��rnٻ�3�>:eĄJ�&Sc`u{fs�A��J�5��~?���dFԄ̐4!���Ez����4a��R��q��ڵ��\	�$����_+xf~ɠUL	5�������GV�o/?��\�8r0wwK����G��p4�M�󾸺�K�����3�ݯ�ʿ��_9����wx,E� �ם��)LB�~�鸒�}��&�������9i�'�q�2ִS��I6*v4}�k�=���}��Ԑ
�
�h,}���@$.k�����p�_ҙ�$U��A� ��"F���m�o�R��D�xܫ��JR��f��dL	��8�y]%ј��F���,2�B�v)��z�يf�|�'7]�D�q9 �}�k���j����
��~ε4�7b��(�#����=�gC8x*�/�&�I��48�b"g�ّ7���R��߲W�
\�ȯq���V,���5�%z��ﰾ8�ߞ �j�����}96�9x�0�/؏H}	M��~�E�Ϲ�"�hZ5��BM&g��&�!�]d��U��#�ѥN,��7d4/ː�MD�.,��μdZ��Ue�f�9~ڿ��<YiP�xy��|՟���0�\Q�iJI:5%zd];��GFR����gñe5K��^#ƪjSɪ[�֞��w�����NN>p�fY���ƫK���\-�l;[9O���Y-h�a�T�=��>�Gn}�� 
�����A�xBv6��f�D3~sd43��|���EYK�s�3�B�P�|l Y:9;�*E�Ml�xÁO�;D�yLt��5'�*p��ט�r<�lކ�dֻCaYp8 V��d�]3�>���^�i��;^��_�S'�� �A��r��kq���F�r(�w�gj�R���~%[�E�x:��/�7۽�$gΎS*H+�2YܫTΟ�!�k4����z�
�|���u����C��,��fƤ�~Hf#{<Y`1`�Wσ0s>�(�Q=EQK�$�S�=��;�D ����=�TB=�ؼ������J��ý|� ���F��U����Ev<Hr�%}�L�ݚ��X�fJ�*5һ'jo�_oi!u&��c���@힞Y=��i3��a���E�Sz�Jo�Od}/닍��F0�W�!���y	�@��wG��SRI���9��zp
Ò�����c��D:[���Z��YJ�dv={KJ4vK�B�@�|/�4$�����g)��UAx����Y?���1vL:�tѫ�Ӿy�{y��˶�d�����w?Z'xn˒Wx�U6R�>�yػ^��lX��}�u[����I���&������&�^h��b/��s�Z�S�������d��=��<P�61c@)sZ��q5@eu�G�')���,�WH�:����{w��1��I~���/��*.�����a2�����>�O��0�p���kA4K�����b� ��b��j���T�U��U�e�h~�ޕ�,��d��jH��`r��g0�W��o2��Ą�1�\u�L�I�,�U��~Gm3`E�	fL� �fd���]a@��.�&�/W�d@�1|��R̄��O�"Ȅ��R�VRl-X�,eb�'�S�s&��;Y����P�t�|�� %	J�m�S���곝�vZ�Fo���o2x����8fۼ��c�~�P>�Z�tҙ:q�����J���֊��vș�v�ҎZJ�/)���5r��ߡ�Z��w�̔ټZdln-�І-?o�;p�Cw �0�g��p=�QNZ���h�2��7C)�ܞ^���D-��,��¢Mѽ) �B����UL��� t�TDa�ϕ�,�j�s�D��Au+��_
ZR�8*����JA3�(M�������NU��9,Y{�L�ڰ�=�*�̊�7�O�~
�d2�/�x����>�B���MC�{�Z�\������m@|o,~h��y��=VH�@�p?[���e�����Er:�Ϸw�� [�J.VT)B~vs�3c��b���5�E@��9>��ax��!�� _��g�+��f��98ڮ�ˆ�Ǔ��3���_�ͫ+���wrs�*��L�jQe�g1�Ȑߏ�ک���+/3��\=��Σ���Ơ" ��D�'6A֞�\	��sJ��'P����n�)���V\1�k6O��o.��k�<�<�Od9�hbg��ф��}z���U���`������.�I:s8��M������>n����x�w�fa�T�Ē>���oJ	8?\�:^$k��AU��W�yW��m}�-���[2S�D�	������t&S���f�I9�"7V	*N��,�8����HT���_�F�����zs�A�qv����[I����%�S2�읊�u��.�0��z��a\e<�:į7Aym�񐃂������m$$`'���@HH���r��W���t�5�&����h�&�9�v�?)|q��y�~�P�7+i����&�bi� A��̲��|Yy���C���g���}YO�0��=�,>����r������Or�ݏҡ�+=u��*tѵ�
���r�]��c��<s���|�ɂ
-���"V&c�S�o�K��bm�|��m0����=��Q��{���;I�$?�������@��L@��p5e[|��h�す�`�w~�/A��Ͼ�pm���e�jJ�\�W%_ς�SⶇǼ߶�p%�C�ῇݎ�E2�7���mT9��L����I-�Zur����&�t���qO�F'ײ�� ��rMp/��s�k�%Ϟl�i��ݤնd�M�O�߃~�h���?�>v�%tR*�����Y��=˳у{��G�����vO��XL�`vq���μ{VE�-N���;Ua�� �R�C��@�z��pi�bp�<��|b��s -*�Q�� �7�c��	q�WZ|/��U�mg�,.��v���>0QB������R|��ɰ�D��<�&��Ã��x���L.��pk٬1��U�6����g��T�=�Ns�FI�x%_�QtP:�d�@�s�0�#�e[��l)�vTG��4y �ȶ�vY��yp-�!F�̶��@��J��iLZqŸh��R��՛��*jo|@�U�(VPӔ�h�9��33@��)�ϲ�}��L�6KΡ������r�ީ���KZ�H�B'c$�J��Ē�-�¥ ^m�'��%��)�1c�\|�c~Oj��'����Ɋ�T_6.�/^�=q�>!ٕ�'F�l_����6*V�Ǆ�9���o��:T*d2��~��TT�W�3�g[����>grnL�����(����z���{�y4����2��4��$�����DR�,K�SСΠI�{�^�v���+2���W�ꉆ�X�t�s�sM%���YUያ�O�h��Oonk��)�īKfN ɒ%d��s��\շF���x�H�`=;в6i��^A���@���;���2���6���R��̭�Fi4��C6���@-\�\\9�"�k���`�F���k��ܑ�2�w�]b6��R�o0���lf�l��d<wux#�wd�j��Rmr�)�LIXx
t�0�l�� p|td��[�X՗P-#%5Vj����m����va��\����	q�SB�d��N�򳺬�J�-��unOO(�|�"DK����H�ϕ/>�~��/�q������>���g ���g\�"�:_��;eEZ�`W7�c���z>2�c�����5�ʪSQP@����+��]l,C3\=I��Yr�=�fƵ�$Z��*h��:T���f��I҄ �)^�"+�����?�@����,���k�՛�l�����h�{���J���&���"�^�=����u�u)��xO�����V��s l�x0>S�=��VA1����A~�����SSi"hHJ�����\BS�mm���k+�[_����G���\J�X��(�_��a]�w���O������ѱ�?#�z�ZSݵ�;������\�P2�g�.�m��/f��RE�x�����g05:O��N�#��p���s��T�����2�����7q�KdBf��r�d�Č�O$S�^��׏?T�.M����`��z4p���M���k׹�U����|�}��(�R���C���%�B�yt~!T���2.��&5��j~��X���D{�&����=o��0��+�Ga��x@�-�aT��5X�$��.5qNR�z��E�^�DFT�A�O;���4V���\n;%_k����3��\�TX31��s��U�Tv(����j�1����0N  �Yݲ�+Z"Ľ7�UD�S�Iw�w�k��O��۠�Ay[Z�3$�g�����S�L��.�ߨ�A��	��$�� �[Mؓ���R���0_(C(_/�?J�wr���C��k�A�xP��}eg��m�
U�1��)�#7[��N5�v��n�S\}I�|i�ڀ��<�&9��}��:c��\⎀30γ?�sb��#[��q��oz|�՟�X
)�G��U�t�_5����)yi�T��� 8}�f�iQe�0&���i��=U�bW��+���׫)2^c�A�SS���~p��e3�$�a��'Ԉ$s�"ݐ%/{�SY�R�V`�[�ݛk[�R�ŧr��h�D��Q���s!�k�f�ݔQh����\�>U�P�B�e��R�PMQ��)� h���(�]$Mpq���
�a��-�Y�d�����bN�
�֤��SY@���>�5h�����Aއ����׬b�W��D�șU�^�R��X��6���=ۑ�$Nz ��HLPH�v������D�EJ����ѨE�R�핓\:8�� @꿭���B/E��-gI�S]^/�,h�7�����~�}��"��� ˏ�y؇y�\q髁�W��rh��es��o��*�/)��JC��fh��3^;��E���N��\{��ݮd�H5�@��	�ivy��Oe��܀n���lƷ�B K�us%�͚�5p��;c�$q!!I�􁨌n���`�����eT�cW�5�b�
e�%]�\+}��S���nYu�-Ǟ���|<ˋ�*�d�;X�$�t��!��k�K&���{W��i��50��e�����??g獤�.�g�m�8Ja������������uX���EL��K��I��,�������o�~��?��~�~��P��5cE�r�Zg�Q�c&�'W+������J.�}� mP����Q�-[��<�&uΘ���!T�8Hwڸ��	.�Ӎ �	Ca��ѻ�`Pq
�-���;�����C�AI����N:D}�C�l���\����3�Hy��ަաڣe�LAUU�F�s��8����|����y{EȭP�ER=�n������k�IhP�5�4g ��:���ʓ�.gҤj�-fs��Xv��b��~su-y��x|����(�?|���&^U�Z�i�2H�ڠ�M�� H���Ov�_b%�#{�Qt�N$ڃ�?Z��$~|F�G��ķ�^@rvMU�^�3X���SZ�x�%��F�ؤ�U`sC����&s<�a�,�xN4YQ�f��jc4Q+�HȞr\p�ʠae��gmP�-��w���a���{_�LQTX���3�$����3URb|�?UA�X��(�!�@�q���V�'��9}΂k
Oj@�3\��� �?��Q��I��G}_��\��QC������<�\&��SJ�����Xc��&0�
���c�������)(�TP�����;T��b;P�#�ss�x��>E�/gc�i|H�*��礪*���z.q� ��U˿�?_�ԗ��W�R���&���@�O�?�_��CK�$9T3��I�tWO� ����?e߻�f�Y�J���LDU�<�j���]����̊��p77SSQ��ٹ9z��i7�4�1���58۰�	>$[�^ߌ
��5��Ɇ��G�I%���c��N�ߒ�JHV��E7�~�;��5C#<_�ed��U���f�✙,4��� ���.G��٢��`��hNI�7�Ѣn����s�*���C�A��./���%�bd����Z�#6�F�lBp�\��(�% j�9�����������ߏFī�\_]�	IQ|#M�u�g3?�>)m��-:�93Xl�ר��-��
� �[FL��#��񈔼�س����F�ݞ2��É��>��9D���@���"��>K�́LF0��O_K�NY��("�N]�^���`�(��?nМ*XO�
'X�qz�������O
���b7
�+��Zf��Ҏ���j)܄��b�sb����յ�E�!�x�dgߍ��:���/�"��3�'?�3 Z��KFI���� Fu��E��T�˩�^\���6*]�"�3�9r�j�ؓ����
��`�_f�l�7H�	�tk���������\Œ@�HZKM�j|�K���G�:O焍�F�5��=y-B����<����xO�.�8�y#�������+������[�z��,.	Nv�瓯n���:�4;�=�@�_{�����1«���q7<@朜���I�}��&�xzu�\^�|E���הs7zr��}|�E����N)��p �ެ2�y��:��%��&�̲/X��׽9���s���
'�h= VT�1��,�W�`�-�i���3�&6�?1�"N�n�����`�S��4�7���7�7�Y`"8��W��W�����7���Y�!-J=�����O��i,s��/p��a�m�k�ߴW�Nm;�R�!��F�u�˼'é?����h�p�߼}���吏�Π7�w���A����=6�3F�e��Ok�$�y���4XFl0GxP���ǝh2`P�m���mѾyS�f5����?ȇ9~��p�O^T�3 2�%C�_�(��OGf��@VҜ��s4,=Q�@���^��jZ{�u{���TB��Vi���$m̀[��D����G��뒶*�Xk1���'�UG����D���+�Σ!죳�}������!�+E��_��9��%@�~���W������ ��>�K�O+����b`�"� kPN�i���i�2�ӖL��c�l��T�X��P>_)���,Z*Ƣsӣ�x	�s�9!��9U)����	+�,W��_��Y�!M�zҞ��� ^G�o��`i}�������߰�6�3:�P_�Z���٥,�+F�P��S�>��F1&&D4"��&�F�i*j�4������݀�7�/���\�q��t�>�L��1ԉz�M��w�9���Wx�~����}kc;e�� d��d}3�����)h��'W��:�v��ǄH�6�H�1���Ӊ>UЃa�ltgT�S�l)ރ,�J7��A|�C��N�X!�\X��y��ח����Ռ�=Ң�),Z�2��֥�u$ )�o�?��	��yc�F6#<`�j��?,op�\��3��=� �7b�Q0���D& ����������>)u+?X>A�H�}:�-�M9`�OV����Oʱ�)Ԑ8⪫�[#���K%rX�27lȦ��9�͏$UiptY��8G�6Č���yL��R(�,ܜ�U�^蛓f���$����6��6��~2pf����勯�甁,U,<0�Lr�^����Y�S�%��2QO�4��SDߧ�%�r'ބh� H{��m��{ˈ1�C��*U��_�n��z�N�˓11f?�t�ui-�ԡ�w#��>�:K��wn��z�Q$m�T_�y�����ڑo_��7r�?j�C��ͽ��ʠkC@���W��?�y����E[��E�CӼ&�K8_��h���|1����8.��ّ���������F������|�Z,K>�`
�-��1��]�;2U3:/�����>{�U�[�5�����Y��m�l�ײ�Ju����n����O�y�c롍�SLki�ÞȀ���g�Qp����#���܆(�4�����y'K�Ox��R�3*h*vR�~���)m� �A�W}g�{#��V�h����QmH�pncoC_�������Y��l)3Г�0���m�efcA)d�,��.8����#[��AW�+���i�	�O�VϗKf8�#T��k7�����[f}4c@�K0�ϖ�@L0:z	�"����5�1zVp�x��x�R�!�`~pz�f��R����拙�ǜh� jn��?����b��!K�Hk�
1�C�����&�Nb�v�s�(V��u`��5����y��!x�$�y�f|����`%U�N3�ؗP� ��v������;ƶ��	��|Q�1A3|��ՙ�.��ޑ=޲UX �=e�;��1P,7a��ľG�z����`R��짣��.2<s�ֽ�_1���{x�9��,)�H�1Bе�l=�xJ�ɛ��qvZ<�~)�����3ڈz,��){��ϓ��9=p��ܒ��
<�4�ͨqS��	��@����ږ�~��N�fQ����s�K�.1*�Ef�R����.Ι���uP�8Y$�Nn��af�r�!Z�e�{k�Ձb�P�2�vX��Q����Hu�o��3uPd�W�Nǳ�%��8v� )�'���,V -�O��4��0\G��9jC�õUB_R�x�-f�g�AT�c6>�g��4Ȣ� (6�BW��6}�,�\�)Jl���(%��Y0����r������|Eu����KÊ�¾U�.���nyo�{<{D�w�f���w �ǐ���T��w�M�����o���r�5�!J�,t�~P~z�:����) �,1�p4e"�H�i�OM�_�N�/�t�ӯ8c0�	�/?��O�kQ��-yr-�1���2o~�A�N����q:���vk���`�0�k�42���]�5ևvD&��A#�6���9Cqa��n�!;� �LP+��J��T%H) ��.j_9|�w51��M���,�lF4B�9����6�Q�E��Z��m��P�&�ڵ��]߳5//�N2?���S����)�jm\x��v
FWKc��1����$Snk�����ɻw��O��9�~à
V�c>�7o~�ۛ�l��Ջ�巿�g��o�YΟ����LP�6XfrˉOw&}>%�N�j䆿1��������ĩ�㓭N��ƜYu}M��s5�M\�5�q52Z�9An���g|��}�*{LQMuH�;��f&`������e��"d34��R!Ԃ�*��lˎ�:Ps�"��b�kQ�Q�c���0o��ɚ��"I]��diF�3à�d�P�BԑP�O*��۬���0��'��5�U��2`|@9���`}.v�
v�f��`JB�D�C��C���ޟ��n��;ᇨ֠5ǰi�S2�{������ƲaZ'��e�N?Me���k���]Q�'2J�,�����/����4{Ɇ�������fͰ�wV� �A���[��?@��l��}&�ϲ���`�h��Y��E����ㆽ�0@Yl�C6���_���/��-nt������6�53�]��l�T��ʞ����Ȗ�s֧�����<&2��N��:ou�R��0�w~���/_�����y���l��-j]m��j�= /��G4x�NY�~u��Ky���;RQ��w@O�hkQ�ɭ�	���rZ�v��2H,v7��[z$��:~��P���AjK�ﱌ`�V=W�߈��y��V�,�g�fy�MT�c�\hA(�����K=0����Q���X����E�����g��E��h���]`,t�0���x��7Vk�!"�������Tx4>vS�-,�9h�(f=�!*4~��Aտ!��Q-�!/r�~�T�#>b�[�|]E~%b��� �4Z�l�sn�6�,�����IЭ�[��T�.7��ߔ{;L�H�^q_a�	�}�xK'j0�� �3�r��ln^m6P��`�I6�,7G�l �qȋx�&��7�x"�닂�,�=v��N������|5�j�9w:��Lv���������B�4�~"&���g$PN�5p�z<�h�hY�0h�-����,u���}L���c$5�'[�k��w�KCsi����!�G�Ny��cU��egC������H�9��d�u}I}LA��:�&xD��,�3���ذ'b�"]Dj��KB?��c��;:g�����k��3+�v���s�BJӳ��m�F�q<�?kU��C���Y?}���Q��@��AOb����M|��0h&0���7 �<wE�	����6�h:v�H�!y0Jx ���L�vr��%hs��v�qKr#�w7�yx`q=�c���1;��)n�����޺�\_'t)�[z�q���'���'y��Or��@�ԡ�a+�>}�O�?�=m./^}+���?�/�9�|��5��:�������P���ts5`R��AF����ܰ��C��G�����~	�^�����S��,=���l��L�K!�@�
�����y��k-JXZ'��8�۸ Ƞ���Zn?��O߲6�+�}c+}��}J��21J��Ƭ���Qk��`;۳���[�,��@k��ǁt8-��g�YK�����j�
��9� "��\#��)�%T�ԓ�r��L�z�T��-��Mk�&���b�b1
z��D��SĜ�Q4�yM����荈M� �3������CG�<<HԞH��G���¤xT ��~��<yMU
�^Kb�+Hd���i8�d$��8=��E�8��%UXD�Kġрy�Z|༎��עw�j!_�L��O�����F�Md|�����Y+n��7y~~P@��>g_����D^~u%���7���E��6>�"�C���7�(6� ���eK�.�}��?A��7���'7��n�o���z��q��e���>RP���<z�����������J �hX���{����y��5�d��H��?� �]]�_��噼��y�ꕜ��dM�G�H1��uJk�{�L��R�R�F,l1Z��;
��d�k�2_;4)�
�ym��d�Wt��}�*F�� �
���@�R����IZښ�U0Tʝ��sN3sU#·C|W[�_I�ZiԃJ��U� _^��FP���h�q�Q���{Fl�d�Z��=oD3UQ�8�!BD����*�|`��.�
����S��f�m1+��i��%��ݥ��Q����i�S��uk"����t�����L�|��1�?�P:Z�}�Z-D��y!t�1uJ�
�t�X�ʸ��(���4s��t�8p��84Kг
u[�)�'����i^P~�S݈����G>7�GF��W�FO�t��U�`Qaݞ6]-�>7�#xUt(��j̛��U�~��By���F�Y�������cgu)�
'@�l�����ӳl�W*�ުL�`�������,g�?6��鍖Z=�t.�P�j�}Q�����O_�ZJ<A���ou��|a�:h����2Z��P�F9�
�j0g�{0��PA(z Ĉf�K��F(���h꽥�-��uE������Y*��Hn{P
ihvM�K�+C��ޔ+w��F�����Y23gL��Y
E�£u�3���}x`1#�l\vnv�Gك"�D݁�<�Ӯ%u#�	5IJˇI�͢�n�Z����n��!��ȯ���w�`����`�r&Uά�C�'ɺ�9��6��|������r��}�STo�h�]�����A�ׂ�V�_�B~���_�����7�z�y̵w�*?�-��>��|���/_�9~���j��{@�S06B�_:Zq8���l���I{��%����I��Pc�vo�,r�~���f�\*گk�Ufg;y��G����l�w�v��XoG�:�z�,b�"�EU�H�4�����1ѹզӉ��{�!�p� �͚̐EY�Rw���r��:��:^?�Vs��8ԥ���<6�#0�U�m�hjm�Hl��O�5-�Q{7�����n�l��hK�*�5��҇��B�Ehd���Fʚ-Þ��4�i��_�ǋt>\�j�5��
j�o�M�p�Aw�����	@z�;k5���T~\��pN�����*����ݑh�PMQ_vqy���Y�$���/g��/���9�7�x���{��P���k��Ƿ��=\ʧ��<g*�6��h.��d]˫o^��5Tg�ƦJ�����ϭ���#�.ϗrq�"�B���{P��@��L��a���aK`۸���{�@�m	�Ha�h///�׿�k���xN6��Wd=��|��g�������1��I\�b���%Ye��<�yi�`�A	�[DW���kO�t�׻Q����7��u�c%�F�.H�Wс���2iſ�G�S�Ϛ� �mk�&���d�:�[�u\��5���Z�5�� ު��2Y`��t	�|��������"��,��8��g�'k�' uJU�6�c��h�{��k��-[���,�S/ܡjh��L�t2��Dٟ���4V�U�V8��_~���o�������@Vp9L��������:�>�M>������fo4����,�$�и�`�(([�$�'�D�*�/���90�&��z�=��?���J�P�;t40�%��U%1ou4�M�kE͸������ �z+H�L��q���L4�Z���E�9k��~�lV"�����N�|�A�"��9��+ʫ6�Ri��*H���P��>�GY���ѬH��<��B��~(|:8�\i�d���y�A��0ٹ����=p�'��z�1VrI��el!"z8h}R��8�s�Þ�)�1�\��.���:��d���Q�.��46,<�I�i�K��E���{����
Q��f��b�	��z���P<f Y맒�w�����kX�$�H��}�ǈG����xO�Ú�9�V~dr�kkא�<>l�����|%ϟe��:�h4�\ǁ5���駴�p�v;Y������������Oy�w��X�f��y ����x����~/����l}+qz���6��0��vu7_'㚷ҜM�����4���ƻ�����S��nں���j��͔곚s�1H9fP_\�K�t�����]���ʙ��E�FC������?}/7��g �����������̋�6����(<�Z���vMTy�H��R�{)�>d-�m�9�z�}k��GjT����41�M��y6$���-�se��&&�,,{) ԳJ��>0�����eï��q����\����P#���As��~���c�Ǥ��l�+��c��@�]}rV�^#k��b~��O	�m�&� &�����T�hcRA���ub�*x�BgHCFe��_�����V��M2P8���:Xf@��c;?��5����7/20�f�����' ��
������<�`�c�Zh�q��q�m���Ys+,2��G��?���g1�|9���2_��[;����Old�� �>���:��`�Jeǽ��
 +�fp�����󽺒�U�eE�9}���R^m{��᜸���q�(�2�im#)�G����B�K��t���(6�D
�R���=�U�S^gq�E�m\}�3+����(O�q���O�ʗ��hBy��^X:��C`Y3�E[�<^�쵿���K���i�v�pk
��k=��>1Z�:X���#.�ɛ��i�+<��3��gSЩ:>�;*�ә
���15���2��zsȇLE�ރzS����U�uz�N��)6s����Hz�<�F�?��)H��5D�&�����i�ηo<@gz嘓b�8�P%Fob���~F���tÉhfǮ��
a�`7��Lb��8���FtF6t��f�D9� Y�ȸ�m4��E�]���Y��W��7֏#o�a�f:�0��z�~O����83jƛg��|�&�>l�x�3D0�>d�j��&�
XS�C�h"=��OOg�)s������3��c#�j?LŇ��=p�U�ln�ѻ��l���\M�۵�z��7�qg�'Ч�XR�Ը�o��:���"���TJ��'2�j��:O���)�j �<{�Um2�8���һ� � �π�aZ��.�2���uټF��Y
�h���?��4#J(6�L�YPg�7;��>�#M�9l��7[�������#p��G4!���?ɫ�|���`y:_�:������ڰ�]�4�5>��4���r��묶����sݭV�;���yxP������򗿑o~�ٹ�ZZ�`i�c��am@�,�EK}���~j�Ւ�z���G����ӝ��_|_R�=��pb��*���F	@�w��f�Nxe�F�T����o^,"<����6l��o_��wod�x���V����]���qG��R���m��O�Y�f�� NL2v�JX�[;6�F��e) �$�)�{�c���Q��3VG�s˝E<�6�WFL�kјE�\��])�σ�7��d�������RyM5�@j��X%�Td V��3:�B��z���IUlK:m7��l{P�ۇ�{ڧV�,��%җ]V��R����yv*���jk�ط2h��h��_�=^�5��8P�=�8�-�y!�sv~.��_�GY�&�2�f���_r�dx̊\q�Rk������l�	(d�Y�X. �����i���W���Ōn��`Ϛ��݃�s�ɠ^v׶���^�6EQ����t
����W�4@8� �Y{�A�����Zo��[8��lB���A�hGU�N}(�'��ש��,�����1�Khs�V��>����Ģ������85I�40�k��@07�mX�����뇒y+u4R�U�Y�c@!�ڶ�s�j@��b��,
\��C&ݛ�`�݄*h/鬫MmR0�6p�t��a%х���L�7�|�L���6eA��
Zm��˩Pm�l�l����`�Y�t��K�&E��}H���XP�B�:2�ɂ��`܁��P�$)!���wc��6�{�ɬ9��:�{���k]���?�i��$��qha��'JO$���*ܰ	�;��P�we��� �d+q�����jjMͣ�6;9����:߬�*����ک�u@Y�
4�܈�.�Zj�Z�BFy�Ӆj��@�=�GfzR ���h��d',�:X�B6��Ns�/[����D�M�c�w1!M!d��nJ
)�P�W;DJ�j���f �y�ٳ�4�򦲀J��U�b!H���9���+i���+����ct0~.�3y�=7�
Ȱ C*�S��Hʉ��G�����A#VL�4�R��*Q�Կ�2/�Vc7������8[�N��Q����۪PM��R��u�S�68�%Hi-�!�HXKiTݯu}ɨ�[������pT'��u]d��<;��7tgOF�������=K�MU��ȉ��oF	�h��,2U��7���[y��k��6>[���"6} -$�sn��
��P��u��O��q0E<�wi��Y+y����������2��f�	]��G�E�wQ��˛�2;�S����>��Qg3A4:;��Z&qi4^(��2�D��x� ���ݟ�;i#��Q�������|�+:9-��-����P6��kf�S>j��&T�f�qS�����&��4LV����+��?��<������6�3�8����ȍ�Ӊ��2'E���siZ�u%����s0��#M���}�����3d3���Q�p �:*ZO�k�i���J���H�ebpjs�Hm���"�)WzT�����d�g���ո�3) �5�M����;�y�F��w٩��;�"-��w[U����5J�y��6�܁�Jz������OC=����r�1�͔�1�,����.��oe�Ȓً�o�DQ�:�,a��y�t/�32 vC���Tq��v=�D�� M4�
v�ꍂ,6�r���;��<c 6��rw8�I?F���+*�n@~��Jx�Z)ɔT��<�
�`�����X�R	+���~O��j>���{��]�=瞾�{�&C���F�[�`u"F�
C�>����������oH��Zl�m���²,�ep�IF�C���j�E�״�;UG�����,�R�l�^��J��^���,����j	*�NX��@Z>a&��t��֊�(h�����\e@wq�˶s�F4p�q}Ԯ����� r��w;̺�!�j� �}4��3�����<��v����W�6�GZ_ �����fy?�Q��/��3ك��FՇ�L
AX#��r� �F ����l�E�%��`-!�����(È��V��r��΃^��8�Ʊ���
R2R>]��e�kv��HP��ۇ�|,��rCŸ�����y���,�g#��u6��)��H�u�T
����Io�%��S�_���
�x]y��������-5op\��$B[�5Z�̫,\ICx�^��b�4Zף	��a��G-����a1�Ɍ~M��v�Q�螚�6�'��^R����M��x��:��pr���0z�_�m��Fs	��R�P�8�����uag`�R��
RGO�8&!�H�P`Ȓ��QT_6X�K-�K�# @�%_89M�?j��:8C -��z�(`��έg_���6D�=B�4�� ��Ӽ�e�2o\(;���l��)\K����0@ %Lh�Ue�n3��żh�:�� ��^Qk�H0�djuX-W(
H�e��a��됝�w�gz:ѤR�xR�H���1��&�	p�S��|i�$��i4�N$ǿ��<=�/z��BcE�
�X� �zτ�BYCJmLem���U�h�yoU~��L��vj#T7v7FT+��S0���F����t֛5i��SɌ��*{;�N ����E�g3�����3bg�dqn��4*��gM�A������s����Ǳ��eb�|4���)���
��0��w�Խ:dv�GB�N��3P:���s�� ��U�$�����<�G��衿�a<��2{2y���ŋ�ôg������uv���s��jK�\]�6���T�l8������)~a.��<���[�_}(�1�B?��g���\D*����E+n��-��9�0�i���f?__S*�4\Ѯ��k����y���ɧ�7��N>�~-��C�dN���&���ǽ���z�E `Ͳ�K���e����wL��ϋRbVFGb}O�����Y���|�mP��l��"�¡l�Q�Z>����W��6G+���*����; C�~�?ț7���^�u�,�W�u�;h���M��8aQE�<���8Nk�:�޲l>������}�HГ��wwwCz/�����k�}����Z���r��JR[�	 +*�.����,`���XX�&���xM �>�`q��'��X֜�[R��
]=� ؚ�j����l���p@�B��!��?��О�~G��.�	3>�~�A,-#x��m,[5�@����$���2 <h+�����o���H¤d�
�'g�w�:fuG�#ج�Ɖf�&S�X�����m7G�� �dATc�� �|���
��j��&���Ȩ:`�9���G���o�<ۉ6$�����J�@�_��<ڣǁ۱�*~B�>B����he���Kz�X�Mtgńs4���$V��4D҉bj����ɭ�C�gч0�nx�c�3���3��bL�r'o�a�Ũ���X�,��dr����c��
&�I�B�.SK
���R2_~��oI������va�aH)�@q �@��^n�g�@�J>iN��/�tH?;���~p-�����s��M���-�Z�!_�����C�gD�{�{��^�E)|Y���8��;�k�ҭ�h=;D�f����N�%@�cDG`Ў���Q��|�I�$h��l��$t{����^��)a1�Q�<BJ5&r3��(�Z�Lp�h�*�ZU��"�ABF��������]�t~N�մV����d�����_��S�=�����3O&�gP�L����������_�����������z�ΊR�����K-�[���`�ЗC*��#F�[��
��"�JK�l9Bx�����hI)��X����+�]=k�zG�J�OuFp:�t(�ߧΜ�&ݼh�|�5{З"�A� �T�)k{�Lp�:��v�4��6��!�&C�NHK�d�{�G�w�$�\s�(��"-4;��ܛ:�'{�픒�4k�3s�jf��N�@��t�c����ë����7ry�\�|���q��q �������.,�j�j1<�s=��s�H�9���S��9�Kw{�wD����t��d{/C�F�_��)����2��� O���N~�����ݏr���PJ���U��5���C�9�L~�!��-V��9@b<�c����v�ӱ�&�j���oh�F���Q��L?:Mj�f��ꉠCgj�̒N���V����:�e�1���IJ1L��Iޣ�8��:d^������OpN�I�/�2��Yk��
�:���̠n���6���Ӝa���:u]���VM���Z�=���o��7��¡�[]^���Uޏ�}��%�o嘴gr#���������JOg̾�Zfs�������ācd�����)�����F:LE�kA`��{ �e�v=c
6:GVe*ф�p~���j?#��2�4U�O�im�,�
����G�Wx�vt#� EG��͎
� ��CCe��v:�Z����Z�0@Ά��v*��d0|O�X��gg�TD[ H��|���kʹow;*Hb.�*���y���J���\^���6����",Q�O�d��aR�,���~���O�G�v��ۓ�8
����T�QQ�՗��WC�,UP�Ujʓ�����-���Kll���S�*�,Ś�bm�t��&ڳ��F���щ�[;�6d��S��\���ܨ�S��xh�m��EC1�|e�W~}Q��QS��%]�,�]X#Z{�Ji������T�.��*c��4|���7w���<�X��ȉX#<]Ч��Z1�T�U�Y����+H	�"������zyD=ݤ�)�c�>n��R8^�m��#���o�|wk��Z���)�
a�E�x՚2�V֠ѢI� J��kN��>�R|q���@n�e��0d�y����j�9�Y��o�q�ip{+U�L�G*�El��RXӠ���| dQ�i��٠1d`մ��y��3�f��c�dW{~���_X����q���┋݋I��y1>���gK�#������ٱ��3���_y<�ѝ�'��A�P���T]�qF)�q=�_�վ��r� � �2����;X�~�P9��#W5�2(
�1����~�0^��\�,�6H��Ǧ�f|��3K��D�o�Z*0��s�6Xj� ��^'G��L��6��}v@[(�5������b?t�<\<���aOZ�:��Ւ@�9�}7UjTP�36H`#�%�d��d�	lJ�MZ����RV��0�γs����@P�\�ɳ_ɋ�$B���4�ی�y�,����z@� �������wuݧ���{J ����oQj�����p�Zk]o22B�?���A=�{��1Њ���9����6�w���������a��\_̧�(!.�f�}4�͂�Ҫ�(�h���I��$߁���v�_R4��{~f7,�X��L�Lv]��ubNs�1Q�����<�k��׀�8PAk.X[n`�:�A*
N�T�G!%bj��P��������΀+���LV���N���.��ؔ�*�d*�B�u�uR�L�	� ZMM�����WJ��{�j�����?�(޽��|~	}z�C4BUw��㎵DTVE�BP3fa�_�V��W��]\p�S��БN���`5�(��~<�T��_��Izo�GR溮��A�HZ6�͖�~���y�{1��㘛�A޿� ޿c���l�l���ݚ�R 2Y�)���#u�/0`0�Ь�����pc2�J�����P����>���������(���� ��L �ڬz�sj5��R��>s��}�]��n)Ȅ���W_-_�'�eA!�o֠����|ͷy\���R�j�;yX?�x/^�$���r~���|� Z�C��b;^�F��W��"�2S�p���s�?נ�x�e�'��N�OX��b�j�5����V�_\.���������#��Y�T�G1=�dbn�Dx4;��D�,���V�`�q�`'ۛP�)�e�2mëtAC������"xm�J%�`��Z�fjOǮ�?!��E5�u���[�{$$��ot�ް�RQ5S{A{�X]��k%3��zo(<U�iЦ�+؍'��~���?\y�*ԧO���M�ޛ�~EwU�ӆ�j�;�R�5�n�y,����>��x�Ŗ��B�(�:��������:[G����~
@T�e� JpE�|��m�1R��u�A�� Z��9�=j�v�����{y���j�A֑���k����^#���`�l6P���U4;����RM�����`]�ۋ�D�m�L���F���)G����A���Sh��2~�y�k��ƗB*t����q���(�)@�Me�j��o;���ʔJ0A�����x5�P���ǥݑe��C�b����{D���Uࡪ{J�q��%��{PEl��ѹ;���:!kEQ���<T e��h�B�_F������kؔ2hAt�2�L���k곍�<.(&��Ze�����##��ث�o[SKYx�����{z]����	lB��Y6j��>�N��ʑ߇�.�l~Lm��v�.8s�������*]��`�u����<,m`�F�*�cSfKm�`��7g	eG���*)��/��s>j�Y��s3�f�O�eǝ�r ���2����R]^di���&m�L�� ��3&z��*���y��;y��G���l�2�����ӎS�_��Q�"�L�c��$��;qf^z�t�-oc-�Q��Ț��Ԩ	1�v�=�5�\���=`�;��E  ��IDAT
���Kט�>kİ�Q	�^{Q�~/v�F��D��'f��h�����/.W���,;�p���l�g�ryq)�٢�T�Y�od3@e��ڂ$7��� @俛8�Gq���g  
F���{�����Gy���||�>��5A֡k��ٓ�섣�ؠ(��*��#	:�7
O��p�:��_��_|�fY�S $�����d����)��Eʛk�Lg~MJ�-�O�� �
��s�k|ǻ��3��*��+@ ��6�Ǎ���;���y��$�0�~A�J�n������D���|��~�=����`���hʜk�%<������o�����!��TV�:�.�Ȃϖsy�A�*� e��<�y_�w `�|�!XC�����zG�5���s���P~ߋ���X��N>���g�����9���p� ��n2��/����R�5^]�4ϱ~Ҕ��DU ��#['��PVY mYW��x.ؑ%{��_��Nn�D�7�߅��=�����+X2GjIS*�B�Y^�w�ly$$ ��M3��ȲKl�ْxk�TZ�κ�žY�	��9�ީP����l|�y����A�|V�]�p&�u7="�zf
{^i�d���T��J��6�C
<}�^;��8�E�As��EX��*	��Q3[Sϡ/k�Q�JE��C�����S�d�g�D�ר�9�|w.Ǝu�&2�`cg�X��:�)5���6��TiF��b*a�l�v"��6L��&jkEUh��8�DjD,����G� $W'|/TP@7�S��b
�0�ٲ�GoQt�&�~7<?%o<�<��������yq���Ŗ�Y�&���x_�p�̘�#�~̖�y��A� [PJ���<;yyk ���^`5�f�߇�Wiy���B�O�������6֔���{+���*kS�� j��9R��� ��'<Q����������x��_��-6q|0T:
k�#��6�fa=Ƞ}w|���������A�%�RT��1g�j�F���mu����(3�*?̌NRǐ k>��p{�4��f]|Cϕ�8A�Ԥњ��?�E����L��M=�/E�@4���F��5Q��,�(�f�T�W��5j�{Ly�#*b[�Jm9�*�m��U������M�i�����();����Uv�`���`L�?�����P\���=��21ؕ��x�����4�
����uAO���ҏT�).�� !�y��-������8�D1�ҁ�v4�V������fr�B���G���u��<<�ʇ�-��G���S�
BF���Q=lfq���u�pD��n���q�׳2dP�k�C��{܁&5��ݸQG��A50�c��=�a'Ѻ,d�:�5��
aZ�Ʀ��˲1nYS���Ę���
#Ѳ��LTZ��˚UE�/���f���{�Z�ƚ���'��Щ,<����y[3�Ϛ1��6R�@v0u�(���d�	�=J!>�Bd�A�~��}���R(=�?pO��?I�]��{�vhJp�*lJ�l�N��	c�=��o��F���g�״��2�C f��G��u�7���T[Ix�YOn}� p�	����m����F�Iܮ�h�q~a�NZ������_��o�C���
E4Vs�ZX?6i-۱�2���ŷ��7��r�Tq�͖���[6�UEb�8�\�` ���N���oz#���#�y:����^\��{�4k���YM5s� Y��/�q�Cp	}7�{� 1n��L�����?��$�#��b�0s��� `�V	gh���y��ej��R{B��߲���K&ƖdQ/��Q���:�=N�3v���b���L2a���R�4�2��̱&b)�1?j0�l��K�k6J[@�yB��6 ��q��B&V��lnk�*ۼ�[����%�=+۟���<8-�� xt9�S�.b�pGt
�X�hh���&g`�qF�0�ЋC�AG�4�ѹڃ�"Ì2ܳ�L#�8��RX�A�5�5�ѡ*�8fv��V�z�
��s�LRu<�&�>f�|L��`���(�|^�q�Ae"���z���P95��j��	�7�lO������U���dA��C^<���������F*C�e�t���yѤ�S��>.=�-�H��s����>�0��Fě;��wT9Wԉ�l��3��t����Z>\?���F�<�'K� �F�b��Q�lPe�Ɣ�4���.rw�?�m������k�BX��	��^#q�
��������Ą�Fa���h���l��X���?=Jr�o�=��^l�-�S|'R��?��y�UA����wD�Og�����WU���Sq'Щ{�<B+PNw��ԫ������������Jtj`�u-Í����`�����"�#eSp�����-@����TX�N��.\_�;�йE�Ԗ4V�_�'J���mM+(�@ 7v�9Y^L��JVX�qj�fuI���}�&�l2���A8�Eʾ���Y	�ˇ�>;>�K��&��&���|d疐�������ј/ϳSy�G#І��RQZ�n��E;��y�2������bw=��s=�>��s�;R���u�Y=�5m�F��9�%Z�qϰ~��{�~ g
bD�!Z`��@tt�v���Mv�2����$�w���x+7��Sx���fP _�@v�Q	1�UմUU@��
i�������(��G^W��K^'S^���ݩ�+6��L���d ��
S���{�C #?�{a`��ꨥL²��Jڼu�cP���c��v��*;�-� 
D-��3��`����k��x;QɌ¾g�� \p�l�N�< 5<�v��Ƞ����}µ�{~�pnf���n3�ܫ�3*g�k�&�G��";v�iBg�������E�
�*��a����Lu\�(�[�O__\��/���_�d0��,�yP���ꅏ���k�G颩�N�`����``ؾ�2���>v�ұE�*/���a�����@c�A�Al��>X�K�&��r��o;2x���w��g?�o&�)��6�;D(:�m�MI�?��	�Ǐ����w�~��q7P]��B��+X��aM,m��S���z��A8���ʡ�a���)�D{��c~�}�{4u7�3Ւ3�C�1_�jz�[�,�8����)2[xDS �p>�38>�U��X{r|�g-Ͳ�h+�mr1������b�R���Wh���2 �=���b��U?�4Д��;h�~�YH\I�5�t?�`Fu;� Ö9^أ����p������мc�_�Yo=dkYp8�3�һɱ�I: ��BGX��J:�Y(�pc�m�pө��8N�(�p�"z01��n����h��hL>U��R�jB�
%
nF� �����Y�|��$^8v�G^��KD�d�5�^�-��
��m�wu�:Ȝ�T],��>Tf_�h�U���@}Z具�6o���V#Ǎ��&/.�L����q�+����3�����NiMC3����.���)�X��4N͐u�>O�l賡��{�8��۳{�rL�g��y�_���Y"vySɛg0#��nv��nuȈ��lಝ�ͮ��5V�y�9cp��ǜ+��(�؈.1����P�e�b���i&��Y���-s��3Tp���4�?a4�N����I��	���O���[��U�-���\������/y|�=��AZ��c�}`��e�`P�@��X̚��<�U��O�23T�"|��,��~���ܢfރ�;z��
�<�� ��`?�:� �H�KC�3��P�)R�5�Mc��vq��H-Ƴ�M4P��S��N!dPjp:�ru�t0b1��dC�_
����
�İ�x�,c�k H�;��� �C4e�)#�g2�-H?Rc�Ö�q��Y?�n��c��?����?
X~�����Qэ�_|8 Vf�� `�w�{�@z��^���Y�� G�гM����m��zK0u�o��������[�!�0cV�e߳����@�]R{�9�R���H'4�3�=����c�M1���{��5ګS�~~E궂��}�m��6j�Rè��e�U�@Vh�N��.�4fS4����/�eu���tG���?�������1Ě�(�t��G �J������x����|�ͯ)@�����`�{�Me� nw��Y�#��%�e�l-XӦ��z�=8%%#�1������~I�;��6�΁m��*b4�TH4�XS)�/j�,�H�D�h9m�l>�m�d�`��R>]�����Q�=O�>vJ�H��?�k��{�1�s�|l�e��
x�d��&��(t0x0���Aګ��u�F�_�|��7�y�M9&���Zׁv0o)|���	��T"���6�5ێ��_�!�&���(h�"�/F{d���fų2��E��6V}��H���; �^L��g�yo���$�űz(���=>����جVK���`OQ̏��N޿{+��ޡO���)�IT�=F�D���(�Q�V�4d�`%g�IՀxRg˵\H��,���WE\�j:����ys�Nj�6��z��(ˬ�@��-@���[ ��_�^o=���p,�Ye�z��� ȃ	�V�7ު�5�&ME'��K��A�4���PT��Ib ���yl�r<��R�:��ۖ��lg�JB挴���{�4�`�&k>�강�����
�Z������bO᯼�>�ƴ�'�m�e0��ǻ��|8��&��.9&�"�a����wy��1˛e���C�p�������e��NJ��.�)B]��V�̈́Y��3B��
�]���Č�9����:�4Y��٭,Vf�28�E{0P����!�g@����KoQ,��6���φ(oZh3�H���e>ތ��ݼT��z
J�Mš� �+b ��J*7otOތp���5�2[c� �Bq2��*fJ�/}:���;O���0�ˏ�}m����_Ƌm}� �O�
<���d��"��M�&�7�um��Y�v�|��(9X�5�J���zf(F�5C���2�(�F�bDA!���Fi
���>R�Z,*R=�!-��h8`aƵú3���ht�zI������fź	��=��Pk��4��s6j0��FEeHcW8�H�݉��=�$�P�}�0�b�� S��b#Ga7����Gm��uXr2�Og��p4G��'/�?�#���G��ˌ����~z͢�� d��� �~p�@�YX��p�X[�lhv�7�J�����u��CaG�"���술�-rP�멍X�V�p%���)|vڸY��*u�(P��d�Ɔ���+S!�)�������ubM0�C̉����̪v���c��iِ9��|����7��o�9�X������O�5A� T/%�2^*X�u�u��o��3�]���7�_�^~��o�b�b"볹'xe$פ*��q;���г$�_����`��@�'�b��j�	GFc��'��Γ*����:���R���"�%3��nCQ�dʸ���f�p=���k�4�i�~�gL"3�	�O$�؏��} j�kC�Q�!�L�R
Y��@�L�*�7�`uLPIE��/� ��2��!�L ��p�%���GϟG�a���6fݐ�Ǭ���9v�� y+3�0��A�G�1�J*"p԰�X�V�X?ݠ�'�<L����
ޢG)�}���SlD�O�����ybo�Ή����5��.�&C��ŋ����K�	d��e���w��?� ��7yl�V�3�J�x�{�`Tq�$סq�5�QdY��"$VAV��c�B�1;�}���Z�ڒɟ�)U�&�C�U���<�<�T�ͣ�+�=0��OmK�R���ӓ��^�/����ۓ�o1��.Ν���%	�X�U�|!�����ۣ��ѦBp�O)B�_&�ֺx���I���O֤D��A�c��B�=��g�c2���V&�ɪ��p2\c�:�r"�MPT`v�#x;�l�����
�]o�3j@'y(3��RqZ�T�4��PNn�\t�����%k��*���������TK����?�%��J�:r�*�"� ����95@8��8N>�i�Ifg�a[�ٳHf�4���)�� ���c���� �]��u'�C ���JܙCH(j6m�P�	^FLe����q����tm��|���T��h��k>OǇ(N�	��\�QU5(�lr��Փs|_��:(��^�7�^1���(���W8�p�N�+c���5�R�x0�j�W��w���Qc�@�\/��U�}�c�n��lȕG�q���Rg�V�z�t��2 ZS4��+���9=n|)���i�N!� a^ӡ�D�A�Vc�`�i�@ �kuc.,��M�Y���:Y��v������6�Ҟm$N�ST^��:�W�De�,�v�W;���6OXd�� ��T�BZ�>+є��{�x�yȫH�?��A|��g�U_z��0
�����f��SAF{EP�Ez�����[��}/������D
�^�;�@����bmn�Z'	��Yv�����z�MR��E�(����fdjƵ)T����s��	��6�Q玎x����jpE���@���I��TĂ��Ԏ��� !3̒�
�Y�a��>���s��?�V����_��������B޾{G�����٬����bj�u��F3qbYr��B�J���R����e�����'�E���;f
e�罏�}�T����9hk2�����]��	�P)�A5{�M,8.Z7��}uu��!��@P+

//.duu)]��е�l.&�2pCG;���6k�L�*�5��w�P����Μm� 8�3����5і���h�uCI��h��S�l�נ����p� AV���7��!���|�LQUU����?�Ȓ�I�Rᇨ��,A ]��w)�ŒA~
� 4{����o��A�� ���^�i�>A�me,$�^��	���'S�����΂�(��2�(�N�,��	Z3�G��^�D�.�ׂڳ����������Oyo����O��G���?�f��4T��?ʠ�H)�Q�T�
�o�iK ��ٯT��	�Y}foR���F��VK�Cq��ĕ�8�\�L�O�T��9�>��H&������c�e�9���=�z���*�a�9em4��h&v�~>��zv�C+Yv�N�����߼h7O�Y�A��F�=���{:ܠ��6Ml�2녉�W#T4ǢD��g�Z�ɮ�<*��2�\�؄""y���[j�����D��\��i���7_մ5�\}	�76OPI�>���1j�a�;��R��Oo�)��z^�@-�l�S�Q���ΩMBCՃe�I�mZzg�9�nt,,D�3���0͆	uZ�-�i�T�kM�%*�a<u�� ���v|�q8^���B��ų3�}��}���' ZG��u)�6��c��E��l���,;�gr�,��S+�|N�l����)�:2�dw���w����� ���m�}o=8؏b�GfZ�v�`CH ׇ�V0�e t=�<�e8S?���R�{=1�lk1'5?2h<��ɾ�Ë����~E����j�s�{�ؘ�jE�z�jEe��s�����SOob��H2Jn���
�ݬ�nK��H���'𜡵���f�g&v�b����6����@��Fe���)E 6T���Yo�M�.i��Z����g�A���}6����J.������c�f����L}��&��=u�G� ��͗t-���jf5����2�7j� : i`��4oZ�#4&Dl���(�z�TG�����Ùǀ
nhz����GF�Y7�(.�,۟ q�EB�cǆ�I�ŇQ��}p�#s��Ȏ
8�=k!v|�f�5���?������ Y�:O���g��D����#�L�}�w�>K���6(���1�Ί��ا�Z �(`Q�����dP(�3;A�u8b�����v��:��f�p
���)���lI�n��
�Q8��r����#�ċڰw�b�ބ6�Ԭ�jC�᠙�#)�=���?��L�^�cNLM�����4qf���M|�4g���A�g���zٶ��<O��6�._(�P��F�9[�����@盯���˙,�9�r}q)��K����x)_B����&8�43���������ܾ}-���M;P����|���?����7��#��R�t*Kȼ��AFu�������A��20^�]jk	쩇���@��fΑ��6������;���{�B�9�u�q8t�e�u� 2?xm��Ы�X�.�wj��<�k�|�BV�y� [�������G���;yw�Nv�{�'��L�2����RX`��U;�ڽ|/���,C��.��� :(n�Zo!�є�R<���9�Z��!�c����f��/��m���m�7�M�1�65{�_�ǡ�l�^��v��Y H��4x�/�G�_���fPx��������_�6QA�����!�ƪ����?�z.IŚ\�Ag��v�K PQ�̬%eu��޿����]����wZ�����&<�od�y@R��W4�>N������`��jR@���'�y6�l$4$i�����]b0���P��2�������s��^�20��(����Y.Y��j}�10�vU�zw�c���m��̆6y?l������H:	��Ocڪ�r5l�F���1ϙ�i�j�՜�H3"d9�����)th#ݨ� ��D6���K���#���fRS��nK:P<�e# ���Z��(�jd�n���}%��R���O�s[PV!��F��|�|L=[2:��;r,�,�A'v�MZ����$Y�iM ��e���=�c��k<:<j4 X��&G;�ߌ�x�kt&F�	�̋q�#��mhgr��ec�I����{�9��a���6��o)������'f���Z�͑���wC���4����/�5X's�"����e1��R�{�Z;5��x1h
�����s�Ԥ���>{������a��P����`��۵��5�[i��T~/G�S���b��8-�e���0���ef�'��@�u:��0|b�2�!�&�C�xo��#�@g6s�٦��� �#�r�����J�z��sZ�Ė-硣m"I�o�c�-ApQ�Ų�y���V4��s-�f�`Sc�	���|�K�؈:; ����hO#�@��L%e�?)Bb�`T�4�f�Q��T�)PM4���EY�^��1�*2a����3{��-���ʤ>R�B�������NP�����'�;�_�C�0�O��Ga�:;T��cv�d<���`ak1Z�Á@�~����K�4��)��0ڭ=�hD��NX�ٞk��`�[�`�Pܠ�m%�f�2�+��Q�
�j:��q�zM�^��y.��x.{ީ�V���bBi�T�lb�@��~�
 �^\�����C� �ѿL�?hߧ`Y��	����?��������+y���w�������e+�q\.�(p  � �-T�p~Wo?e�s��eI��lā�Dl�5�b��+?|�GJ��T;����y��fqI��h��TFm��V*��k�/�������\��/Y�������ޮ���AֻMiGe�h�_7���z��7X��w�=
�f:v*G��0H�j	�T�w�}�o촷�yֆ���c҇)�M[�mJ�2��٫EiS�̶����	���'T������Q��x��-'LR����`�Zo�L���Oը��Xsg����X�T������߷�5�������'�1�~�N>~|O��M�~���r��`�*S ]ˀ�2T�f��k:o�Pɪ@?�V�dt�N���V^9��cR��Г��"����a���)}o{�2����FOdN{�U	����2Z��A�C���B��Kx�Km�i$Q�$p�$dx��Y4�Ds�A�-̦I Ȋ���8|&y� Id������je�ܞD����PTG�=fXɘfĉ�4�14�T���=�7�	�5R&�x1�Y:�l�r��1+m�@����]�C��cNw(����o���@j��R	��{ +�=���J5���0�&��̀;���^!Xh#�Qd�\���d��,��?�q����0jw��Ɇ�B��M`q1��������h��M�� �]��v��Od���F�њ�4��`t��걐U�d�C'VemxS�H@����ua���2�|�tq�Y$q�Y�ˮ<͐�~�T�a�FɁu=G��I���~�E����:)���LM�r񧠮�m�F��u����5����Ӡ��3m6���n����v���7Oy�NY��D��^���ыX�L�ޭ٨�Q��������҃�:e��:�4XƬ�� �<�,4 g��^Ay�Б}���{v����t���j�b���$��I�3OC��� g����J�l	�ղ�h��� J�M�-����t�/�P��ϳӝ�劁/���~��)��O����ޏBc�jQ�eD�1wؗm�=�H3cS�	o�4�v�M�&��߷'�X�����3�:��҃��j�p��H���t�aZ��4��-to��@7|��SgE?k�$~����@b>�i��W2��U�e���9�꯰��eʱ�M@�꘼a0��-�q��a[��W�p�~�:��M\o�1"{h���?���k�Tb_k�1���Bf��2�߼��Х<{v%W�V�my|�s6Q�S����wrww����CB�(����r~���!��î�ml�i:G(�8E����������IC��q>�w������	GU�����7�� 0�jJ�M;��"A>i� L�x�|��^�u��9�:2p��Ľ�6<��̌��;��f`(�_T���CK!��\�.�%����w�b�������L"��R?��߱G�W���{\��u��i�\�l Lܣ�b٘���`"!�;�J��9hd�G�f(%���ɏ�/ۇ�d������&��{*F�u�����nά�D�?�OܤT�)BK�3�%�0��}���ȷ���%l�-I�+9������t>y �1y��h>���u�Tx'��ˉ��κ���=W�S������
f��'�N>Vo�s4����>��폪'�PQ3��$�ba��x35J�7ڇ���Q,r�g�_�)�`����D��	����ТғJ��?i���KC3�����U%�Δ�9���;����-��8X��������:��<m�>%-RӐ�DM�F��ۊ�ra��|�{����<�0Z;
f4Rn����!9a��#x����Ngk�,�34C俣�CdŪ覾�d�r����e�ǘ������_���ҿ���(34�t;F��w:WB������vF�� ��Y�%�q"e���=*mF7ܓ$>g��C}���$%{r2��sn]%�� :%��_��������?��x�!W}����J���X�~R�5��)b�]"����;y�\7ߣъhyF�6��L�о���0������Ѡ�#@�ev����:t�XSer�ɲ����S���_D�jT}j_�����f���b���촠>O�W+��LI�
�<r�Go�[=dY�����ͧ�,b~@sKP��v;m�<��ܠKz��d�dl |��!�9@�8���L�+Ćt���甿�l�X�Y�Z�Z"����J`'(4�I�J�ҮE�if��,�`b���J�A�*:�8���̀�Q#�՗�U/��(*}��;1*]�މ��eK^ ����� �,5�>%I_�\��(l�ٞ���(@V�8B*�5b�$S��4���׹~\S��p�� ��z���"Jn�X�
X_k
a��Xw{wKY�ۛ$�����<��c]��
P՟Q�8�IL���2<�U�_���>�߲g�:d�
�=u6�l`�γ��v~!/����7�$�|�?=�d���"����:�&8���6�?��{A)1%� ���4�����<�.��9���yà���l�==�@��t����:#��d$0��A�no>��B���Hjv���(s �Ժn�Z>���M�M�Sֽ��!�;Ơl��Y�N�p9��9�/:X�O�K�3� ������J�2����t�̀*u�D�T�1�!�E%�c��K	ȡo�}�������{Y��]��п��h���ޛvI�G�j�G�G�U}�	r@�p��~���'��rH�htwݕgD�����aY�@c�/��def������������6z
��=2E�4m�]���L]P<���Kk���O"E���.���R���R����C��X�rB��-�g�Dū��i`2���@ cCY2kz�����7�n�E��&y8��(�AȾ�ޏ��wV��1I+�)��.�Z���TD�S��k��沪��)��CN�)7�p�re=^Ir�.`MsVf^[��w|�$e8|�����:XgNy3p�ǳ\��}��@IU��Xe����O��0T0�q�a�R�.< �[�\�\�V?ҁ�ACT=ϣ�%Ҵ;�f�{��J�n#\�s��>�XFWՏ�6Q<=��Z�՝ț��UO�'�%UEkTv���o��EF�dcE��cȗn�X26A������4`�LÕ7�Ø�ҦyBuR���"Q@D�|(nv��܁��14`S�?���wv��k�l䷳��`8�hn-A #@^n��C���;f�A���'�I���tP:u�A�A&��|Uek[�PI�Yƛ���ͱb*����f�|V��&�O�-֕�,t��S�_��3����^��Z���̶S�;sp�N�us�h��j�:�G�(D�`1���#:N(�^hmU�FT�Wpv�MT%�{��*�܇�޼�I^��}�c����\}�"�^_@�b�ө�YdW'nc�F�5�NJ�V3m��i+�
��^v-�U]/�<�7ƿh��z���qiR$��L`���衆� [Ț��)����}
��ޖ ��/��5�H�'��W��>&x5����5WGk�p�I�QK��r}�ԎZ��Jm�o(�j'&�қ`�G�E� �TD}�ΐ�o���)Kͨ�|��_R�ِv��7IՏ!�o�%�$��S�|��v�0�� ���\���aA+m^������f{+�o>>Τ�b}u�DhfY�w���\���L���}��^>~|�>h�6QW0��q���އڧӋg��������%>����/�!��[�X���l14��.�CPkJ�V��l��-�!�t�컂iک޲XYw^�0�2�,�d"�b�$�1�����f~����x�_QȺ����ț7?��A��F�Mk� ��F��|�,���ߢhba�
����㙀������&� ��8u����k��j�Q�!�y�DI���Z���t�-eHa�G�@燏�����C�#�,�K�OϬ���B=�r-h�s_��{f�H��d�Y�*�O����+A��A���H�6@�Ƿ���|�� �}��Œx� �ӟ�9g�x�L{b���	�Z�����l!^՜X{�(>l1��-k�@˞_��
�*>h�^6߲���H���u�2���坧�H�c8��G��U�}5�,)���:��^�"MZ�Փ��kt!>+�����h{��D���
n{;����棑*l�#J�{�`��MW�����;���6a�hXRˆ,b̵(e���/ћ������Q~�F"�]��.���A�d4�x�(�G�!f��F�1��?��b�� ��؂Yd�U�;(�����F�7W�n���HVO@��F�T��O�5�j�A֬K����¨�70k��Wk<D;� b������?�y�Os���j ����s4(8h W���UhW��,~`?K͜��a�1�{6�W���E��ۇ#�����hk�-��i�;u{n�1e����b2ۡ�Ś�}�T7��uF/��҄��y�3�y\��#�+�1����x.��R��(h�%��hP��ܭ{f}�ON�����sy��qqV/��OP��J���#��&:��w�����l���I�c�(jq?~x/��A���&��_������V@�{Fo����ZU��l��1S��/�M��J����"�tD�k�)��5���<���֬A'f��z����Xg��W�χ�ɶ����li�@i2�����r}W �����(����3y��Uqx_���#ʁ#��Z��a���< ,�q! ����Y������h��l<Ojs���GyI^�����M�?�6Ս6
�7�c�,��φlN��t��j$����g�^	3�P�C� ǕH�3�u�CmA��=��8`'D��<�ڀB#zLMPA�� �_=��d]��+�b_�/cs}s%��[J��v��(K��]���?K�����ڟ�z%���������݇�$��Oo�Z���<nT}����>�b$�����^k���W���m&�����������T(���\�r�s��>~�F���3�A��8+��2���J�.���-��ךi-��-t�Q�����MX)-u�����x@�hu�9�������L�
i�9�y�}�	)Xt���u���鋰�^ǈZu�L(�	����Ş[�ܓ�F?O�I�,�fR��J�#/sb/��ŭ����J'�0�3M,t��P���s�>�����u����ߒ5½i&H���X�}�J�s_�?k�߅��E�=���u]u�U	�r�-��)�+�'�YZ�'*p���,�p7�Et^v�� 0@^��3g-�j_������l5���<e�dX�+q�L�Dz{�L�K9�M�e6�E�g$�V��C�#=�8C;僻aS�1[O�}��� ����^%�}��6��<�W�^�G���`�.��<C�%U�/,F�-_{͑M0��H����s��� �p<kc��W�;S�3����٨a��rҚ,��6��f�O��2g�QnU�U��̈x6��P4j�Z�-���n���rWvW8 �I�|(�` U���6�d��5X�Kg偋8��L��y���8���f��-aOr������(��/�� '݂Rnм�����>e��+�u՝js_���&~����4y�����Jr�� ��g{�.�a׌�z@�FAi�]m�`����2�m��9W��N7p��]�-�Ҥ�F�;����)h����W�Y�J�P�I� W��С�f���e���5�5t+�r\\\ȳ'O��z�葜�����?D��P�x_��>q�V�MF�ϡs�۔A��t^,�Sȩ��xZ>��?�'���PA0`�NF@�AM�҇U�w���ُH)�S��¡���ZQ��M��s|oMxV�s����7:԰��8j�PK)�y�)�l����T����XJ��F�Ăs{V^�rR�qzvQ�my_���YN̉�hF��ޫ�d[AE<9D�NH~d p�	Y��W5ڎ�@셓ѹ�Z�:�dO���ni����?��5w��
{t!ޣ�'a����Y�Q��Y���u�W�D��le�H,,J�b �}4�6F�M�A���$3Ca��{��~�_<\�$?�r��7�j���Э�e���u��Ky� �OXW�꺎!�`���b�q֚V�����z����!ǥ3io+�Щ׻�5�v�BATGƞ�=�8�[�-��G����$Q�2�*�q�L_b�U�>�}Ec���1:�#a�؇�~L&����
E��!_�gl���!Z�κo�m�<P�������c��������IU�o�=�]G��x�l��l���3[�k
-$�	��u�}l<#�*��hD�-�։$k���G�)�Ï��6�v`�4��uk{=�ϝh_"Qt����%7�]Ek8��7��L�5��H"������Y�3�)~���枊Ӆ+��_&�9�RJL�Y��=�V����l���;�����N�Ŋ�Vw�d��\�`G�{�A錞���d�ul(7Z�7�u�%}҂q<c歷�8�`�]����0�J����������Sة
S�m�D���<����$ޯX�����{b�(us6n�b@�:wS�����&��@:�?	��GC��*8jF�4�d��O1�eQy�V�N���_(�Z.f�)@��p�r���I#��
2H:Ga/�#]��6�se)���ԞR��ԛbe�
l�*�e�s@YT���/����H��D.����0*#���""�}��ɨq�G�@K9���U�Q��?��t�4�
�r ���'p�>���Ժ�v�٣߷!��zTc�sE��Z|�7��<�٫���p @忽=S�>�C�Q*a�|4�b�Mgs�w�u�(ѰZ�s�^ݮ3It�z�]Si�ӂuSj�����o���ò�"
�Tqm�P�����L�=���Źy���)������Ab�;4�����.�8�� n�Y{ o]�⢗�aIa���@]>z,�����������e�|��1��e)3��b"�Nzs@)�����n�[@�׾�����S�b�QsF�mE���j��z���k���]��E��3�D�AoC��@UeS8��hVw%T=z�T�=&�^�(��iq����?��bO�p�1_ U��(�7���A;������'y��D>�-WW���,����sT����(�TV�5w�C,���2�����KY�)���`������IY�K����YMJ��Yd�[�	E&��& �������.��$�^����^jGq�u;�V"�l�֎�#�պ ����������D�[�e������s�<y,/_>�Ǘ�T9d{���(R����f��]�U71ѡ������Y;�l�g�Ƭv&Y]h�ɂc��K�z��Z�,��ur��Ā;�'�`�]2Ål�ݞ���%��{����!�m?RA�������f��۱+[.���gv�O	�����*%�p��=?^ �����b�;�ƨ���jE��gi~����o&�&�G���={f��ԧ���3L����g�,�l�H[��kN�@�~�k{�ϩ�	��˫�V���%[si�{?��>��~�J�[�ӂ�����w��:g��>m�(v�`���&�$�B)��w��yB��'К-�7��`'^��a?��iO��[�Ղ�o��z<�BN2h7+��m{���p�{���L�}^kv���� ��ww
�|y�=�=����e���U�y�~6oP��_��>�gh�*��hiIO�ɑb�~F\�;>���IW�jޛM�S,2E.���*����~�;��>C��F��j��E*f�N8'^�Q�51�� �~>S�VP&�0F&�\�be���fk�G�ͥ3����D��Mf���ؔ؜P���R�E��hJ����/.���G��S����k�u��%.��]����K�����Y�|����OQ������
��9f|���[1��ac���lX��Ҧ�^�T����ڳb_�S��y�VKE'����. }JQ�>��7{"��5x ����V7�R���tD��&�����갈ӓ5{5]���RU����L�?{*�^=��/���Ǘr~z�N@]��=�f������)3�y��4[��4�L��)I֦�lڨ�(N�is��X�pŇ�&��^�'���`u�l�FN�g��Jm��h�1�<�e|�l�E���m�W�����G8T�*$�t�#�]���Tֿ���J������ﳗ����/�8藏�	��Y�| �
_q��RNjŢƫa-���"���R��d�@���iw'���nS�e���v!�~u���:kh� ��Z�eMc�o�O������ ���� ɯ�z%��`ise��D����\m}�ހS�2c�q3����q�5��k׋��<( �@6�]9�T�n�V*PtЂz؃� Mَ̠�.����ޙj�4���4Z~��9�MՎu�,��A�=C�@���v�O�A=Wv�J�#�[�,8��:�~W��={�=�3�h��蕞J��������M�?}�����m[��wĞ������ɓ�p-
x�F{]w�s���c=�]��N��g�Qe�7�5R���?�C职�0�{���j DI�^Z�Y6�4�5��dL�(RA�5�uc;�m�V\��kj�q�VK0� 5��d{y�����?�w�"{���3Oݙ/$ܿ�b�s�S
V��r�o�������S{� �~��|��J�f����	�����!b�Nլ�;����q�@0z�-��Ɂn�$�H�_0e��W��T�ap�	�<w\Z��\Xj�0����"Y\�xVz��{ƝLrY���Q[[0ˆ�06b�hA݈Ҝ�J>`����,^oŗX��/7�ҡP��3W�&�Gb<��4)��T����:0V��}~a��Z��N	c����VExtJL�ۡ��G�����]1�ҙ�����ZlP����#�Y�;e��vƆ�ŉ�)�<$���ٶ�� �N�����}��-�ivD�Y3fT�lY.�/����6'�=�z'��ٳ����9�uq$k ���{6K,*���OA:���h}L���������^��������QAIޟ>Ԥ�G���DV��ȁ�C0�~Rr'BT%(9Ht���(? r��v��[:�;(q/41� EK�������<�(��1n�\����X'(Q���Ś=ǥ��M�&���\so2�n�;��s������(<?96j`X_�|��+y���\��R`�i�:�F/�F3�~I��z�}d�qn�b�d�ٴm�����T�旼7DY��8ro�f�Y8X��N�$.�ް�L��of�HTڠ֫�{أ��#�Vqj�������^��"%܄/�N�꿣�B�m�W��)��Y֧��ꫯ�٫����%��;�����:X�ԁt	
R8W{K��� R��qG ��9�m�����*�a�O��V�YG�ב�J���z[-vX1��[�s�f�i%� Ԭ=.@t�3��A3PT�ޝzw�t�AmLb��`����7n @�^P����e��p=T��mTcW����V�­��3Y���G�^��n�dv�,�%AuC�`�An7�E;9�WG1W&�A��N�E!x����c���Z5Ss�-��}a ��`
��⧱�j�򘕶��URw� ��\��D�c,nٲ���Y���0��I./Ni[���X�ݤ�X޻�N�p��q���BF~�ީ\;���)֍ʣ��H$d�!��ʩQj����l��k���G�|�}��y�F��=�,Wʦ�O���	���l���^W��z�Zf�����gQA�G@O�W[���l������)��̆^z|hvR�k��Ҟ,{�T�E�?����1�P�wi~����q^� �g�yf�R!�}��W���/��\�C�sޮh�~c6FT�������oBG��ձDD8�9n�F�u����ά]$ Y6���v�����~
�R����. �f"��H&	t
7�bu#�޲���3H�.:NfN���5X� � 0��i+��b ��8���y&�
��d�M���d�r�Y;k��}���6��>y��{eOvH�-9B;i��-�����CW'D(��N|����w֫!�{}Q��G�X3Iϝ ��_����"d�s������ׁY!`F�lP���o���;�����)+GMU��� "1��������A�M�v�4�|����=���%m��;G ��p&��̈́�-��X r
��g����)>�yl�������� �f�Z^[�%�RA��̧�Ԕ�ZG)���r[��:�\0��P%b�}}1`�#��]ҵ�ɳlM�f�pũ�hUg�������'-E��P�P���7�p�AMr;�� �r�̋��xDT�J,G�.z2���S�/�7)�<��KCAcvvzV��#��ꇲa�f{���C(j.�<Ԓ5Q�hr(�ݰ�r~y,���+����;���G��<��&��1w�>QHk�'<`Lt���y�z,�~�QL�8Y-��ꡘ-��c@���r�uq�.�s=!`��~_6�[�ͣ���sQHGe��2��D]���-2�-�O�;,��␽w�֙�ᬀ��S�[���-����~=���Pf��b��һ><�j%��o?ݖ�E�J�[����ӗ�ʷ����ꫯ�|�k�+t?���z�ɽZ�������\k��JީpK�^Z�Z1g�=�����|��Gy��{y�����9w���]�A�v�[�!��a����W��D6���S@8N�A@�n7ڽp�onM4E�뾀"dz= ���M�a
�GuZ����;�Afmպ��398|I!) j����M������@bW���7o$_�6���JUU��< M�7��V���-�@��_9��U'����TΕ7h�{L��U�g�-6a�� �[�d���o�(��)-�|�!������\{�����7���ig˽����C��;98�,���>�43@	-Y�����Ʀ��b݁�D'K��Čx��\l,��m�q7r0L���p&������rv�.��Qtt�D1��i���6���>&���ݎ*��Q��
`	�$Cٲ��4�E����]�Cwp ���B:B�j��G���(�Q BE����Q:�!�L��0/p���we�ܒ��](��ttRa���g�Br����Y���eVYrf|�L[�izFF�M�a�O��q��v\s�͞��YDV���LN�EvJ�Yk�T�JL���k�g����@0�ݻ���O?J�6���o�(S��W�J�,�����T���3��3T�O�9hS�>2�?�Ț(u��<!�� e�|qgbl�ECw��`���去�<u�%������]������dΪ�B#���9�bS�Q'�i�mTۣ�����B��T�PQS!���҃����2�W��o��� `�� �8�l2���&�<��H1��2�ܩO�p��/�;���بƿc�SU��|���zD��Y#������J�X��<+u��'P�\�4�0���0I��Yу��Y��p�:�0K���1/;�r=�r���-,]������F�L�"�ȩ�[�y�D�>?Zw0�
vP�E���'��J>!j��y��2��ˇS�����{�,o�1��ւ!����,���ZFM�(���w܎T����=�����M�WĨ(3��(���i�Qi�Z���Ȕ�9[A��^[Tf��]�_&2W��82�	�/\����SU5m7j��3݂0Q�*�C��o��F���7���s�����M�v�}<�:�Dם4�?G}��� �Rd�?�����K�z����7�`4�e�J�QdTtf����b!�*F���zcu�(�����wZu�}�������W8,r����uB�`�]�f�w�@*�&W�׃�y�����^~-��HdH�2ʘ'��H�INR�4�
�)�A91�������	�2j��'��B�AB}C�2�w�ؓ0���ق{��:�(��m����9-��-A��ω�MWl@����PUa�O�kEPggM��42��l�ɚ��yGt_}����Ϗ��H3,�CM�Q��T���3wwJM.ˊ  �g���=K&����K*�q�&�P�����4�����u��_����� ������ƶ;N���Ě�Bx������-{Qݳ��=3Wo0��4Z��4H �ʞu�ҫS�&�h����xd=V�PqgbB�
���@yFCȹȩ2���3c� x0�6�0P�V�+�b�|�<���(@E�Λ�Z��s��kb�kd��	h?DfA�X N��=!ڻ4�{X#W=�Z�*�V{�m�����Z���܇�zo�U����;�F����hꡏ�����E��e���f�4���''��֢-��`o$��@ߤX�c��]\��G�7��}�~z���l�l�J��k���X荟��o��~���k���}g����$�2Q����C3��p5��Y��]{���$-�f��UX��ʉDg~�I3��i'��2�j`ܙ!7|R�6d[x(0_(�oޛ��>��d���J=�)!���@&�d����p�5�ҼvM�Pr��w�lQ�Ȧ`�d��dU��\)��y�i k�����&��Er
f���UM�2�\�et���~U<�m���T'1ل'`�5svu�Y�-|ŧ:1���:�h�X�C�/�1M�*<�Pm��}�`��R���sS�<��~_0�2g{n����_1�b@��� h���k$$7��0���Ek�$����ȸkZ���:n��"~�Ul��c?���o��Xr9�K�6JW�J��n6���7 VC����ޔm�c�\�J���z�D�\m�<�t��ϔ�����g���G��d�+}N)��~��<}�T���[�MX/_�`����EFC�=9ծ�-q~�à��+��A��^�����R�F����K��@�x�����L�={�\�Y�Rg�3�f�^�@�Y@���l����뻡�|V����8�>�f�u)0�z�71�`W���5�@#��� ��^}]��K
�I��j��dbEa� �>���]���|�L��3@(}��~y���%�:>}@�e\�p��6���p�e�^�`�R�f]e��8d3��7^l���}�,F؋��9��ƍT��0��o��\��ȣ�c9:X�:�I}�m�<p�{��߉~M���}Y�
�&�qj;i� �=E��� AR@e�nP�1
�n�6��?���_��:.�:��A18���<�x�>S��x���8�6+{X>����.�'��2�]�VEș�Pd��sk��
<h����`D��!1��s���R�&���9�?�vl�^�9��3jo)����{��k�Vt�k��z괅lL<Rᨀ���g�a{�c�YJ�)͕/�Q��J�	�{�bR�qk��y�'��)9vZV�gat:�Y�����Sy���B`��Wii��X�Zq��o��"�:!E�1P!=\Z=��X��r�dMdu`��_*�B���!���O�G\�������OSZt0����w��v�l���B"Y����$�R'xM�丢J'�g��!U1���_�K���G�aB��s5,I�V��@�Y��0JcE�"�nc��x�8��dè#�������3V��.&�;��5��L��-2Y��'�ff�T��ˤ������/&������<Mw�����|��=��j;c�����Ľy��`��N��^�-{n��{ϲ�t��s�@Gy��b_�HmR(�H�9�3�ڴx�s��lO�Μ�Y�G��g�*�k&��S��݆t���r�S�I���x�(|	�f��e�c��Q��������t���8"��O)��]\�G�T��t@�k�޾pd�~?�?c�!���n/���eٮ��FX-d(���L���>^Ζ���m3!M�-a�D��Yk������VW��NuXR�}-����͛���͛b�oxNR�;�Nl����������u,���w,�Gt�5��5�A&�u�^W���<�����Cp�Z��}�-�.���`��ܕM�Iq~��G�}���I���o�na�(1W���4=X ˕:vhl<�}d�kjv|6F������z�q��vj����*��K����i6(�h�������7��W_'�?-�bey˰�')��<�&�T�^¸��c������>�4I��z/vxxB�J"���\O�ui���`Td�7��+կ��:'�����n��6dh��Ḧt�2�}� Ԛ1BpԦL�X�.��7_ɳg���l��x;-翥��"���_�D�w����T�r�=ؙ_cYj�ٕ��ׅ0*�!�t��{��PҲ��n)�1˻�e���MX׷SrG�����< ������#@�g�#�n���Ь̤�0<Gd� ��B��9i���蘩T�lR�8S�b��7�jw��?YR�@��zqY�-��=����k�@��2�*(�d���&U�_��(�����U�s�=����8nQ�Fj��Tj|����|����7�����e��@@}��"����e�P�d��@A��eR��� �{`o�����0P�R�,�1֢�E�an<A�N��5xFL�j�^���;Ȃ�DrPS�L����DK���Z/ ���qr~J�����8���)�#��h���|����MDI�����>@����!R�b���+lkY��7���4d v�A��α�%mF��A�"��E�I��os�}�ȹ"H�RD�HI �l�I�(��z1��,ݭ|�F�<m[��vP��n���8ږpξ�����p[0^ǥc�f��O�/M��9���ʤq��\�����p�;��ͤ�o�~K,�U^����9�Y���lT��� G�.C��A�ܤ���n�s���)�T��Yh���~���Z4�{J���"*3��½����¶@�ǹv�l�����gG��%�{����*w�s���K�w��f|b<��4�l٬zM>��`|ᚣ�D��>��R���!�O��TgB��e�S��g�3׾;<~�fj�4�!�Ա���(P�B�k E"����My�R|�]�jX>���ȕ�s(G��T^�f�������������Mq@�	wF�Ȥ�LlR�:U���wT������\}M�uqqIP�~7&��[U;�RgX�n-W�w�ƸY���`?B�1)`�̋ٿ~}$��˳�������2m٬�tA�`�x>�ޱ��iA�Vd��I�mF��y}~��C�jU�̩���Y�ZB�{)T���g�X}-�~�;y����S�*��_2� F?���&h�r��َ���ط|K�ȉ(81D��
Cq�?Nl"v�be���{r��wS���ǩ�Q���bq[���Y�s}}#WWWZy>�Zx�B]�&�nت���\\���HP"�Q+�wtt*�xl��W	�&2���ݤbO7U�c	��3P�g���l#��tpt&G��rV�W<���������v#�߽���;�����>.���˿��r��ب>S�׷;�v uX�8�O�D#S*�Q�PӃ��"��-cY(�H&���@
���T�LXK��Fv�p��ݵ��u������LĞ��fp� ɎJZ�4G{�%���nŹ�֨���Mz����Q��L��@�1�r�ӵ6G����_��o�w��G9, ������������Oe�F>Xp�&{0�)���(x2j��̀ͧT��>D�\�O���+
�v����˹��ތ��J!l'�R��s�>��Ku3�I�� ����(�� �ZG���[���T�������������93Y Y����&Z�@0�ӧO���[�����r�~���vE4U�/�A�zp�IR��tu��y���z"�S�cP�|`d���7��}R�$���F���#�h	)'��o��u�kf
�x�t�LE\�Æ4�7 f�.9���Zj]�5���pq��ױh�CU���7�*�*���!Ґ���;�9��t�NM��Nj���d�����ԺQ��Ҥ���sj�+mX�_\%�qp�]�;`�i(@qp�1u�YJ�3F����Z+ب2�>�F��s,�}Q���Z��?�����(,��'h�����`�R� �.�� ���i�mn��gk���\i5��ϩ�����)�}\�T���]�����l��B��a{��[߃�1����,_�R�̾p���Ј5YL��/3�S_z]�ݱ���(�l�'=?�S�杣6��&���dJ�ؼ(��i��Y+�T���U��餇ЈxtSm�g1h���9U�� �'��7��ŋ���P�%�L�E�锌��B��|u�j{v�	}���g��j�NrA�h-
�:�x*��Ei�Ooe����z�Q��P�X9�&A��%��en�5��>�h�S4�g��|a�����s�*�k*8`�ҠK|E�!�W��>�/_ɳ�/�h�_*4�؄ZZ���[�~7���s}�Yۏ�?�
��'����9zj�b��`{�� �Yv^��;Ĵ�S -�&���2��2*�D��^��J�3&n�Ç���;���f�؅��G[:�~B�lZ�ܬ�Y��2�R{�u���Um�둭�B ���@*�Ԗ�_���Y���z����s8���~�t�l��ɥ���;���o(k~us#��G���;��G�~����$I���܎tb�h���8������l�!�zp�H^�y���s9)��7v��	b�hpJ�X�8mw�B��y��ѿ���3�q�y�@Y+sta�1��C]��[e�����:�V��[�~}p$���W���J��[Y_�9{�(Zk�YO��i<U��Q�k�� ����;�o��7������w��;�
���T����y�>��z�]�Z NUW�4�?�3m-j�vcb6��R���S�w�h�=�0ؖ�N����4��l�|���M�/'M����i�8�(�➲\�֋}O��,;�-�}u3�(A	<<:�^���R�\��ݚs��䈪��Z�ޱ��`r6���i��{M���}��~?���OIF�(���Bk�[�&�f���r��4R���I�����u;Ō�eVg�?H�P�>-��L��<J�à0{�}j&K}�CW3Y���A8�q���@,�����hIH4Wg���EQVj�C<L��|��I� R��x����� �N�^���f/����ݟ8�iGι����?7�[̃9�׹y��A�g�d����d���7�v����Z�߈͹R���0��Y��^��o��L����ך��g��]����¯�����H6���k�K�T1<�Y��>s?�m	���߻�K��ϧQ��l,D+6�`�q�^�_����f�|je��M���o�R�Z�����"uA�q����UN[����~/���v25+���\"-�����������~Dϩ�dF֕�2v��;�y�P����Ϟ�����^�
T�B���e������?���*�#fX8��������Ã��k*N���T�<{Y�ʷ�}���i����v�gF����ةd�F�%>Վ��\���I�Iu��z�mu���JZK-6����e��t|,��g���#9����6Ŧd[���{�8{g��.�������mBj�u���T��܋��G�hu˾8cgr~q�:&�,� �6!�~[�5[�A����� ��Ȁ�S�_oj˛��J�#�;{��㘩�ZiP���ٴ4a��oG�c�>T��ї�x{Ap��4ؽ��bI�I��:'�s�g�����BU��D����O�eq���5!@��'��鋯����=�/ �œ���d��U~|����?���G�n�r}}Ga�rY!,�B�]��Q��G����cy���tPOD&H�6�N�i�c�kΓY�GO�ՙ������G!ȚI%�I�ʀT9|I�g��_a_�_�-��d�����4PWX>{��T=UL����)��Wy�@��zDu:�UL�@8.�����o��W�� Z��(��?>B��%�%櫊�Z.a ����ބ>�PҞ,�µb�*�&�LE�E䬊� H�v�J�>L����^1I�5jY�_�zCn�����&⢭P �У/Ԩa�x{�շĞ���qy�M�] ��5����1�c��j����m���4�}u�����zf�3����x�y�ڞ�2W&��u��鸣U �q��ve��r��.K���T,�Ҁ�=�n�>O�ۙ}���rB߄>�\}�܈�D�������`D�1���<*�l?�WǢ�����sL¶�y��"���ut�������V��C#��=%�qrpA�r ��p��ƣ3ŭ%\���ߝT�I�V��Ȝx�@�X��ڥ�z��s��,�+��z�*��f������C�f<c�k�+��>��?�xꢠ?g�����goƻ]�����N�ٙxֻnn��&n�O�`�5P�����	T8�>��ᒆJY{��x �{Q=��/׀�_T��O����?O�,��YB�܊t�nG�*�TZ��)@���񆾍��nL�T��� �
�Qs�6h	�[�A�{d���j9��-���D��_�����wl=c��b2��Q�5bFۛnW�UW���h��k��7�����o6���X����eƱ<~�\>~|+ן����J�W���r`�����.��d�H�e��k8���y���W<��K6�K��ۯ��|t|"���]����A쉔r�B�b������9��E�w���)4�Y��>��:M�R���]:�9�2�z}$��eʑͺEC�͍t��O�Qzz�d/�L��������l���±����74 �B8��r"D���q9j��5����K
�R��DGLfG��:;���)��{�i��{����$�~��4��N,��qd�@M>=>-�)�����rT�긼.?�6��.��y�����n�����ObP45O�~g�d��b�:m�o����O����ݽ̻����ē8KƩxT[�}�/�7�6��!���� *���p;���P��j������ߎJ�Ml��v���"O�(���)*c��uHg �Ѕ����T�h�2`|d�z�`��\M�$�B�jړ8�s���9{��RI]��<KT�k���E��Yb�=��%t�waݧ-��=e�ҤA
�'@�Zګ&D�xF��)�UV�,������x�:'h��f��w�^u�t�=���R�V���N�w���k�{�w�L��76��A���@����j�:)�����b���4>�s��>�7�����7��Te0I�t�U�bJ46�F&F�0�9M�R�%2`�Y�������gs�5T���ubϮ08+�5����lZ/"8Q^��7�<�����'����u���[��)Ա�ӧ�\z������\RS����U��Ţ�Ցwu:7*���Ȣ�H��X釾���!2�-9�S��1P�٬�u�۩����Ʈɽ���\_DX�J��w��9������������m��д�.{�Y��*����_'�� ��~ Z:-����
���Y�NnlS����~���Y�)l�C�k�:���9�_�����Zb.(��T���v�7to�������1i�o�U�m!b���0�t�ȑך��qO��wf�'���Yur| O�\ʫ�^ʷ�|] ׅ6T7g4��pP��c=��v6׋�X����t��^���� z]�]<��O����|��Z��=k@�X�&n!.,�����xR�J#�}r ���&h�%}f�~=�Gu�M�&i���e^�v�����C9<Z��_��ey-V���S��Gx�q�ʙ�Ϧ��q{?o��N�l�}ߣ̡���Nb��D�YF�y�(��5�J��L�z�s���f;��=��WVŐX炚�)�s��vG��Z�l�{Wkgݣ��t/hM���]@�v��#�zv.�F_�K-����%l1"Ѵ4����N�xN�C,��H2�3�g�T �G:�l��i�u�=R�l��
"g/ĀٟT�UR�\�F�q?|����������rc�A:�N3�f���1�_�\�������ǰK��o�=�o�8ժ3kbY�R�o�Yc�f���mWd�_v%�I�)mM�2��Y�A��BvÁ�W�>t���0�4�0O@Ce�
�se�l��և���*⍣��1{¹X�&�f�'����5�+0M0�̏��~ ��p/�zi,�L�W#LW3���\ɰ�:�5�b+b�2�z��Wj��ٕ���m٢��R���m/���+��@Kt���H���,wcm%×٪�@��K�{��>s��}�#P�����&��HD�c1�RY��']� �Q"·Tt�Yo�����V��\�]cDdM
���(�i��p�Mj��Ȟ�>���γ��h�xT]e#I�K|��أJ��s�m�땫d�ß�U�}�Jߓoj��'Vj t��iuPg�O�MeN>�r�2���� 5(�-'B5�nr��?�G��Y="� [�T�M��U C7nG�y��lҌo� �<�D�U{q�u��3<8�(pcS�U�*�'5cs�z�ώ\o6��;����_p`��a_�>��zOq��k�K���R��r(�
��r�4<�*�x�Ѕ�=뛲���A����C��޸E�&jv ���JS�x���l�+�v�!�]���d��"[�id���� �G���sy��4��f�e-���k[,�),f[�}ۃ�s���̴:�$�����l�f��\�v�H_�)@��&���3�>c��i�9w>������\��L*����n��C���51�Nj��ډ�1���[:��t��<�Y�9�c��Q'"���猂��� ������NJh�}��Z��rMjhCh� �>�Gts��@� 2Y{v&q���쎘�\��Fڹ�5�5��q}oz��ĳ�!�ӥ�_|����P�����~e/,�V"Q�"d���Wc�S� b�q���[y��-e��PS:#%ߋ���AD�,Ț�h8=���
c(�=|2
������e���;�|�P�P�ޙ��ĠՆ��!����*����9�P��g�TI:�rr�VRb�A%;:<`@�3�.��`���Nvm�Z&���,�����k`Y9F�η��Df6�U*"��q
,�����@~-�?�,���xt!x����_���s�~��	�&��v��6A�I�hDrg5��~��(��'��~��-ܟ��v���YN5��[��7�c����?�;�o$j�.l=�F�MՇ�+Eu�d�=�@G��f�܊$�i�j�j875w���4+�{3�i�AUq��b��B��fk	�@U�����d�O�C�^�!y�(_&S��@TE�r!;p�Y�T�B�j��*-�c��l��)�C4!\�$�8j3¼[�B��	Qj�вr����}��=tX!2��bD4�@��ⳋ�4w�I٬���f�x$�5�Ɯ2'd[��rm��6&FE�
����YPұ�|�t�Ns<ub��X��]�GM!6��3t/���9�� �_KJ�h��nTC���I���1�z�^�����pe�Ze}S�J9?�$�g��H>��b2���ih�K��:�
0tC���9�H�j� �Yu����k-���Ӭ�̟�l�x�J��s�Ei3>v�]�^-�I�����_DL!���Pr����LS(��\h����RD���M�?��]52}�Tzfn�ۇT�����J{��+�@��vb;�4(�i�t]��T�>�4��3���yK���5 ���g��]Y���6o�lj$��3i }��4��R���v4�#�XL�Hw�@(�0����O��꣡�9�5��pA^������o嫯�+`��s�xۇ"lD���_��O��q�����d����c��l1G�~��Y&�FҲ�>�X.Ξ˻��r���7֠�,�����F;\����	T�m�����Z�X7��J2�j��|�Ty�?@��x�������b�j=m��垏Amu�X�1@�l)%�滨	�7e>�i.�"P�*{oVaq�H�Li�j�.w��j�>B�e�hg��b9�t�sb_��)ڢ��ڌG������侇��=�.�C���R�2�V��rn��G��a�=���2��%v���+n�W�7��E����D��d�Tij�t�Z�Z�Q�\��Ή:��*&6�}��my�/�.6�����iq�7z��:��lj�`8ve�G�|w��M�@��3V�5�&�a�>B�=�?6���]q,>����z��;�S�#�<o�~��=%iX��#���؇���5�(�޿���f��vh6�-X�Sx��8�
ا� v��h���.�ݙ-*svBM�z%��SY�ɲ��ږ��������õ���^������C����h6��ӫʓ��1�W�)�gt��y��^ {Y�����E���<�<���.��bͬ�fl]\�������o���\��� ��HI� �ĺcm����㓓2�sf�.�'f�'�8�\�	�X|lPD<�Q����?[�c�{U���J�gMt�����rgtJ� O*����,�zRv��A.T���e�?��S5�!@0������I�3��F�\P��1on &�=��uf�&���!��gSFƕg���Po�\�l�T?!�_Yy_�OKd��t����/�� ˘�7d�TYfs�,������e{� FX�#��%��L�Au��M4|�G�_�&����G�����b�m��x�p"�H0�4�w���I�d��v�9����1mF智��h!�D���.|2{5�a�� �fʏ����Yd?�"�g���v(�q��*L{��/d%rؤ����k�w�͝9����N�y��j����d`+�]~������� ��\I�Q�1�v�����p��G�;v�_�Y�p��tC�q4� @�4������q�qm�)̋��M��x�2�{͚�?�g��N�"���U3��9?��zbf3�q�i��?��8(�IB>:|��8��w�{m�ȷGD�o1o�^:��Y{��nG��:��M���4�"j$�fӫ2�M$ڨՊ���z��� ��9��5�q�r�+�3!l��8;����rN�zT3�i��4�:�u<��W����|�g�m'�=���T[Dtq�If+4B�g��=��[�8��W����̬�J���:�Ul�>?JFC���h�~ͱ�c?�>���e?����S��_�<����9����-(��Y֖-T���� �xM��6��wR�Q����"�Y�S�,�~�}�`��]�~z�� l�M~ݟb#�ł���(���a�֎�<��}|�^�����X��fcʺY�a j�v���8�����;��@�����}�Cg�4#Kvw{#'�'r��q[�|�����%����l�R�#���Ϡc=y �S��6��ˮ�<������MˡҊ舩�nC��kD��m5Qc�6.���>e��r~8��^m5`���뫛2We,�ɺ�nI�+��X�����2��0 ���#�C�_�
)�����x>�g��ށ<y|!O�=�G�.������<8>:f�D��ӓ�����vs�z�G�1��9/ټyk{�H����f����|�^�x̓��b�����_�����?+�_k�zZ�+��\kn��~Z]��F��=9[�y���U�I�\�� �Խ�AӾ��-���B+m��J���7��~�q��=f�:���������9����9��#����y��� �����n�)l��!��YO�b�4z��X��z`�a�P��\/h�1a6}C�2��k�*��z�����(jo��:)��9y��̘M��٭J�#���v�*0���Jw��ͨ k�Q�@��g���|��M�f����P�t
^MzXD.�D6K<�������qH�*����?��Zp���j�T
�E�:�T��[�#���b�w��ߵ��E!�?}L]_����T3xfT�	k�c�<��(��F7m�ɯt���_�[-�L���p>�\m���TR}F��q��h�\���:�v��w�����s=|\���L����Rj�+5�F�Ѡ�=�eS˲ِ��YSC7�i��&��5Nco���
��6峃^�^�a��r�鬗_��T<��(�

r�
�B��ڛ�w���>i]jfg����3HE�yoVy#i�@�7l� Z֧�TR+�FM*���}�>��^���Q�^��>��<�U�[���I�Q3��e���]ظD7�iχ�%��Z��	���j<�Y�Zź��8`�,��ӕ
̜-�	�7.�(�@�o6Ƅ��]]P���PU�?�ٮ�3�����ac *�ۻ�>\����@��� \wduf*H�uy7Q<J}�����i�� @2V�߫����O�U�RE�P�=.=��/_�����EP��}� �L!B�kR�� AӬ�����Ʉ�R9'z#]\^p�h$˾[�
��e�"�gF����_Raʫ�����ᳵ�U@�gwwI>�����#�j��i�{ (v��Z��ψ��/�f!^ٛ�\ǽD�������/�DL��т�	
������`h��c�򻻝lFd�(�RΔ6�g�!|�Lq!(�<����|���)�~���9n����|\�䚳ϯ�k���筡ݗ��l�G�%J��#S��:Ν����+հ����v9��g�l�� 
⡍Av��0��R�C"\ck���j�ic�y�5�:j�:˺�i7f���&hЪoT>��P'e����_@��j{O�C��a�q����CT1*�����1���H�h$3^�T�i���j��JG����U ʴ��s�s�nD�� ZF'TL��H�/˜3��̲XU��g����G���~<�v2G$�4�Y��~3�����r���iD��*������c�x;�䑅�� �>��A�T�ܹ�E�D8�9��a�yd�QH���<~�`OO���Q��
EuJ��x���>�$Aߕdq�������@���z�g��z$�W��)�WZ�{���c�C �pc�z&��!8����&��@�q�])�S���o�r��Z([Si��6q�X�����=��S�]\a�����E�?(����~1��ej�������j��ug�MYµ�2�x{�����M�ܗ�s���8�FBqޓ�S9;9g�+�U3��]�6�e����ڣ�3(�=�\7/���s�Px�����|T�m�<����sr���]g1���_A���ث��}�]�vp�Eƅ��_{�:�U~���w{O��9���V�/��{���~֫zϮ�j!Tqaҭ��}�"��k/��{�"�0سP&�_^R��0P�U3�����y�}����B������?~/�����+R7P�5(��H��`�j2K��+��jϦt˲���������ȧ�t�p;+�ׯ�uvϯo(t
 {��ʂ��2�"b�&p�s�2V&p���X_48���;*���6@><>����7�?��3�*i�>�g*�d��|Rk.@���F}Y����-�N槀�}W�ɧk�d]]]����@) �8Z		�5�eZ�#��sVd\e*�n�{�l"���y6�ԉ�>�F��p'b9p?�?Y�]�+�XQ�c�lX6�S��b�=��|�@^�����|b�/t$H{���NE���6�Ȅ�����k��ut�ۚr�I�/���L�L�D��P�m��T��.m>�v_�g��`���L��[��_��b�`b��@�Z�xO��ʝ����.
�"$cv*�}�=3i�V��f�C�{��� �����7�l�1E��0O^�YeVzA��j$��܄�?v��E�c�\Dc2lԛ�;	���V����I	Ny��<���9� ��}�>D����.�`FYrYـ�Q�9��E���FH��
��ި����dlm�ʓe�P��o)7��(~���ؑ)�e��Z�ǋ��o�J�W�	 �Z��!2X�'�LFz�+��:?�ʩO5E� ��㾛SsF��d��AC�(���믋u�TqMih!2�$([Ɂ�S�<�����,�)��D8@�ť�Q�v�z���Е�86��1x���mwJUL)�>�É����0��?s0�x�9��{�
|D$ސ���`���`_�^ǯ�Pџ��(LY
�x���N���O~`�l��l�r����_���6�jШ4��?�$�d�>h��.F��zf�:%���Z�Z��ᱬ�>���vM�e_�?G�l��/E[���? �S=����Y�Úa'��"�.��3[_�(�	�q9w�+�k����mǭT�_�����2Y�>R?TD�\z��fUf��Z�q�:���?���>VŅ���z'}q��]D�ToL�{9��?W����7���/��k�:�<xUo)����0�T==;!U��M��o	j�)� �� �����~).�A��n�?p��������7��m!A=��2�o�Q��x�%0C�n;+k�6[�$�nd]�R"����M�5�{�������wpzB����R-���gJkTf��i͚o�ò�]q4W+f��Y	�D.�:DC���2~��g/����Q0?f{F��s��d�˳\B�@$�G��;�_I0��9�@��w4#�71�E�*��Q�U�q�g�OX+A��ڣ'��^k� ��}F���O[�zl��M�J5ɤ*���㼚r�ޙ��TQ<�9"`�5��*����)"2�G_p�ɚϝ��p�8m;�]�ŵ>���8GǙp=#�����,�8d��ss�gԱ����A�N)���v*�[��V؛T{oj�Μ�.���*����߳�P��Iݰ��XE��j�����d+�@���G��p403�`]���GI��,��9�.��ua�K's|r|� @Z�@\#�{t�ĊE;:�J޹�dW�����0!E�[Q'˝n�JRITU �Y!w!�eG�v�,�i��<����ɴ(s�"�J�hz2�D��12T�b��;70�����}H�'�m�=~�ؼ�(N�R|^J^��W�呆���p̶����ţ~uR,l�6���d����y�'Q|��_�l}�w&��s�#&P?W*�3�!�g��]3g���~R8�m͖��թ���i��0Ek��)�0�s0��:��hC�, �ay�Ge��V��<�
��G^��1�i��9�Z�@&��]��g*|������_Z4H�ϼI�W���u���ȍ�p�gVl�6ť�*�ϭ�a]�n��C���sA¦(���*w�n���-l�h�I7b��$~�)御�������+گ���d\����|�Ŋԥ��C�l���:$u�7����}?���/r^�QE0*�r��5XK
Z4
��$L�����X��f���X6�\�f�_�6~=D�ap�>K���������~�"�lԝU-5=�����+Z�%"�ޔ��sTq�ۊ�w-��Ņ��*2���k�/�=�8�� evQ_ͭ]�l>�ڵ^Ջ�T���_�p!�g�O
���d͞��[-�_��l�����?����O?�H��,��s��o�H��ܹ�Z�)�־HUz�+��2D�*���������� �~z-��t�"{L��(�M�jP��lo�lIdp���Z0H_ ��l�P�N8=��b7O�N�����2����N<7]L�`u�AEy:J�@�-���ڟ���E^���������7J�BM10��;�^�S]��p��`{��9+���|�fS@�튾 k��L��z7()�c<O�D�Iǵ���Ӭ	@
h����䘊�-�*PS��i&+?c��`�9��L)����7"�l����z�uQ)րS6��|ϷCs�|�}�R�{jcX/m�8�2�\JӝB�>[&�Ǿ�,�e��V�:OV?Ϭq� �[��`�ݔ}u�we}l	�t�o�X	
�����U5Mec�@X�=P�j�M�+[��M ��e���
�<�3��ql���H�����+bc ��E?�7��Q�Z<jÐӜp��R�㑓o�ۚC�7�]�{�wk�����}�Jm�D�
 �燾B-O|s�����ެ�+�g`��]��%d�N���.��2�4��Z�L:CɏHB8Ǎ�܄L�Er�(��ek�[�3�7�,����57� i;Fc�p�Y���I�]��b4[lNc��i�xeaC{��- ��r��٫���>���F��d�^w�Y,����bqT��h�2\�^�(�?���$��y���?��������֗��c/�)���g�y��	I�������_�\�<#ѭ�p3W�h�Ƀڐ�=�����^Ё;ݤ�v�6¸�x�v�Ԭ�=+���F�:$�L;4�L/��<����Z��cS���5c�Wk4J��c/���;I�z��<�U1��?����_[?�aLͻ~�Q�=��s�.��R���kY< �5��t���$G��mU�Ƴ�]\o�H͵<������R�j�m��N�5'�=�j�݁MDW�hW��cv��V��l���~���_\�<��f��X��Z�*���Q�Z�^�iu��h��	F�i�h<WR�%y���wl��lV��l5��sfS~�x�s 0���ׯ��� a�N2,��������,ɘձ,s_l�2;U~�YmR?��b��"�;��Sf\���,Ӏ���ͻw�ͨ]��O�*"�5�ّ�>]ק��M���ZZ�jzb���8����"�R��wk�PiD����D�v0,��g,VZ���/��B���Μ���/�-�|=�����nHY��#*C��n�4�����dB4��ܗg�!;	s�q�~I�!���D
઀:��������7W��?(� �+����v�VBԉ��^LQL���	�^gm�4�51�Z*��������W@���Xe
��g��,�E�B����?�c�p��ZCL{�f��cW���'�vv;�ۮ��Z�\��g�k:�Y[��D ��r"�X�m�Ѹ�?Wb�z�^j���Նy-�ǎ��ΆE�t���د��������!v�ǥ��쵶n�ym���Z��:/�g&��hA���(S�:du!`�M̖v3� ��y;3�����6	����k9��o�w -{y�&�$��Q%�%��l��L��{d�D� �4C���{�ı�`�P�w~?ձwG��H�Vog��ŜϠ6�g����2[��:|��~���y�3�Yluw����at��p���g���F؊hdO���k ����H8�>m�?��~ƻ��v˩���q
�'�:�i4��Ѱ\ύ� �Y�%��y:�� �V��7F�L����Vx#ƽ}���z�%@�3'�����Iu0j�����b�{�e�oZ�<sr@]zvPn�G3�n�s\W�,!����	�9mY/�}]��OJ�5��e���@�Z�/��I�ߌ�$�6ś'R�h��6�	�(��8��N�Zg�c#�kܩG��)��v��	 <|���h�#���9�g㞇�
'����"���C��&l�8��-��Ю��{���||��R�yf�ú��W&k��0D���1ƿ;��KuV<H�$��9�۹�ɟ;~�
��Bb9�m����F�;��v��8mI�X��8��ȷ��\A�FX�́��iW�&Ev��R�gc����G^{n�sx{{g=���Z�<>k�P�� �x/w�3o��uO*��f�ww�,��Л�ɮm�rpo5�ڌ��Jݚ͈���A�z����nF��� ��rQ�,*Ou�I}#=����^�9==���c�mW徆�|_ ��n�v�3�0����O����;�Q����d]�u�cS�1+�c#a���:��-���?|�T�����h�#+�{����k<+��'��Y��2�<w5�HȺg�p��i���'O��wh�qp$���d��TY<, ���Gc�M�g�D"`��A�P���e==����/ 3��	k�F�KxR�����*|]Ɉ��_�}�Y��GreX�m7�B�du�RcK̯�^�a�[��}������Sx-�[�G��/f�<&�c�g�+O!T��褨����|xm�.k���t&��g���f�=v)}a�} ��hpfd�U�����P`=ˌ/[7��Rt��"1�T�Y}���:��=�\iF_�¼�L4� 1c�����i1؄����& �S�j-�D2���h佯-7;���l���F�*G�"v]PD�bӁ�+�d����*�X�ĲX�/�֭Ԛc-٩��:�����A���5W���Y�b���׀0��6�}��M��h���H}�7 +��g�R�Y�u{NR<�m����"�s�ID$5#��f,���cU{��}���dͣ]�F���ňK��R� $[@�&�����ψ�����%׈M\k8)�H������PK��hr�h��%�+��e��Op�hM4�s��Z���㽰��p�N|������{vɒ$ׁ�)K�z�Ո�$8\�=���������E���{���#�^O�  �;_eeeF�4�k�Z�7�dՊa�qk��^�if��a�&c���P�z�Dk�u)"�!����BA��[����F�Te�q�W��^��� HN9T$����u=�`�y��s�w�x/�Wq�|%�066`Z���n�����j�F�]9�������������Zd9��)V���0mX��#���a{�^~��$��D;���i=�ek�/~fM�a�i	�hh|	�i��6y�Ɂ暹F�YӍ�o�ę�@����z(����P0�4Ѡ�:#����|��R�ې�����G������@>���	?�<N�(�ٷi�=%������;zĢ���5@~g��"mF-��i$�®��M�[��(�ͽ��>����L{�x��W��6�s�olOfS�~��] ʸes����� �޽�>ȏ?� Wח	�-�����gys�'�dY�,�>�������L�*��l?�q�zx:��<��t����D�PF���f}�3;�4��`�S������1����7Grqq��5��?�!�a.��Q:GƲ���AP����Q���3 �z��`�؞j�>)���[��KgJ��	�^_]�^��c�lX�n��%��.t"t���Qy_�q�4��5l�Pp]��D�C=��7}���� �D"A��fT0��ɍy��_X�2(0܏���hL�QCdGX�Z-�=�/�b��<;�$�<��jYy��렮*��$����*:5�5C��m̸.�5����$&Ѽ��� ��t�r���l�.��ʠ�O���n��Rs�w��R뽇�4V̫�c�{��B�l��l��Iρ�T�|P�$�ܷ�YDc,r��nX�1�cY��3���@!\Aaw2sEJ�Xϡ�X�	��k���&T=(&�F�21�q�>�����V��6_�Q=����`}��[��9��\�� ަ����s��n���X�E]�U�o�2|t�H�7K����h�\�=c�c{��I'FO$q4�yw�>O�-k�l�2/.�2�ɢ3���~L�y߈�C��\F{�;�pw������Tժj��l~)������_;4�ٗu��0{nP~�f��6+;P�:)䚚�ܼ��S����x�p@���lbTL�ӡ���z�k��C
��&'䂠K���[����p0F/}�_�@v����8�X8��X-���G�{�����Rs� ������d�����k�J>��Py�]8���+B���
�=��'YV�]�2N�]p�?�R_C�}(�Z��0̽q�_3������� dP�0x��iq�S��I��'�
���}sL���ь�q,�
vߠL�S�e�>Y%�pyy-�}�}w�Yޓ�����n��C�s�N���2��Ś$�����~5�֧�O�`!i��	s���m�s�b�:��Q�ײA4Q�����Aw���/T(��A���R����7r�qD��Q���@����O?ɧ� ?'�9S�k�uZGU�m�'�Z��3���E���" Vy�G \cu�N (�?@�]Q�v�pA�Rb
�K�����,PoJ#��H.^�o~�N�����ߦ�o.N�X�ό�Xt�O@i��;�?�»��C���`då![�WOOO�u#o��Uj�L>}z/?������q�Y[40~��͇�F��[�?t��U`���{{-�˜ʝ���eߣ���B��@�KjPe{$���"Sh|臞,�,����,�9��j�qKVE�##�?�=j{u4�N&�ز��H�۵'�Ғ*������[���b:���U�BN59,��#u�s��GD�D�ک�=z~UG޷Yn�}��j�pcaSGU�~��B7?ߠ�L#u��^�"��z;-��H{�-�J�L	�k4q��.	��*U��%��hnx!evk�}�ejH$�#����6�h9� �.�mzo�^l���>��u��k��6k�_�65�V�|!Q>�f�Z61�벘o*�p����Ҋ`[�-%�jG��͝���h�g,����U
�^���2�+���V,���9X�ףΊ�y.�W`�wq�W���*?m{т� H��:* �xG�v6�y�p&��帔�]6E���V���^�ԝ�7�歾>�Y���A�a�mshÜ��p��l��J���f�!RP�{b�6�<�}&=r
�e�5�,�8�Ep��V#�PS&�j�w����h�����
���t�UبB�Q5��F���|�y�A7 @��G�iB��=�*ܮ�5�N���N4�^��b��I���Om�"�r^Ы1�P�dr�: �N�aZ"3T+�8GC8���ԛA�8R�����y�x)�O�z*����~-w��.xO�t�]���Q�{x�n���	�o�M����K#���5��7��������,�n�aM�
m��#�ðj��s�_��jP\����a���5�>�I�X1�m����,eM�HC±��>�FV����:玒4�͈�5����|�iԵ
��Cͻ9��s(ӆZ���F��wy�	s��s���ó�n&K��J�{D#�T�,�,i�3��Ԛ'e?��䕌QȔ�ǲߎ�pOi��x�6����jfX���g�Ʊ��Ψ��bp����?���Te��.2��BF�D���A�̓����Ꞓ��iN}cO���W��Sրl���$�e�b�^�˓�,;RD%� >���H�d�)5a���⨕/���n>��Ҿ�tk�d����7�K`�i����Õ|��`h���/���y��AD�M��*��~-�ܶl'���#����\���PB��@�$)�(�~vr��rƁ]&/ �2��vq+��#��r@�d��gg"�{�̔�k��D�E�M�Ԏ��,t��@w�H�ZN��Y�
���EyLJ׏W���㍬�	T��2> �&j���S��y��A����r�X�f�g.�."��*��9��a;m�X���� ��0��0g.���W�y�=�����s����_����������w�ͯ.�w{���\9f��&d���=g�C� �7=&�O\@Ο�>��7�ҭۤ��rz�ʫ����9�o��&�m��2W����J&���x�����xȚ��d��p��(�c�����D+�ϵQ#n(q���3P&j$�h:�I�5M6�#�N^Wvo�W�U6J����9��t�N��a��)Y,C�\���f7O{2��}����������O�wL�K�zJ�5�:=/���e�p��^��!*�;fT�{X��H���Y���X�,4<��q�a����.�õ<<���cZ����_<�������B��2��Vqw3�C4g�N=:��219|,Z8���H��Gc Q/
����xp�gG���Cw�#�(n�S����_2��2·q�O���/U~�)6�4���w�t=q(4l�+�>fv�����0*�E#e�D�2R���'�k�4����,Y�/&β$w�߯�!�;��1V�ە��|?�kq���$�0�yr�c��e�@V�L�u(^NS���Ub����;�k8^������Kv�Js�j+��1��s�r��u��J�߈y?x�r<�t���;\���h5�՗�LU�$W}	e���֦����5��{�3�<!ፆ󕰝�3owa"Ł�v�rYX�{��I�/�P���3,Q�xxUp���eXZaA||L��ݝ<>=�y:<%�D���R9���:o1�����*r������k�Ƥ�w�<���(�lD@1�Ő�h!V���z��+�����,R$�S.*Y�H���?RG,��a�()��g���G��;e��K%)\�� c �Y+��ђ@V��՚FѨ��2W�!���Y��d$��?����́���XG���%�
��'��3�v�[�5	2�qPJ�8�T=�ai8cA��	X�I��.��>�i9䭑LA��`4��&)z�Ղa�0�b_�!)���̩����H���Vn���X���ͽ�(i�Xm������XE��5�:`�>#z
���*���l�7ب&o�@����e�+�'k�������n)r�@� �ԗUR$�Ifд�A1��
�y��<�-R{`.4��ʰ�W�2�b�)�N:͇�;�2���e�f��$ܓ�s������L�������N>���D4�v4,DK���IY3�^hЎ�1�5޾��o��R~��o��涏����}iMm����Z�S��іƛڨ�J�����a\k&\w�?lR�^���u <3��Z��Ox�	H=X,������,��O?2��	-��1�����zNi���u����}}/;��?���X��"���\E��pb,pf d��	M�X]�)�[OX8{�\8�*'YĚj��1��Z�q�� !��|1M�u�ɺj�_�Z��*��^BYѓZ/uCQ���0Ya��2�췞��@�s'�7�Ck��6�.�z�x�$��7�>��]
 �+!�ui:
��t�kڡ��E��a�r�b����x�+?�|�`��>�aط9�6�:UKuŚU)�~�BibA^~S�K(�ޛV%Sܩ�Xa�h�'H(e�B4�F�w�Ӷ�?��x��rc*厀���f4�l�U�6>�l�YMY���"����a���U�*{�=T�&Pպ&U��L�J��C��C�ߒa��ئ�ƍ�'���
�ʂ��yT���	Ӷ8�k�h�A���>Ժ��=��J0�U����~��������2�Ny�D;����B*��0ǘ���5Ro����qXkNVk^:�^�5��5�����G��sP/r�k-�����8�u+۠d�G��-��{&�����_��Bf�y��|�e`��j8�UP��x�fH�I����c�{�o�jͩ��Z�͚LVL����h��M:+)����u�4�ۓ�=f���Xy�����d(�������!(�E={��4Eb�>�G�x�60�@oD-;M�=5�&�YRz��Y���	�N/V�,6�{<S���j����#�ܘ��Ł��Hhh��sn4�>�~^Y5��
$۝Fꔼ�rj9͵��w��@(0)�#C��7KJ��ɉ����L�VҊ�z HMo�3*��td��b:�	�Mh��M�
{N���@���#Î��,�kG�x'f$�h-��4�!J���@��r4�7��%�V05b�}����1-���	,��X4 H�r���yR|/ ,�c5İ@�ab���ZSG,�h��W_�J��N��I��Aܓ�˳c� ��/�J9ˌ�y�^��atv._}�N~���"���ޥ1=M�="c�O?�(�^n.e�|�w^�Q{�c�] �#�ـ��&����w<��>L��b�"�Cb��?����5��7�b �CdD؞�7�Q��FI��~Hҥ)ff��߻x��JL k)�g�H��T�ʺ'J6�W}����Ϯ@g�z��Ld���.��d��������)�,�J�e�< �����  
}�f%ќf-����i-���ŝ�K�p}�{��i���ؗ=���i�W<�g�'��5�	��P��߂�c[	��(��H59��3-�/�0�}���F�NɨGK+ɏ,sg�/6���p	.&#
3�-X9�qC7+����C�D��g�2���w�6i�tʊ���8h������@+2i���{�x����Y��I5���:H���jomk��ht��GK6�uK��w|nj5��e5�����
~�Qd�i�g-��R��k�a��J��z���L �0��)��to��"z�BȞQ��w���T�ԁ�)����Ӵdo��`��벐*JuVW0U����{38U}v�U@�3��2�_u{�>	���U���� �Jm�w6*\꿘W��0�`ޫ�I�����s��Ǽ�Q�Cɡ�u冐�8#����ӳۨɍ����3�փ*XY��
��N����y�L}�5�L����z/?~�o�-�l�/�E��y�].7��]�2��QQ����?|4�Q�{ F�����R�Z<&�fE� ���Y�:,�NMM���jg񠏵�]-���[&籦�"��D���Og���O���S��u�\C�8X�޵0b��{EalX������=	H
P�kZ�^��͕��w��z�֯��|/2�|h1��&?u,�� �V�K�6W�^k��C��k*�5���ԉFkoƨ��D �@�<��Ue�I<{���o���^ߥ}>�ER ���Z6D�P��t�@k�'�z,g�G�љ'�=Z"
`h��}��9���B��)D$x��/� �j��m����@��`/�ZW�Ր������.��b��e����q����C��˯��w�^��z�z��r$g	d�:N@3��P���V�>*�5�r���Ǖ���R}��$K@� ��Z7f��Diӡ`G�����];9:��o����{��39??����i/77��� �����5�2p5z�&%LiS{�A��2�b0�kޒћ���`��>�|t�m���YZ�Q`'  c��n��t,�w�c�� {z��&̟cI[����m���^z3d��8�S����2i[z����8+}��vʡU�@��g�+���.�o����w����,��A��It*OV��6i�x��2dN�e$G>�����0��l��ԅ���{�u�J�ƀ�3��2�\��ڜ*R<\�g<X�$��A_)Q�OnM���)�x�T��5�Iw�`���LP9�5�����3Z`���SC�*q��tU�G�וk$�񜰟Tr�B}c{"�{� ���$c���uccYY��u��Lc!;I(v-Y�4^TA��	����5�j��*:��sn�(�uy��	�(Y��	����9��\�gm���+~^�������m	�6�{Y�����%T��?�>�J�����z$,
kX�T-�/��|��E)\Q,��@sԤ烮��{h�d�W]��tJP�+��W�fj�/<|d�����e��9K����91R�Ɣ����'��/+������8\ �g!Z��
`�N�I����"����@����3ZE������Y�P9�vF���~ƃ�xP
�O �����^�G�aT�ω�"CPi���B���Ƹ�p��E�]7DTb򸘂���K�d�mRv��p+������(ch�e�Q��ɞƼ�=��[��d42B��|sH�&�jΞ)��f>W/��3�c�?׊<�v��fE��Ai���k<"�8��qt��$C
��"W��i3�{'���_d�k�B�V�`jh|��;��m�ˤTo����0rR��d:pI@�ѭ�kxOj9+:����s9NO��AV���I�ۛ�o�?����������k6-X�
`LC� N�g$�8?;���T��^�o����^��ޱsN��-��n�тl�����崵�f|�˧�� �r _
:��h�(딂2}Z.7��Ӎ\��Q!�q���	$ _���/�x'�߼�?$�Y.e������Zޤ���0cn<J����H��ۥ���VF�O�L��(��{#��:�a������0VG��[�z@O����d.�|������;yu>a�M�݆9�����_>1Dp� � 0����<�Qt�埂�vİn�>(Ad����g~h��v��\�+�
ҽ�62��|�9�0I����󮎏�i~&2M�7���~GX����\~����dR�bt�re���5��Ѣ�	��jD������)��Q��)(�s�XL'�|S=o��<&�$�R?'46�5% x��Q��	��f�2mS�'��5�+�۫�S}X�
�}����[��Pi8!�Ź�{e���AG�����G�!��\,.�p���\W�A�~�ĻJi4>K3\�Ƕ��v �� b�k\1� ]��9H0	P���::�0���B<S�� ������M�Pe�<����Z7/Ԑ���wa̰��N%����7&��X�~�D�\Y۞M��L�k?������Sj�L|`LQ��2R0���-��`�4��Fr7�/C�"�s|�W������<����ǮR�L��m]y?b�->�o4>G��J������Qj��k�؋���"�Z2�Cs�B��T�\*úQ�w��z`m)K����B��m|�Q��S#8��o�h�?1�W�Ѡ��gJ�����P�9}��2���%�g"�	��A���&{��e�Z�`��Y75�B��
���52Ku5�Qg�vLC�<~�C����#^��'�?ؾ�+Zf4c����[�1����4)�٘�#� ��mv�%妏u+Wt�ZیN���s<^�|�^y�&;�O����6)(��
��Q���ljn����CI��X��j�l%'3�b��a�A`d>�W;�����2�X�����=�:%d��� K��cR�"�«�I����O��+��5LT�(m#���f�����/Ƀr�_��3*�!�Yٱ]� @�S�wa�,ӛ�[��Z�M#O����#��`r
v"����˫�9{�J&�#l�J���3���'i�_�]K�́Z����x>���S99J���DNX�B	�է����&�������X�A�@B�^k�\!�� ��Tka��S�	��=$��(�t�	��O���kh����Y+ƞ��ܟۤ����G�:�Ӟ���r|t�{�����9uJ��e,��E����C�h��0T��S��r� �� �H�͂�
�X3������:ͽF4AO<M�%���A6�4���(��4�g����1k�����mMn��M %��i9�c����C�ϧh���G��q�k�.1酞L�U��J�'���i��}�_}%�/X�+�������R���#=��g��ka����a�����S������Ԟ�ݑt)*{54F�=V�> pz��\��K��dG�o8�I*/��h�l���]�3�(z9�P�.k~D����''�;R��3�9�~�
��TkP5Z���یJ��A� * ��Ъ��{m�v�8>����[ZnJ���JE8㡒�)(�\��sp�Z�s�uؠg�=0��F̛�	��� e��	������%�,��y�Δ�>��U~��ؗ���łoy`�f!;��?��X��8*��Y
�-V7\�
�pw���$�?))�g�,��.*�&�o��]��/ K�W�kb/����0+7�3�eJy�و�����,E�Dܙ������5�B#�����ӣ�9��ٷ����b}=��*'�&ThZ*�g1Xڋ�C��Y�N�C_���x�o�V�Z�ý�(|8f�B��p��zԆ�C/w��P�7P�۵q�z����K�	1?�5�Rċ�r����G�ڝ݂�u����+��K�S�3WD���R�S��d��rz���Ԯ�7�[�'�(��&�U��5���}g�DAs��Y�-$�B�WG�k;���Y�{Z����?�#k�̎fr܎�1��<�qQk�dW�a�AY�C9����y~���fr380L�1)���y��'*�Z4�	��1��U��݆���jI��E� e����
�_� W>�\9��.��a�,9?�����A͟�/��5}d��g9����Z��i�&��r�&����F3�G#x"���5U���$�g:��-ʐ���i4�W����޾�[`-��d1�U
#�57���`���%߲v�/(�s(�� Yo��$���1r����{�.P�W�/�,��k	C����<xg�����G���ݠ@m��O*�؞���"9��
!T�ѧռT|���RVoi/�':v
�x~F�i6hs-����� `�M��,�o^�K�$�8>>K��1�
/ ����َh�-_S�����g��q���B�����YS�7G�N�x0ڄ"�#*��o)V:�p3�G����ǬJ0r��^%y}BP�Z�7���P���b�"�܃�����g"%�Co.�X� �yO���% ��Ǐ���^�>�~(~@Β���G�B�I,.�|��������@�>-���,{�c�TAꎁ������I���iP�{&j>l�w�=fG�pg�Cyk`q(K���>&zG6�uI�#�y���>J�dc�v;b�=滟��`�;l�1�3򭐃�{5FD��!��s�f��<�~�ެ�;��,���EoI?�/��7�Ku�X�Jc)
b�J�"�3���G^U:[�_R�����r���������� u�i�1L<6:Ыc��l82zd�:Ҕ�u�L��Ǻ	�<r1O^�N�z\ko>Z��yp�"���=�����Rɒ�;h,n���ٴ�S�j	�di�� ��!�j��W��݂"��#�מ�]���i(U�y�Vot��k�#SP=_N�!Vĵ׶�`�����2h�Y�cp՟�xs줮��+6+��AD��,/)op�g�UDr��^����u��1�T�����
B�a1�9=��byǸWqxN,1����E��vą��n>�t�wQV��Sb�Z=�ҟx8�
!��^ת�ƪ�?w���HV)C	��P�:$�"r�1�G�c��Ɡ[�`�o��>:�����nJ��*J�
d{����� i)��#-҉뀹�O�==���lF��uzz*�'�L<7��,�ю����:Gݖ�?������w_^01~2�Qy(�.yϸl�	+sg�A��#�+�|�͝XiXzb�
�Ý�\_���me造����r�D���Z���l����k_��T�z�c^�zf��c��%�`ya��_��%����������s�s �c)��&�Ɇ^��!�k�Q��=ʇ��$�e��sۣ|�F����Ϸ�s��z!@!Jƈq��	�{������5��z��(`��|,�{Y�A��+���P=��,
��숄��w$�N��Ę���	"' �w(8�$Y2&��g�S4���ig� 툦$���Pdo��f�8�"g2�ڇ�ȥ���o`l`@�ӓ�ř��.5�vX�vJ�C0*A^� >�Esgf�eԨC0�	F��#�`�tY)�`.����<z7�u�$1X��+r������H�� �� s�^ш�hy�hc|�g��K;�m�caX$�����rz�f�>���o�0Jj�HV���V�Қy��ׯ���u Y�|�����OW�';?U��W_-_|���J)n� ��V��W�7������;�8�����|�tGO�(,xl�>���2�z?~�$�;���h����� �C����:gݰ�x]��oL�Eux�b3��%gg�G�d���þ���6�ZAp5�r��Fn��w�c �b�5��j�����S4�u�-�/�R%*�>��T�Ò��@�8
1�Ө�(����de�ʗ�5���ڞQ�;!�8&�C-<�Y� ���+ �1��F�샩a,�1����$��8���jlU'���/�]�S�*A�'��5Ȓ2F�q-�)����	�9��3к4e��HO�Dkd�ᦗL�7Qť.��Zr�hQ>/�G���h�����/����!����c@�9s�G'^-பW�BY��~o,N�R�Ǭ��Qr�hu�Zz��uwF���=�y}: ��7fe�=쉇��G�[gd#ѭ�ʤVX�`i���89ȳ��lr[@Vp�� �d_��"y�*$��j���1������*){V]�����2�v�!U���]1� ��f�(�6�Q\��aƕ'�p�R#���ǝ����-��>�'n���K�6�PCE�5ގ
�~c�)X#�׀�2��5�h��i��I������׌��9�CL�P��յ���I~��7��_��ٹ#�G�BX4��-�j�����?U&���>{�)��=XA�lq���
����;�������Aq1�����m�� ��t�%%wI���p'ԥi���`�ͺmul��)�C?֋���Gm��։�=~�W�ޭ�����
�[4C�<���}ь�f�L{o-m7���`%�aa��zPy�L���?1��o-�F����l�v$�����L���֘���#�o�UfAҥw����T�K�I��1��n��#��5�x̢��u�h׃�עlF�F*(�:z��$P�х}[�5�̕Idt����_h��+{Z32"3\t;=/A���H�E�A���e\�</M�%+2�M��HI�?��J����#]O���C
��}�Kc�6!S�:�aoN�ѩwcЀ���W
a��nF�m��"�1��}oҪ՚��j4�Ԇ�r#�%B�P�,�Ó�t:[ߜްh�%�6O�pB1X���M-��0�Kk�2� ���$�'c/7�|�Y	=>�-�l㼾{Lkd�Ί1�Xk�浣�Oruw#�u���r	 uMV�h�����2 w���k詚ع��=�:)�(�E��}�.��`Ώ�̋�ά,�*��	~��;��}�]5�L���������!�, 
��h�>5��z�1j���(��wv���_�Wٰȫ�{�_ڧC=G*�� +O�uɺ�{�X��6�����*�U ���ˊpA�٥�H8�J��V�u� �m�jɬa�M0���� Kk.��`�V�`�Aw�o՜��GS%�-��~����[~A�}�̋��P����@ dEMF��Z���<s��,,�`��fMH�̮�G���ݪ}Ydq�<��4�(2g�qb�\Rj���.�h +�5	�l!�vP�A ��{>TΘ�W � �Y<�t`L����{ȣH��)�g�l-7���k�uS���㡟�H��5d�h���zb�XzH`*#�؁d�,$��Lo�'�v>�+��%j:����u�2M\��g�Ԭ���|�2DJ��T��}�j��+��Y���]��2�B;5��[�9���ql��a�%�j�x䣇
�'T`lokB=�m��j$����K �.-��_����h�����z}�C6K�`2{H���O����r}{#_|�s�#�1ךN]<xݻ= ��!~�(��RJ����9@L�x����9n���N6��8���D������=���uR��i�V����^e9�B<��D�X7�V��Ó�t������:��� �,�3f� G��G����:���Ѵ֘��ؠ�G�#d����vȫIj-,%�����g;c��V�y�<Q�YC��Mٮ�4��d���ub � �(Y�X�F9�<:'���`ax;����߿OJ;��N�͛S9N2�r�WEk���}�7��u[Z`m�gp��͑�e"�Sk�1�o��������X�X0O�������i��k ;�r��k�����D��cPe�ۛN��>Q?@�ℹ%�#G��i�1-(�k�P���~��X�S����rv~.g�@5JO�:a����$����i�$`Dnh�W�9��t�2�q2�indg:�7������X�Z �N� ��e�d4#��q�c�:־��i�D-��I��So�����W�:�ʌ������ˆa�;��gD���dƼ7�؇����'�O�o�\�~��&8g����N��2���j-���,�v���0lA�����G3-!����QG��nZ�T
�ߎFD8v�����$��K��������ܱ1|��ɘ@�����u�&����YL����XT�댝�����(/g�Tf�^?�~��V����E��\��Po�Y��dtYm	�"��J��x�;�Ԏ�F��Ieuê�-����ԏ�x(��k�@v�Ec�se!ZYA @:2� !|�Q����� ���=-0�����:�[��ڐ�f��PO
Q��!���YX��Mg~���PA�&m��V_綞�Ã�ژFtRB�g��~EM@���E$��Y�oo�I�37�"��� �Ӑ��AZm����21c]4� ��@�����%��%��}o��.*?H��ih=�DQ�G�`��z�t�Zi���|����	7���P��ƽ�~cnom�`���s{!dm�N�gfx��2�zX��m_�*��Lr_�h�Wl�ҏO�2>I::$���FS(�G�ux�����s5�`��ƪ�m�k�!��h�����0�R��ԍr'*� � -��$��������F�^�b톔GC�j���<b�|�%��AaJ����ێ�R1�Uz�Vci�Z6����������j�)�b�!�i��iR����c�� �%��	OOw�\<� �и�zQ�d�'�������4�w8�Qc��6) ��6��>ȗ�|/�_�!+ֱY#Uy@��<��H�!{��-Y=\����`I��zJjmLqǫ�D*[ht�5gskY��$W?�An�/�y���1KWt��i�xZ�P:�$���; K3��rq/�~��|��"��,�팊Q^V�Z6���iB~2TH�K�f��D�L��G��C��g���!&��S�,�W%�����>Cb�4)���!i��k�'=���#�
����(�l�0�>�lX��d�4CV�@�2��dY���r����]m�'�{?��dn��*� Hl���I�x%��KY��aƈ a�7>�QY�BR���'I	��r�� ����x��Q�~�S���N��S���^=�o��Z�������9N{Y������c�3�*˲�t�uG��N���w����$2�
�	�%��n�7�C{Y<���pN2�����@�	(���4��ӵ��m�t^���/�ի3�w�|���9C[��c�,�� ���T {�ў�1�,���C����s� l����i	�.V����å|� #�G��g��\�s��z�@g�޸�SO�;�{�c��W!���m����}J��!]��������ߧ���K�Hs�	C;�J�pW�Ñ��QМ��,0��Q��J����0R�C$����e��IZ?#��mǒX��������|H��kR�dJ�k/�٧%ϗ~�:�>�J���	�p�����;�:�>���Cc�3Y�b(�(����喞]0mB�@ݠ���w��E�pGj��]j�4�JuШce~����b:B�3�qE�S���Ϡ8x֘#c*c��E���^��⌢�6����*Y�}�4E��x�p�ʮ��>Oل�2B (F1i�o�Z�9C��&�7r�,�jM�:���2EWD�ZFe��f�!<�d��Ж�\h��,� �=��9,A��d����Ԟ,kB-�eGo�J��
{���m�W�Le��;�\���Ў5!3��,VǑ4�lO����d�h�i$�fE=Rm/:��1���`��[��m��-/���g�V%��UFB�3T��4<Ӂ�Ȫ۷7�U�l���%E���N�-�@��Hm׾|/:��x� >�!��2�ޥ=<,��B�9b���>9��QC.ԫ��%�g�G���Oge]J�Y��|�z���^��s�����C��nL���D�ޢ�E�{�Z��DP���t��P�r��,����y��f�
�l`���'YC��^�Qs����IO9#QC=�� I%�~_%E��q)����?� o/^�l2�//.Ȭ���[��u`J9�*�^�Q�,�U��f�\�K���ZQxQi��֍-qOF����Or{�))��M��>�M)�<�s�/2��v��?=0��/~�[���V�ŉCc�AZ�c���vU�����j���/��g�����P���^�{�FqK��ɘ@�zU�A�Yx,�S�O�DMhh��Ы���;.���`bƗ>C�� d���@�$z=K���>��#�
m��\,(�0 �[5nԣ�F`��Qyt�K͙a�Lg��x�;>e�5�������#�2\]]��	]�}��!o�>�{)���Ч���;y���܀8?9�S2���^�W��R���O1G6�=C��Y��L��p�?��b�G���E�Tj0�}�wU�g��A=-Х�8�"�0f ���tnd ��������K��j��ʫ$�޼���u���V���������t}�~����VsZ����%i�8g��'AGd�1z�1��f�?<��?�(�G��b��뱜��bN/�dŵ�S�J> ���۵XƣZXn40`�����H��L��1��6��n��q��������_���Γ.;���ݧ�#���Qc��J]���,�T�U�ҁG1�����z�Gj  ��L�g�P:�k4:�v�P�T^��J�ZO)����$R�"3�f�*��r$������v�)+��&dpϒ��M������I*�ꖍ�y{�z�ٸ_]'XJ��M���1�0:?#�/��U�H2x����k����R����sQ���>�V/��C�љ%��|�>�����m���AV5de +�L��G�mAٙ�����刪Vh,�<=[�c��'��埠*L=�w�0��j����vd����z�]}sH�Ƣy��a(��1�;Z��CX��X�o���dC �ʭyC��Lx�Β��ѫW�59�1Ss:w�{B�3�Y��u_��(�Ȗi�co�jP�ﻸ��`LpՎO��;��
��F�Z(B���Z u�>��}���e�>{��@�.�b����=8�
�T�?Ǽ�F�J�BSR>[���ʲ�����!�����ُ��s�������x�گe=�A������LPj�PC6*KX�=��
�f�3?=����Q����Xv����I���>���Q�A�����[���[99>V�x4c�#���[I�_j��%�0G6�Q���!�)�F��mR��t��=	/@��1Tu�ZV��J�����7KU�4x|�';�SRzQgJmE���l��Wh���z���?\~�1.�/e�����մ��$�x�smŦ��j���@$!����2I k�r� A u0_!��<CIk����Z^�(�Ԓ,+��L�S��I֋%�= �6�-����Ez<�86�e�$;f��fC��@�2��eRV�PO쁹D
� �9k==.	�v`i�mx2����,�#��u~rF��iGP���B�7��>�=�9��%*����An0!K�\��5<�`1omϜ���>]ݱ�0��jo��N�Ӡ	��A�	�Q �	p�;��K$��#���uYwi��,*<�p-''XGaz�{`�O�@xd�V����h��|5V�9�Q�
���!t���E�l����+��#�����o~�M�cQ����bF��#X�SB��/`�enb�3ʹޤ�}
�j�,�nQ���3u|���F�JC��w2���c����rys#wi�m-���D��&T[ɜ �gM�1�-�fyBQۡ�u-�4�>Xy��92D��5j�vc
Ec$T�6�����a ����z������|�2��u�"��F�����d;��:CE� ���58*z����Z����D�^�xf�U}�ڥ�E57�T���7i�G���F�ߠaV�
A��q�^�P&7�h��ZI4�L�z)t�1+�,3����N
s�)OA�u8I;\)S�%���&%	�o�z�$HV�Ռ+��&�»bQ�<.`���U�eNJ,Jl_y�
�k}���¦�Ձ�(8&�Q�ɼX����Cs�%�e�)kC��ڃ�Y�UO�g�*ZM+�����k������ d�^��ܒ��0��v���+��yYM�j�Gi=�S@����l��;)!Lk�F}��H�5�o�b0�]'Ŋ�ݏ/�5�w��>�Q{���X	�X�<��h��yͅj߄"$k[R��\P��!�;��`3;�1�g1�r���!�[�&���)_�cdy�b �[��QgV��dJj�)tP� (�x��jp_]-^�����\]��?NZ�FBj嵐��^�1�O�=���}���E�á\|z,4,�}QY+z�7n�{�Vw���-�t>]�C�<�>���u�'j�b��q*}�r,�yhf�h�ہ� ���yR$�R?��T����e��g@+�����/�8��,��G'~���%Ca��dm�J9�`��D5�� 8�8&�a�&تnWOOu��,�냴W���B㠇���Y�2�р�:���K��jϺYA�&�v](��� YC2���.*�Y�
S�p��a{`��W��� s�-����\kH=>>I�^�N��J�ms��Qa����	Ev�҃;��-D^s�>��O :�4����Eҋ�I�-)��K�'�_ǱQ�4=�c�1��
�x[��H�0�iօL�%P̻Ҍ�$c�щ� �K����"�
.�<l	ܠP�i��d)-���x���ӰR���ݫ�V�+p\��7�s4�|
������ �Bw�e�"�@#OOVo�e�o����I����� �2�	��EM㱮V�
��Ҕ��zIY��w�3M�Q�U�_!'���Vn���Op4�E%��9⥅��A#.2Sft���oX��H��4CI6�$�
�zY ߙqX˶(�C�1d7�95r]�X>[�|�|�3re�1`����5�_]S� ,���J'��(�͇��秗�%׉�v>�J�E1ÌEtl�s@ϲT#'�Q ���q�2��C.����#Q�W;I/�DB���m%|���� ��E��b�Y0[�
��
eJ,��z"�

��^C�k�.�:�����}S&v 4�T+��=%���0]^$��:��z��luNޥ�e�m��zo�?~��"�z*�H�Es��hy*���r豫�R�^� 찊Uݭ�qׅ���b�y%�V����T �>���钷�}����tM?k�	^�ږ5�a���Ê�{Q�Xh�IQQ����!�چ-B�	%t����\Qn𙁩��Ց�on���1�UB}/W/@�h��w�����G^hq��U��A���l:���J!�#+`��Yإ/�vS���������˄.¦��;qr*'ǙK����ǧ'z�������D�%z昱�QA�c�ɧ��|�x#S(Z�F�G(���$���v��Z12:R�����ZݣYO)/���k�\�O�W�JQ�n+���m��+���r�ӏ� �&���AA�Ӈ�tDj+�e[��{�?�8���Z��u?~�Qf�G����D���hU%;XA 1׋��O/�?��_�[%|�*#bQ͋#B��IY�W�!)���� �G��uR�7+M�'�k�"P�sm�M&�����h�9hC�T��� K�൪x�&�P&�f�G^��d�B�����}z~d遮�0G��-��Q���ހ9@�Q/3f�Ѥ��Ë�5��2ax��A�Z���7̉M8d:��~��t���d�-��d{O�,�e��z��G�B�A������3⼂�|����6�Ol��K���v��j��8a@��Ϧ�{�QBX(J+`����������ҲfӔCL��!�P2���ʖm�FJ��h��@Ly7jC�QС3��H��{<�џy��Wgȕb�$c@�q�~�Mߙ��N`��z[dzt:��g!_���0��k��#�$+C�����#�z�F"�=�!q.	o ��цm�\8P���-jсq;(��v�f��$����rpݠ�gpc��X��]������T/w��:+^�kx�~�<b)��+���"]�-��~�l 0LN���z������E��T}Đ#�>�p�&;����ϝ�5G���}5�B��x���i>�As�+-��r*�F�_�2˻50�����sS�-�)/z�|��l͚�kzᮽQ6ƾX�5���I]�~;����
�L���Dπ��`�?��kI��K�t�� ��+��r�nw��S��0�׌ʚp���@+�f ��}(o��bȎ
�D��=d���4��]�Ԡ��J[wb�"�G�WW���<r�	�[�?��u�4!�H=����lK�X�{��N�a��(�ZQKkd�;���Ƭr*�bUʔ��^p�^p��ϏO�l^��
�_������}�ha���O����U��	Xe�8�J���hD2��������1ꪜ��,w�o���N~�(���1�3�"'�]P~�`���ф��P��Ia��NW�.��Z��1�V����I���������$�]���<)�����_������t��
-���#���i$d�k�f���{�22j	���()a��Gy��N����d���Ǐ��O}��;W֜ib�w�	�d�2f׆�$� Zz���O�Y��ݛw�+�˴��((ӗ��=qQ�pd�%�>(���1x����C% �P��.e��g�H�I9���lX��Kk-���Ձ�ڜ�}݃��K4�gkAC
�Ӗ�Y �C�ֽ���)8�SI<bS�ŭ�\�����o/�x�v��[���=����!ȁ�p0�1�&:�PP6�`FSx��Q$�Vhy�&�u�}�[$;��u\��Z��F�R�VB(��Y��C5���9�q;M����[eDM'��!����u.�,�M��cӏ��b��Y8}ƐA>��-d^���m�d��'���	�0Q�=r{:%�����i���3�y�ێy�0RAv�SwO�i�iabqR/Q��+)�=�%�@3�D;h�R-=Pf���#���_����,���+]&���EN���|�F�>�$���L���>h0��
����g�t��yQHР]����6��䀘�a��X�FZ�kE���h!�n<�����$���}�n�����b~q'ZC�ɷ���(�ޢ� �J��{Rk���Υs2Q��/������\�h^���𨑲�k���J-�nkMb^�9�tmp�a�9E�%)����T�T���(J��%�B���l���\ $&�b7��(���0
t$�y��M�+�x Z¸���[��gD���Z[Bs�8tF��(O�g��Xy�ie�e�	��nJ�u0yjas��#+�W���P]!߯b�z�g�:�$���b�k��Q�y����,�l�J���|��1�'[�?��#g��Fg��u��i�t�.H�M�M�{�U��%m�K�_�3��q|�s�)s�����d�7��\X��m�Y�wO�|L��6h���J��Q򁪞��+�{�L��6��@����ӱ�X�t��g�9{1����X_k�X��p�d�{˃�['�l> !jF�Fښ��aX!C�Iu�p�������Q #\�A�0�зr8x�,���L�c�s(2�i.�����
��P!�W_�Z@i0�M��"��������x<I�DI	���}.g'��@Hm��L��-�޽�bʨ.��y?M�pB�Aq�� 7Wrs�Q��Ox� �����B�D(&�1����	��j�v4>�`T��InT���-��ЬO�.,�=_#�5lD�p�B&[�>/1p�Q������޺y�!�)#�ޫ��4��Z>&���2H�
�S��2� D�����0���h~��h�_���57AB�(~N� ��)��g�Q��;�e.՜fD#�Yj�V�/?������CRr��X�!xZ���cڧȑY,��f��m�:L#T�5dh�_��dxr�d��j�b�lbe�Vj�u��v�&�
��3�O홐d!`�����]�^Աjӵ�@�z� �f($1��O{gQj���s��D��}0�s����vȓ�q���+�a��(?��v.�fB*x��-Uo�ŋ��E�ݎL�{���k�����=�*�4S�	�:(p�|z�{GH�`��׵V�!�2��FQ2�t41�5���t.��_����o�����L�[ 2X���2o�^У����vg��U�g2��pi��ͷ�@����!�Y���F	���8L?N��$��)��M��s�8�Wg�����$��M0J���b���$�b�x� ���k�uZ�)�|B��K��L���k����G����o���� +Gx�9Z�z�|�{��<xA�U�"��;MԞ	�|v��?Ti�Sn�������qP3:�wL��P(������+ �w�K�j\AV[�,osV�=T�S@���.��YS�|����,��9�/�l�#��C�D4�
�;��IeI4��N��u-�~W<6CI^��j��SR=%�p�O���j��y��{�%�l��1Z�j� ���%`�tj�3p(�^{��7gc���P+��o��?��ʵ�=�_�i_,yU?j�s V����ů=���7�A���.\5Tm=xfi?2�M��@��Ec��_���;� ��B �(@�k��g=�D��Bx���}˵��Ù�}���8�t�e��!�p2�M�����3�:+�;ˋ�<l��s�"kȴi}1TЍ ƺ���b43����+��=o�nw;���ek{����Q�9t��z8BRZe8��F��h29���0E3Z���X͞�����|��:D���=�zq'��g�廕��_0|I��dFO>kE@1��+/�̥&�]D��슁V�'y��%!���%Y�m�'
�.=潩���=6>C���F���GԶiJX��2��a=����t���S9;{#�T��F�}�fSGYL�e<����y���cEn���K��!�KO���6H"n��Bi�,���Ar'P�K�C\j^BdP���L�_u2?��"��a�־���B4�|+�<<��}c�\=V1b=Z�^@֜Z��]Z�W���G���1�����m�ߚ,ߴ]5A	�@�p0݁�`��1}	����y1vc��������im�=��N�fu ��NUqF_����T!v�9�5a���=�'���ab�YO]�z�4�Al�5v�FO@���������wV"�̢��Z�A=���9�.ʾ��1��pbӆ�!��z9 P�&ˉ�{����y����}�1*CZq��Ȋ�SY�v��n*�.�}�D�l� F	�R[v����1;?�ɯ��B�귿J�e"���� �4������� uJI
��so -����czs��6��I�bL|dP�L� ��M9���C�/��"�|6��Ԯ�E�#DE%���酼y�:�<��dJ�?�wJ��I\ҫ������K"jr�dz��(�+�zBc5
c� 9�ǝ�����(׃y��o�K>W]�IBy.�שʥJ���9e��Q�8)\��=#�0�]�1����Y���g�6`���W���נϯg�̟���N�
�Vg�d��������k�(+i�;�X��3;�bq�t�`��gi�+�d1�f��N
��1-Ȉ3��ZZh�R�P���A�@i{�p.
� � U�z1�I�\X�!u��WNLS V0䖙�*To5TZ}q���
��U����e��#��P*���4^��x�i�y%Wcr����˪�)Ѱ��	���|�:���_6���P(���ZT�30@o�7�������`bx��?��ԟ|�+�b�������Z�����܋�8D&ֳ!�q������h�ZϺZ�G7<����Z��P@y	��y��W��w� 8Y�pi�f����B��پ�Qͽ�>H��ʎ�jzU�<�|@͏F�?x>�vL��F����{c{BsO�(q��jb=x׃���� ��GY>��<���ݣ�~�V�_]��+�G� ��AC �666�~PZ(aT�&ݲ�rDHhq{��d��g=��f��d�k����e�b�:ދ���ېs�@+�2�����y�����㇤����S�*�(e�2���״K��ܽ��ܿ����=�`({R��Ƞ�nM�s���#�����Q%k^��%�2^A�5�16;���+tt�H�[/'��G��|ZR��¥`��t�'5ȲHj�A��Ń�ޡ��Ń�_����$Vyx�"�|�� �,�^7�W��Z����N����6�C��N�����]��] }@�G��4M�l�R����P��b�#P�'%u!���t��B�r�v 4P�I��BL==v�Ճ�Z8�r8RfT)$�{�x�����՚X�$æ�$?�Y�i#Y�z4YL�"�ᕞ���$�g	$�S�Hy�@�>ݿo��G�p;�O�{�ahZ�� <Ӹ�A��������#xv(�B&���`�y.�3�dP�y�9.�^k
R�E�X���/�O���4}΢���p���u�}��;Y�u�O�I���3dY�)��z��J;�����E[pʽ����܁�q۠ƖL���cF�$�o�d%��@�I������r�q�HI��B�� `|L;�� +�]&):�@!,�MG�4�3��A��y�{�C�h����Wrh``6�4�L.��LR��<���1��+'��M(za�/0��*�5��~ѵ��4P�9�9G�uJ�za�[J�t��I���>��@��S���W<*}.����� ��8uݙB٫%d:�P��Ua�Q���[<a׽g�&c���9���;@�'�}��R�V�gzq�)���a0AR&���j^�`���mP/UVX�f�I�WX�Rc��z䢟W>��r�m������y����m�D���2���[�k  ��IDATKT/ݮ�hno���N���a��D���֛1�e5�1+���G�[K�`[�o����4U�V�!�L;�{W�1����������*��{��E*oLo�AJ��{�]������)���i`��z�3��C�V����F�wu�B�D�kY ����j��yt@$��J�6���� ��s/�R @��f�d�ް��k���x�; ,~d��`�����Y���;�64
�`ؙ�54�)��#��(y	IK��!�;�������cؚ�����eRB&#Xp�'s�pǛOWr~�J^�y#o޽�Wk~���'d%���}��\��ڸN�\,�dAr��,o?�CW��LJv���{*�jȊT���z!����W�1ו��]%�=�C����[ �7[TT�/?��2?:����dFA7�Ho��֧���)��`���X����d�J���#�A8�#W�2pN�TF�{ �>��{\�׽C��&������ɉaGjn(��ݎ�K�WI�<O��,]�ѺZ��R�<���dp��gQ���g��� �-��ۻ+����eVO�����+)��^fr(��f�<���U���H<I2h�c�������|��~�~7����Bb\�i���'c-�Ke'���޵t_�'AW:�<�̩u��A\!�Z ���`}D�@��D����4��I�yu!5��f�V^�:fAb��@__H ��� �SQ< �h<��@�?A��XQ_�Z��/WY���9�����9n��w�	��W�,��V�iJ"� �Z*���z��8��7e�#=T;�>"�`f��X"BT՗����i-�9�i�����[�P4�Q��0��$�J$䆣������I�s;E�U3�9n���]��5��t�WIw:" �'B F���Ғ^Y������Ju�6bfxVU�0`[���!|�0�6*�m��<�a�d�zQ�P+�'
�L�iL����Q2�H���=�Ub�e�[�a���˦��k�/e��ɉ��6�*#'H>ڡB��M�p�S����)��˯.�.�|u������<ݦ�[�!~uL���U\�A�"�#2P[�*�%�\���r�z�c�:�l�A#7�Sk�4m��фL5}KĹ��@�Dq�3y7q�Xq�	���Q!f8G�n�7��[���:�4Ym��Z~�{�W��DFE$����j�����@���]W��zn0��7����
�s�F �U�ࡱi�%*T��;��պ�&{"ܫ��Y�$姹��� ��b[��h��~d 4b��;������eR�`̑ōm�],�ռ�[*r�`�:2�g��ݪ�ky��U}l��xK��q�PCT�;�0=ؘ{Ϯ-�p}��`� ٘�{Js ݡ���:�C�Ҩ���t��gJ�-�Ż�@�b�-՜��!��lmv�og��rk�G�#�l�2�,!���Л�,B�j<~owdXk:ô�@�I�Mj��7ov��� �������M�|ڑ�kE�a�Z!$n�f��P��P�a���+k�e��jŢ�8�a]!�"���lU�0��|��S.0<G���2e�8��^3aXq�t<t��?��FfHRFm������R�o&IA9���_%%�B�O������GV|tK=Q���e-��G���M׸M 9X����P&��G(.�ɘ!N��=P���%	�,�C�dYDC�p'���������2C��S'WI��%��t�}�d��w�dx��h$uB���ޅ,�F�]^���;Y�ρ�bn҇n�a�$�qt�1�ݧű�gg�w���w��$��Q��,n����dqw���yXc*�P�7�5����>�����7�-(פ%\��>��ټ������&�pF��5���!Zv�K��1Y���<�K���f��m�
�n����^]�f��wޞ��V�I^L�*3�y0�4&,LmEY���������I܍d���>�<�F�����u�&��@��3�y�$�r~>�����������WI~̵H��Q��S{R��(����D����,��6��܂Up��1gs���'F�J���T�؏���Ă���3�^ec��-	&��Q���W��w�����(�o?$�p��ւ��Gs5�@a��*�"�'0��������̪�7w�XГ?y���|��o�_}C��Ï�忏Z���mҵ�������8��i9̔`�gDt�m);j�D�<�8Ð��T�6���d6f��	�@۞��"��p�(��]A ���i`���z�j��e/ߔ2Y�{�ԲB4 g1�t���9�iM�#�uLr�I>�p-o�~h�S9>�y"iL���/�ne�F���'�����5$��k�FB������"�D�@?�f*�n�����c��鄀�kN"��u��Y#,����A>�$�{N=}(j�c�_З�L~}dO�zJ۸>,9���pV��G�SH�K��?�ES�^��_�v%�:u͝A`]�:��EZ�^9�2a<��IfP3�'�i�����	��7�*�=z�����t���u������{0���c�:,|JCl����
MÂ�Xb�U@�J!_h��'Ӓ�5���)���g�MWB�bn�5׬��DC�R-��_s����0t��!������ ���]?V����ߟ+����v5��1���*jo��[�c�C�Մ}'�g���7���n"��+�Y��$nU˥V7��uU���x�Uׯ������>�_����Q���u�%�×�����v{�Og��y������q����E�?���do`��������y�o�zo�V�z�V�u쿇�s����7+w��`�b5.�W
(���A�BP/S�B�J��T�ٚB�d�^s��s�k��E����u�h������j����BnPy}wG� &R]G� �P��Y���oZ�g` �z�ZJs�M�nߛ�JJ�rs�Z�'���i<�Yad��g?̧�Ӥ�"�%������-����j�LV�u]�Q(��Y��H�$����wfVVuW�|�3��}��/�����twY�~�N�������}��UL���  3SSQ��G��.C&�Ե�=�~CS�����ؕqb:%��F��7oа��.�)!��%lT׀I�������B���B�}?�+�������ۆ���!Ɛ]�I��������~ ި�C��~�Y,�AN�u����m]�n�(q���B�l=��qZ�od\ק�齠���ڊ�P�y����Z�Z�g{|~�ۇ���PqC�����Q����A0�UȂ��<b� t���T4=���^����QI4��?�&��eq�N����Wl|���?�zuΠ�3�k��,Ź>���K[w�bmFC�.�]e%Լ�c�yfC��-��!
��|�o���~�اϟ��Ǐv�U�=2��a�� ��wuy^ �+���r.X���ޞʽ�x��~`S��9 �N��;t@ۓ���X�w_���~�#;�=�o?��;��od����ҁ�+߁_W ��&f�HC�LYO�Ƃ��4M�L����ֹ��L�-X�qp���Jj���?[�l����LV@�)s�eP�L��z�8:�D`:8\c�Q������MS��gR��S�1܃�����?��O����iy}�Q�>//c�ȞJxIT^z%�j	z��Б�)&��38�2�7N��41�jK��E�#��+cVJ�*����is���ɘ<�C"=7fs�Vݝ�&����}N��69מ՚��#L����˞<�J!N�3cu՜.�t�Q����`NQ$���U��AE[Q��}*�4�p�q��_�݄p*ZJ���W���pXv��&@�E�w��c���Gl�������j�Xᴽ�z�夏N9�(f�,�1�������׎�k�-2?"^ϧ���&�� w>A�D=�}���;�tR��;��49��M�8������R �a��nk�r݃�KP��xt>��H���
�*��m��&���s���#�`O�j�@,� RA�{8�� ^>r+�H�2�׿�S.�P3a�ג��Ə�f�n�}�W��_Ԥ�<U4O��p�p��G���@�?�k�X�	>�^��(���I�h�x��j�@T�8S˖@Q��[�)�h���M�@JH���p���
0��7j�G�����n�#�,��)�]�>����H���3�lY$긖Х�i�U�XVfW,'�vRݤ9�W�B�tP�=h^h��m��Z����Ɋ]��E��d���(u��3TP�*�p�#�u"㔦p��T�>ٜ)83ͭ�8� ,WW�}��}�S���|bM��D0��cwj�39�jw���`��6�����G����F���[+vp5�P�{եl��ᡀ��o���>��I,J����hn��V��^�B�5=�Ɂ�Ư+f[/�
jP�<�dD�.pbc��]-�٫�oS ����>��h�gP�I�:)���.3��-RP��x�<�k��`S\��}�uW���i�Y'�W��:�K6�!��и�w�������?���}W���Y#x,@��g;87�u^���&�&I���˩��%��/#������`��?��9��F ��K���R����垬�5��j�$ծeFMT��b���'��!2f��=Z"����4��g�wۢ��]�����C��}������S�y���w����S�|ug��X�U���͙Y��[I��8�_؀=�k2a���`���V��]��'��Β���.0��,���H�Mڌ&�_�^�9�	�[f�Z(�%�	�F����DI��af ��_��?��&���3�Q�W���0�T��O;QCGm��F�����NG��%����S|�j�F`-b�}��t/m�}Z���`:����LY=JܻBnr:�b[���y��8
�F2Bo�,�!a߾e��a웕�/�Ws����p�������+�6$��o��¯n"�'�LZ����S�}'4Rz��-��;���9?{^L{�����! (!M���'Hu"���:��
ʩ��r@;:: �������Tk��*���<�"��j�8D]Ǭ�v~�{�������K։���+�z���w�;N|=v�	�U��_=��*S���?Ve�������oC
V�uX]C���ñ���HrR}Qf�^��Vl�ߊH��ݰ�<H��g�Y�n
����Vs�O+���U��
h��_����)�#0#/�~���1JS.NA	\oW?57�Z ��+�^�1>��V��-����Ͽx��L�+�[6�����8>��"[7��1Ò��eaѵ^o��٤ޣtR~J���Q=��ݦQ��g%�Π���W�Ĕ�6�<><�ͧ{�VT�����tuui�^����+"�>m5�ˍ��~�����Z���8zcQd���ڳ�F!A��� �ۺ�b�`|�8q"��N���5{����T��u�M��{�̠˦y��p6i�BѩmU�b�R[���L<d),R{8��2 �����..���}F���4Y�-uN��6M�Y�$<���w����=^d��5�:�4\�g<@5��^���"�Z& o6�ƾ٬)� ʽ���9e��1X��%|i@�"�-���0���������%�X蓴d��T��䬖V�>g;E�I�{�m�+Z����[�q��@�m�,w�,�iT�K��RY���5����6σ�;s��~ �Iw"!�N����A0�ʂ����®__�o��{����?����S�o�����0�ϋc{�L��:P5��L���k�jX�C?_I��Ye���Q�E�k�� ߅뭀$�Y]���[�;��ހ��������� _�Iy3,v~e�K�z�~���}#0���Usk��ݛW����,������/�������޽���W�p/��GR��	Df�g6h.�eݷ�S[4n��k����f����%ڰ������'��/�����B+��A]�օ� �V)[���g`��5��_��[?���1�{R��&��+�w�S6��u��_��V���|�T�}�z:�<�u}�e��^�I�ՙƛ
��O�\�5�#��b�����!s�;�ި�/�������=)]j?o,�����+�Ιu�ng���#�+{<g.}e����k3wE~��Շp0��5�w�Tg��#���Ҝ}�q=!��lVG@?�iU�O�Q�m�:��pL�,��}3W7����s�J'�ӗ���2N�\ܞh����	B��i�9s�&&P9�(�P��UMӽY1d����m��a��*$#gN�|Lr��x�o�́�hڝ~E'j�T�"��t�Z눾�\{����.��xq�- ��N�PQK5z�cLc� �g��oҢ�H&4Ef3�݁��)z-9}N/�	���X�9�S���b�x��%w�&�6E�}�g�k�p<x�!Q�����7�p�œ� ����N�h��Ѽ���<=��䀅q��<|�k'�an�r��ά������7�MtA;2rfV��1��O�W��M���`Fqgǜ��P��7�VΕl��R9�$z����@D��p�ksG��������Q=O����B(�|�����%�0]\\Pq������/X�L
�S���Y�*��8:��3�N�I�&ke�O|��u��x�����ϫE癶�-pK�Y���RX-�VN:���uw����[�}�QiF�"ٮf�tR�p>v���!	)a][�[��uSp����ӯ?�9'
����@�h���c̍c:�_Z����?��+�7��S ,a��P��.���ў���h�h�[�?n�jU�R�zQ�G:��
�s����]�:�����:UK��=���8�;�еy���ꚺ�t*hE�#�߳f��Ӗt�}9�g2�7����P��'����h��w��yJ���շ��=ؗ���h �0V{<�=M�/_,N���͖�Eq����v'd]�o~��~�O?���CD�X3�3u셷O8{(�
�����Oi�Ձ��@0&�������2��Q=3[���]-�}Df��}�%�/��K^��W1�^��v!5��j`��͍y.EHL��Gr;j&�L��nOWvq���`d�����ݾ؞�A��[p�F#^N�*�IBl��N,3�+�ɥ�����@��cp�]ʾ�����ß���/�\��o�ym�IC�fL�8e�3�d -�G�P+�JnP��tLd?��]��E���_��آ�
�3(��IeT��˦��{h�*�n v,y/�N{3Y���R�����r�T�D�����4�U�7�.^�7d�ջi���я��o��'�̻� IRano§�="ƣ&�j��OI�㲁#��oYC����ώ��׾�ο�����L��� ���P��N�4~,�^AeY�����.��H�ٜ�ZQ_ܴ�9(���&����& �(Y/�O88��,��	���!�a��b�)����U��͑t�7I���)(�4�2Y�5�u��&K��d�?f�aAK�	<w���^��w����WSp��JGT�ʝ��bm8��j�Z֤EEm���~"!��(Z8X�q0_����6������4Q��	9�TS��GӒ��;n"D"y���*�Lv�]�d~ς�79j`���;Ω��<�Y~r����y������,��Uv`��Y`�ͷ�o���{�:�^�.�c�yz��S��N�L]���o�%p��˸�����K�T�)'��S~z�h!"r�b~|�!̡v��B� "���6�(B&�J��r0:�E,˷�q�R�߬k�BP���Z5 
,�>�,��"�=�sq�PbC7E$��kE�l� {�q�N2�봕Z��V���#�� �ŬT�Dg`�Q}���,�r��U��p[��{�L����ʃ=o�˧_�� (�oD�J�Zφ���G?^>b��O��������|���F�r��{���ϟ���!��hT��Pf�#�t�ۨc2�ց������Ε˱+P"�W֎�Y�(#��ۓABZ���t�L����R��  -�<��!}������� �;��9�g��V�d/@�귭=l�������Kfl�~tA�5;�M�z1���3�rz��7o��ݻ����9U����ԫ���h�����dl���Ȟ��;;o	Za�P������������� U��-WQ\��q�1������\�L�*z9���w}�ʸP�� ��@%��� d�W[��B����	tυ����c����QŴ�SP,E@[5p���*6<��g���~R夗����
5[����Od��޽��7o���;)����j�����5�����_�6��X��S5�kB�A~\ro���C�w���A#?�s�n4I�x�R&Tle�����3�o�~dT��k}���@t>�;��;���A����7
ʵ�)����iL���̛U�W�+�%s�6�<���:�y�+���& b~�4v߲��N��6ޓ�����U���J�N�89��$*;l���Ű�K��u�7E���[��I�^�F*��^eEo�����̢�=�ᨆ��:��8��u�JǇ\��p�:gW@K�ӹ	��Y��AE�4�"�R�q^/7�4;�u�D�C��u ��G����hi�sN�k�Q�1������7�ۏ�D�_P�,U�|2�he�%���2:��9���H�P�c$��}V�@W���g_���>$�g4)��"P�*p|:���V��"'* ��&� )���D����t:�u-��{gw6����]2����X��i�GN����h�)�7 ���+{S�/[u��d�z͟�:���ɣͷ�\���t�~pś�H�5Oy�u���wў >;�Idx�&()�9ac]�
��E-{�u��gF��~���DM��yM ����Ơ"y���gg'�	��Z�bD��Y�����͟�
�]�O ����ҳ4��TC���jF�з5�k$q��u�2�DOs��6/1���'Hy�|�d�y���~�Z7�+y�#F��n��������	�F�:��MJ�ؗ�������)$���vV���=�P�F�Lӷ���gN��{�xñ���KJ�b����N�.�ў�>��-��/��F"k0�!%Յ��!%M���LO4�Om��Y�;n"Z�&&�L*�&)�`8ǞY!�Yʎ,�4�+2ɐ�mH�ڣ�H���<m5�ȌKN��,T�z��iq���hI����+!7�k`�vPC�,������c�
�������zO�}��ۧ��~z������@ۏ{��</`�}eo	D@��t���X��]R=�P4��|����G�=c/n\`AY5�J*N�gm��>�ZAPtT4����\�A��b�N��]^\��!B�d�BUت`��ic7�>�����=d����ř]^�r~�{ ���mQd��#<mY�E�>��QC�ƃ�S.K'2z`ˁ>����� �Y.������]��|�_>~��b���:�P��䬵��+�~����U�/mS�
�$�%�ٲ㩜��ԅ6�%��������;rH�Ǣ�����M�GP�J��ehى򴱳~m�T^���G��ܺ� ��������m{r#Zy�e����H���3P�[�+��( t_���-�?��f�8&�H�j��?j��s2�a#��r�y�w:3hf�[<�~�ַ=�)����?3m�I����u.�o�?B����v�����-�eȟU$�o�n�,�M���a��	��b;Q�́֜>h�V]�I��ս�^{��4]^��������O�K�g&��i �9q�Ù����V���pƦ���ʳ!ٝ���������̢e�ˁ��[�/"|Y?�1��t���c���a�NQE�rj��jTX�Á=Ib=(��,�����j��(���~��Xk��0d��x��u�h��dP�<��p)oT c�
Y�n�oYG:`���R�`�: �-���g
�Sv*;����G�1Svz�Z�:�3p6���L�9\�\�oN3���#�r�ѹ�|��g�xv��Y���3�ߙ�����w���߇ɮ���HP��;��@�b�E�@R���>��:�̉��+��E>�����'���k{����z}M����O��_~�Ct��U� Y(�n�[�L�nF;FD�%D��v{��I�uy.&���yoTa����u8���m�D=5O�]�ydr�h����vLs��xt7@��t>�/�s��uf�OP��i�����`׀>�>�9iY3�>\�)�u',H7�Օ1��S��#�U�}��x��{��B&�m7wl��p�ޢS�Gd��;��Gѣ"5T;k�I�# ^�Jg�爂P&���@5.����A�吘"j�'29]#�
s�2�A�P�cny�c0]��M��߬'i%L y���k<>����6{RrG��:����uaN񵺖(�=x�����Ԡ޶+���?۟��G�o޽e��u=?l��1P�=
�_��FuMwwvsS����Pv�4��ʦ��Y��ʌ�zƚI���E�?��{5 ��d����Յ]]�S]����c�<b[�ߵ�	 `��/����}�����z����ia;pO.�qу������I}4��MO�P�w¾y�)G0 <������2��ō�5�&��ʣ��q{ԑH*�-[��b�}9��I�PyY�Y����^o��6J���i�Ĉ�r��f}���je��O��!�U��i�F�j�ٕ���y�f��2s�$�SmtP�,�){�Խ&�z�ki��+��5M���e"����vu�yqR��Xl�g>�����(X9�O��K)��b��L��K�R}O�a�#�s��#��K��$��_Ǟ������kKq*�����9�?z��$�����l�τJp�=��U��kMc�Mj�ǛiDy�iGhr���D9�輜���gɉA�;��1�����륒�R��b&ɺs#����1Wh�?ŠL��}�Q'��K\�R8gyr_z��0��@+���ߎ����왍�;�5}i��f�ZռM�����O��e�F�!"���R�l�?��v/Hq�]5 �@���9GZ�*j��+�%ZU�)���υ�A0�Ni�'�dU-��]P=����N�p<3�f@���hu����������&���3t9W aѴ��OT�	v�3$��� s_:�����>�Y"٫��Ǿ2���}��pF�'����L(�^��g�7���Ϣ���V�.Dv���e~�R����Li3ïQA[esϼ��"-�l>h���ۻ��/@�l��g������� �	J��ޏ�"�f��ŕ�Ҳ����ʶ=5;+(h8��9H�+*�<�0�2�VNXO!���C]��`��[\�ͷR�L����@��m>4���܎2�k��b�ECbf�Y��f��-���!˲��eqJMMW�(�g@���Ƽ1��gzL����xƻ��v��-�	���d})������^z)m�&ӽ�uN�M�1�=5b�aES���)��h	�U������FA�#e�_�)#��Z/����*�}�H4̢j���ڏ��ނu�����)k��~k��bz����nl�,�Ǫ�P�-��kGR���Y�"�]dް/��3���������@A),�^ŖK�g/�=�"keR�Dj���%���
�L� �LwrvN�F�1�2U@4g����+yp�`� ���ر�+{��`� �����<k+���1?:�{����ͯ��O7����l!��՛�����J��)��Wx��7߳5����l2���=�Y_#�t�c?`}KY��H�24�ٷ�a���^�s��JȾf���f����N���͵}��=�V�U'c
��Act���2����k�J&&gG#(�i&�����`�j��{��ڮ$��:.S�I	��N�H�s����)�9�$�����U7c�5�I`�R�
٢J�n��!�� �E����*����޽{g������˞�K���j���'��T@�����<�)`{輌@�����Xs�4�w���տ��z���ܰ����-t=���n����?�8P:>f�0AT!�mU���ZbA˗1t��a=���@���+���!��~DS�o �
X���8��ajP�<ˡT[�,
��D�fb�٠d����U�A5��c�2�(��iӚ�Nw
�魎�Z�&�W��o<��&�ɏ��s�(��[�g<lrn�K<���iG-� #��K��9�Bg���~�Q�A�a�lְ�B�����	z�j��Uw3Q
�#`��Mm��
@��TF�PE�44Pj$O��a�!Z��_�����c٤P��c/��f��C9$7;~Bʆ藠��޺��e�8K㑼�o�~E#kl8�g�x����N�6L�}>g�`G ���c��	@��Z�F�85E�&05��~��.�(�P�?��}}��Ѧ��!����R�kz�t�S��+��uAʲ����1��1ќtL�J�撵�Ka#�����l:W���{{��-i6p"P/�l���#����fJ���^,�H�2�޴�]7AF՟�������a(�{khs�<[̀.7���Vr*��+���;�^790���N���ܬ��^�Q��x��REN|��P�#�� ő�גxM��3�y��MyF�xY��ՙ���Xwbw��F8����i�}�o>�{Ac���/և;�\�L�����>@@ ��}��Ѿ|�X�ϔoG����.��vR�pE�� ��q6u/���:�0jB"�j^�lV��a����U������	�����5�s�J:RF`-O��X;��o�l� s�T@��S�T��ۤ���` $Շn���f��q*�I!���k�(=�'[#,������g�姟��#�#!�����?����Q�(��Ԗ�\v���E�#)���=2xD��1 Yp�˱!���7&����b X� Y ��Z��9����ͧ�uЋv't{���;�pM��x2[hl{[~�&�S�U->�w߽���3��7�0R�a�(�g��bC_���X�;�h�(�[����^5 �8�k� ��(�* �2P;�/�.]�����X&���?ؿ��?�����eôA�o�]2�s[��`tt�����1Z��-�9�7 }&a4� �r�w h�_�ER�r?P�38s��r��]�V��$��u�'�-j��c���l�9ja�4�d��z��Ţ�_��|HJq��w�F�W?�����������/�~���_��>c�?QhNmhrMz�)� �qeD�88�~RMdپ	��x�����+�g��#�0�_�I��O��+�g1�A�7����YA�	�4�ޡw\Y/�
+�F� -��[:��e�j[�?�XP$���qb�yA�7w�cDG�N53L���m�zʇ��;���9P�E��	���(�+�=�U	�L���N�'t`z�>�.{%�(���/Gd7���A1b�ҽ���,��Z1�b�c�c]�j�н�tlD���>_���s����I�|ǔ�G�]��9$�O/��g��v䜫	Y�F;��{'_�Uq���B���[�� U������|"6d�-�KR8�&��H������&�=��t�oNL��2�-��5�Q�$�pu��A؈&��z�����P�Zx��k�+60��Ɏ�����V�'���T�p��zF��gQ��biJM��ńF0 �+�b��$FL��q�76/R�(�K�E�pTwt:PD�"H����z��"�\���H�0���
@6�,f�b�J�ˇs=E�=3+<�dvG�C.1=g?v#ʆ5N��:	�݇A;����|���{��{	;�R�,�LrFGϸ�t]�"KJ��zVH��P�Z����:{k��KJ1o�����)�F6�lTK��y/�c��)b����9x��Q���eY{�`����l�,m4�<��@��U����T����Ӕk]df���j_P@��ي��qw01N+�w���y����G���w�;U8o��r�u ��:R�vtA��u�{:�jv�O�{Q<��9t'�<NyN�2�{;�|[�ʒk�v����=3�����:VIgDYM��PU��_�
�ܸ��<���U�l�~�9��Ծ��_Rq�.�V��#d��1+��ȶ.�C(dn�� (hǘ>���8��vw�kX.N�/ű�����w>�q\�FLL�Υ�;�<0��A-��
��4�<_���WM;���O��ѕ���9*Sܔצg�R�d�aP�5�lz�-AݪY�|k}Q�*j5a7�8���y�P�O�b�˝}�C[�3�=��s)�+ ��=�~ ���@*a���RȂ��:�8�}�Ý�O[K�����r�޶϶�lH�ܗ��8~���3^_
Ё8h�����8�-�V��Q���Ȇ� �P�vT[��4gHG��u��64�ʂ��:�ɳ1涎-s`ò�	�!؂���e�M�Y��f���P��q>=r��z���opj���*��ߍ��z�����^]�U@��[;�s9=Kemc��)8�u?.[�/6�	A^�l`n�{iN�Vvvv���A5g}9���b,�]�����~g�����
���l����V���/v����������%�n�T+�^\�.s�}W1��F���3��N+��	�Ц#kz~��z�q��$s��S>�a�-6nSƯ�8[�s�S�V+�[�D�|>�q��ðs���U��m �^^q�q��g�����w�/ֺx���Qg�����×2g�/���
��Z-Z�y��������~�[�>�h�+;0|wsc�7��<Є{j��(��.Y�!�u��K�F�m 1ȢV)��"�����t#��L��ݝ��7�����L`��Ԫ��X��k=w���J���Yqo��d[���m�O�ٔ9D���<.�I3��G��9��H��BM�kcq�����?JHq ��=Atc�f��){�h.ڥ���3J�[��S������k�~m~���i���9F')�7���T��Xu�c�gD��q'sd�I���U�n�!r�6���7��%�:�R;w$��դ����*QC��F� ���FFd|�:U����|c9�{͈G����ѮMT-0�6r�̵ ��C�0�8׌�@W�"̔%��Tub�M����#}h��e���gW�)�MnmR�D��D|č�U�%6���G)/�T��ī~�����u���Q���?���������G� ��d�'�ڬ�؎@������U����?�霢_G����מ"z�N�'PE�;+��c� �i����ݱ6�FkA4ՐB^2�C�����f�s�'��%mג_�<`��%j���+��!���]Tbt�bhY�I���4���2��J����� N��}H������ߩlT��1���.D�m�G�ׁ@�8�a�AZ�S��~�2����#�$�[a�s	}|߁@�1��Y8KpD �P������|7���r��Ĉ�Kh��S7�lHe��4/� �e[�M߯���l1����4����G�A9y�i-���$jk�q����&M`YAD�n!(���|aC�(�gԜ�E�Æ�W��e�,5��#If� �랷*�F}�j�$V��K�J�k'���v���ʙ�u�I�!YP	H����u�Ae��:8�T��Xk�Rgpe7���<��� Md�;��:�V��
k�3��i�.A ˃tC���=kdD�]tq�&<���$�7[���jh��#��P
Ь�X�/VU A=K�e]��4e�j�>Dك9�TH��y���|�%��k���ƴH�/���5���rq(kw_���Vj�YCy�l��x��_��,"x��2j��5����"�V�Q6g_���	�9z�uw-i�tv�AF�8��a#�@3��*�h�������s���y0o�}||��甠����K�V�����{W-f;�욖����m�3X�`j��<@!�
6c�^��b!�S %T*Ѥ{�j��J�Jh�<@�=�Y�S�m5�$��e��P�&���Y� xzjCϘӃ�(�٩17��9) �����w?ػ����=�w�^����MPŭ����5�pr5�ٝ�I�8��yXs?:0G��w��ER"XG5�U0#P�D�ԛ�����g�S����,x�Z���I���#��d}ؤ;�Ŧ=������ �Y)W�V��p2�̀�! @��s�(�j]&�	�N���6B"J㙬�5�!.k�d�Lyv�/ 7�٥�)0�ձ�$��_4ל��TU���{�1��91m��:�ܐ*`�&�����|�J���r-�g�{����[�?�{�P��X�"�����#�x�@�kܨ-���jX��F�2�;Eɂ�Z#����֢�qV�Á!ML򦅘�ThCDv�){�BV��r����qe]y�+�k���uDi|vIY���ѻP�So�aE~��^W��c�]%��)\2�����l6�u���0�:ũ�0�@DE#s~��k'2�Ӝ�y>���Jߞ�/��o=�)[sZW��0��
�<�G��J%���i?ѯit�������P͢��YRTX�
:se3���S�uP�6�u��Y�%��쇑�ӛt�g޶�co��jw�PmW���L�С����L�U1d�[�x�Gk�M�<>�`t�:��[�4��$y�Z7�`�k�q:R�U-��Ha�ܜvr��Zem�V>A��hѧ���e#�<ޱ>e��h��A�|^�ӭO���`��#vs�=���sk�*�fP��~c����i�O{E=��s��<V&�
��8�I��f������~���7�tkw�?�uC�=�W웖4.�����
j|z��"b�����6����W��Z�� �v{� ��=�<Ξ���}����'��$�r�XW�Fs]��CD��f���4����<�@�n[��2�@�CO�A�k�^nZ+̈�$�r6Eu�ߞt���Zxq͠��r���j� 2hE*��$6�ခn���5SgM,������;D�e�Pہ=Υ�c2S���4f-�3)F�E��hX�>K��Ŵ��ř$�Q� u�lhҬAY5��=��2���h*��C�ab� #�f��q���N![I�q7Љ�ga�A��.�����2����G{�j%�pݺ ������y�FvK�t����w�`A�R
$��� #iӸ^$�����"������
T�ڧ\�BF���0���9�i�=�
 *�C��Y" T;aP[�s0בA�.K���t@Ei�p�2��]PQs��M����R��:!3�;r�������]��`o>�`��y*@k|z,s�yf覒mFQ��fa�f^����7O�	CW�e���8����3�~
qV{y���ޚèV��Vx8�DK(���^��Rd -���=���u�����ig��'�k�&'��m[��i���k�U�$R}ɯ�qcƈ�rI'i���SS�Pj��M+icD[�iw��1����ɜ��ɽ�9��.�M1�q���&L���I�o��ș}��@W���Mr�"+�4��"��@�NG���=0�pl� �v,�ǭ~�
��
��O�'�vC�D��f����`N��t^����JQj�t5;��F��n[� R��?p��-}nOh���N�Q��M�BM!��F�I;6vl!�!�5'a
/����9at��&}��6���(5<�׍^�=O�hn�|NcK�H{C\�u\��|��9��1�룉�F�1����S3�y�d�kl��8��y�ά�4)�Mʳ9��}�E�����e�J�Ԏ1 )֍߷�]������><�°3�2f���8)���rF_7mmg�`<pL�$ٳ��� Ǳ�)�u]��ձpeT|I�m ҍS�g����48dO�
䝓D0��q��6(@�=p|ػA
]T(Ħ�N��Y:��WH���7��~+�ÒE����J�#�c��~b!*R�v��cC�:��D�<���������6ٚ� ��z4�ڐ:Cbc(�����d���Q���i7�'
c��jh���H�i}3�ۏ�k��j���ʘg��dڻ���Ё�t�9sz`x&{�@2X��@ﹱ���b=`���\��.��..�'�j����'	A��oT�M��%�!��RH�#;��|�u��d��*�d��lź0)�QԢW��4#�-���)�����*�6�x�j�� N-�:��n�̣���>t���3g2h�'�b�5�o��{�$x�����i����	)m �b�e�E!� Uܦ���b�2(l�`L�!k�c��,c��a`�t��Q=���"�@�I�s�g�vS���L��1�}���Sv<Ӷ�<�� ����իW��(��#�v#�0���.L-�<[���m�w���@���R���e�Oh��ӔY5}���S�<��v;��'�c<�^���Z����cdl�A2��H�E����ͽAUf)F+߄�	��|�k�_R�L���$[�0s��/�1�!B挊䙩&��u�����d{�}����Vo��2�Fm�.�d+�l���n�A�D ���gH��J\.��v^��UZ�7l}�@5l�6��M�wr쇪9�UR�s�4��>E���������9���p0VW
`������<��Ef�c� j�Sd�Q��<-7d����E`�V�u,���`-�|�M���G����ؔ��|���E�*όRuL�nT���tCc�iBµ�:GӁu0lJ�3��>W���gە�?�+FͲ�F}�V���֣y�0��C��7��V-�,�y����y4�K<�y�?C=�H����EV+�S�$BZ �*;={d���}{*�F���֡lƻ�9�D)Pס&�]�&��Ftk_r���DQ)�,�s��MŸ�Vʑ,��)�-��旌�Y� �U$C����^s�)	8N"}���	�%�k� Y��=y����8t�hi�Ȫ�x�"�H΁��l~q�c�����^_k���q@�.�fIY�)33�`N�-D7�h���ϝ��s��2��f���k��q����8���q��,O7����rC�.y4=�^�y�p�a�̊$�ϣ;c0��v�c�>�W_�`�/��l�w��lEFG�۱�ɝ7^ܟ����.6�V�Mv����U
�
�s��{��û�3d�V����|�b����>[��^��6K���{���}Z��q[��6�<�JJ�JL�M3�G���uWƺ+T,48h���~��:�Y��%���K"�;��A6ܔg�����!��_[9����u��x8A g���/�T���"9�2us�YpTS5�S/�G(�G�zE���7e����~�������W'ꕋl|/*v�ysg�����������S�7�a��G�����v~qeWo?���+e�@-ŎhÉoM=͖:�r.m�v�N�8N������V����[���,1�q�:�ǆc޹�%���y]�� �p�H�N�7��s�
p�s'�=��&i;弞˞���`���}�0�j��虫S�[�)�F*�fǱf�5&A��S������ Ⱥ�����+6&U�Gb3A5��s�kE*ނY,�f���E�sG�!��sos��B':
��62��V1�L��4F@����W���}���0��-X�qqqɦ�������H�QB@��%�hg�Q�~�\��
��~<1I�7tL1fk*
 �:���z��-�O�>��h��t�${��0mt��a]�%�v�*�[� ��b0z'��6�U>1�X+�uӲ�׍�������`5A�����:���;��z9��㸰l|�~��IP�l�5��u�9ܒ���S��2�Xwɢ�������脬깝]����7��<���\	\6���QcӞ�kjR�N-�����8���FP*���o
�LB{�J�5ߥ
h��㾒�xG�+c��/QQ-FFqfcY�je5�5
Ta_c=��C�^�p�=Q#��N ���2�t����զ��ɋ����z�o9u*�� JHa8棚����:�#B���f�~��DU�@��;��ݳ&K�8ƹԄ[
�׌���5�ӂ\j�y롵���b��I��4�w�����fܱ[E�s���f8��}1)���g$9g_����	X���� ���I �׳�7\��p��<������5%Qѫ� ��������j�ȅ:N�q�@Nw��h�����&���Sa)�B�^N~��$�$j�P�`9�F&����� � @V�Bz �r/��&I{��M)"�j�Q���ik�Σj�Y�o�7O��@y
�n���*��y�e�䴙�+�1�'���W�b�`�dT,��W���J/ڨgmG�\�@�{p�ѯy��T��3�5�����
6[(+�Y"6M�Dy�ܴx�4�`���>h�"��^/�(�"|A���,��H)�;�%P�R���HՃʆ�� Ri�Ж��	��A�hD�A�>�A��7��
�#˹Cm�+ o'P�D:+xOW�c���s�!�Q⸃���oÿ�݊J(����TC�r�I��m�� �A�������5c\��8Th��=pJY@z�@'u8d��J ��J�{Ee_�}~��ϙT4	 0Ԍ[[]�P�㲜��T���g �=$�f�5��,ZG�'�&��xT
�>?��_/���U��6˲U1� �aO���k0�p��` �{�>c�n~�ϟ?����b��~�D�Cuz��s�z��._�-�w�Q����k[���&�PfEs-{�kL����xǹ1 ��A�)̂������T�<�%���]_��l�a�F i���Z<F�Qˀw�B��nʶ"��:_\YNYfe����M�!�X��۲��=���y�R'zcE�+彜"ƀ.2H
"rfX��9���I��k`�z݁׀ϣ���r�!��57�	Y�F�B�[���;�ô�8[��⣤ؑ��Z�(ID%��r�ܤip��ڶ��fW��v_���U�@=��1�IJ}�s���B�,砤�3U7�'���戞��҆ʋ��>�x�1�� d�A��`�ꠞW�a���э�N�iX��=�Ⱦ<{��ۭ�Pb�<AU@n��B��dQ���ш2��u���LZ�t@��te�>Ė:~P^nİ�=]�E�U��g�jH݁�f	И�|���a��\.$jB�6H�� ?�fk>@o��jN�C։c�^b��w���ֲ�{�yH�vs��� E��A��lc���j���f����������i�u���+��~k�O���T���pM�6��G�H�^^���71�&󩲐4������T��y�C���QI����ɧ	p���&�E8�q�-v1�r�}��ZB�U��'��u�g��B�d��&T�ڊ9�͂_��}���_q��V��3;������E��8Tqv�� }�w����v��^O�h�^Gt�1�	p�Vؠ�hD7@�c㲠*NN�
�S�^=Br��b��������3:[s9�I�vڊ����9�ܔs�$'cD�S�
�t���R��X�i����n�A����~ ��-#"űB������޽}��t'hA9�ey���N -���ZQ'J �{�L���D��=��kM4�Ӽ����|1����Hg���j�15�sG(?�}f6*tc��EO~3��Pו�Y�|��<�c��i|��1&��|.qÚh6u�_9yd�Tl�~}����B��.�Ms6y ��;B�T-��8��/�W���0�CU���^_5T�8���@�w�^Ӌ �%�4M���m��l�\s!�~��_�[I���*�Gʵ��@�A瓏�*�c�x�A�$��O���mZׯ��& TZF�W�_�f�M�LꎞEԋK�$3��y�>^��Műؘx���ݏ�x�>r��� ����|j���"(Qٕ0�ȷ�	t����� ���+�c�\��g�>/�97��I٨�����Yo�=ڏ�P� f���2�OOO*���b����S��Tp�]�����*���z(��8ǧ�ה��P���W��F��S�i��>��2����8���6���4� Z1W#R��$�� ����ԓ�oQ�P�9 �헏v��_���l�>}���O��S�c �8����w?�ή�|g�\��Y�0�%P���, ���>�0-���� ita�,��)���∴�R���� -�@B~��`��v�3A�zѲ����,���C�� ��u���3�����Û�k���gvC����>?<ۗ���Q'Ѳk߫0zp�I�j������f�XH�3@�
�&� �s4����{ 2���1`{��Pқ��L)��5n߼�M��h��'�������@Q��}KW]��X�׽^LL��8-�QC\զ��(Z�α%P�
�Q�̒&���j�H�M@P{�h΁v鴀	�����I����
�^Ӿ��������/�J���7
%:�Fg���i٫Q��8��b(�@~??��� �� `��|���~����}�"5�d4C^���� �S;�@��9�0G0"�xI�C��۱\�U�Mf�uY;�0�;P=O�-���2�S�"|���=Q�����D.�����ژs��҃�]^��C�A(��:՚],BQ4������Z�f ����]�y�@ ��d�<��������|�����~k�߼*s����� u��\���5�3�H Y=7ց>��}kΨ���)#��Q4�y��W�_%?V~���60�6�`�-N
bc����K�B�<X��/�X�U�QoVR�P��x������貵�T�D'mw�#8Y�7��.�fQ��k�6�9`ŮxN��.7��J�;wC��md�Qt���~D٦�zU@��0����nO�|����Bd�R=�T�%���~i2����qIc=㳞Ur�/zfE!�6�\��ɿ'���s;����g�h݀m�eY�K�Dxr4Sv����V�k�z+�H���������Ö�	�0�������޽����}�恐]H��` �V����
tY�
��r ����.�u���� ePM��T����N��B�	��s�q8��Y��X�ߊ2p�Gv[g�J\�h�xA���;�6O�W',M5@�?���	��PL�����h�i%a���L�*�D��W�q��LTw��M��et��h���7̱�_�j��}�<�g�lcvL���G�B�QF.۔�"�Я�k��ee�Ɛ7��8�+伓�Cn�u��\��}���>�l�޿��Wt��?C?��4a�u����A�h�iU��W����Z�r��g4R�e��z-� ٣����V��VJ%�Yl(�<%���{�풦8I�?�w���ƌ��U�� V���O.��^���5�y@5kN�MXvt<�Tv�^�B6"�+v����}���N��\���-)uW��$�`�-;�����������U9�WšQD�y#�b�W��2��j!Md��<��j9���T�D }u�5;�W���1���n��nY��� �Z��B�{�P�˧����?��_��g��� �EGj������</��[��0�c)��o'Z�|#�j�h�~���*��F��0�z@�\��
[����C��Mq��e~�t��nQ�WST�ե��C�){�A�l�K�':�*H�R�� �ǲf�6d�9��64��9�O:?��	����WUA�"��UyB�7�k�.//�\��x}�����OT���<c}�g(]���N|�7H�g�J�O�+�Nዖ�C�g�{=�@U+uD�[#�yT�hjn��0{����I�K<�硵�?� ��E��V���1˿XЀ�5xP������͵u�d�ݢ��M��������z6	��e�G�m��c0�2���@d#ň2��A��x�w���;������?�)���v
���l�P1|_��?��oi8�<����h`ݹ����FX���pF1�,3�%T�쁺,ju����h��sE�j��l0���p h���2s�@�-  �æ��깖����n�%kuq��1>\�ggTD��PĚ���:�?��H䔾�Ð�S@�o��`߽M��Y��=6�1�(jP�E��8�y�(c���Н��l)�2 Y^Zb����������Z�'��~�}�f���t��ņ��ti����/H�;��	�C��q�K�}j�Nm%�p��]W�+þ�ܣtJ ��Z�U�hJ9�t%w�����i��e�X�����(�ّ
(���#N��B���bJ��l��*R�R�u`�~�{*2�=z6� �SiFI O`�d�(6Q�Q�l��dl�3�6�p����,��:9���/��\u��N�	$�Lc��^W�^�vw�����m��qG~�y�%���E�8޽�`?��G���wvyuQbH�f[��z�[q�Y2B�S�jM��ʵ)�s`4��4��:���z-�g,
o1���}�/g�����+ӥz�������u�9��-���ëk� ?܇կ�zw��31�{I)毃+OeO�����c}T�a 1�J��� ps�'�;��������2�>�-��M�%��5^�7Q�׏Ƞ��;���1Q�U�Zŕ���
�浠��P��F��g�Z3���Suo�4?��B{�� �>�b_��Ɵ�N��������󲑯x\F�R㍍5��\�i�Z�Le�&���ʳ�"I�6n?��zϨ6z���ѷ����z_�2[�v�� Z)�q�#S��B4����J^{��v`�9�փ�P���,���溼~Q6�S�'����,�%a,(����4����T���Xo?��rO������a �=5��6�������
�a�:ҫW;9�m]Ωa�8ز�'�R̷,�9exD��Q)X1�g����i}������ȣM�].=��]<D8sW����)�����/&M�W�-�S���^]]�������[{��W��-v�x��Xp*)����@�2�q�ju�ù�B^ڋCl��*i��B���\��,�y��\�RN�'l8�E����x��xɃˏK]��G�a8�O��}��/��}׫�J�2 �3�EF��Պ�wL�
����N�-�= �������kʐc�D)Cq� F���q�55zm��*fBp�;ͥ�='3�q h ���n��G���`M���p!q �!H3Wn��f���N���V3ֽ4��]�D��]B�34HoT���b�Q�s��Z�-��D����1U ���iS��D� �b&e��H�u����h)���5�/e�Z�Ι���l[Cߠ�q9�O�>��o�b?~wn�ם�~u�O�������>��8]�51�$	���r���Ov��^5�!ZQ�U>�ޝ������u��h�p/r�9P@��ၾ�Qˑ�<�t�R���J��fc77��� $�+������ڕ��aߵ�i4�@1���A34Z�t�Ѿ|���Í�F��p�U��yzv�� �w8>��U�������:�J�,d��w�-Ѷ��d�Wʸ;�w����w�{��)��&^R
��]s����3L���?yf.��f� u�/&B�JF(&�"��`"��=�YS�� e��F�:�b��ռ�!S�+Տ٩�����X�#Em"Ǳ�z}S��/��ɪ��ށ�QϾFJo�s5R���xAk��o�/ޟzE���h�\D���W��� YS;�A[ج t�2�.�`yJ1�]��{�we�K�8���^�P��lÞ\�(ҎOϼ�#�8T�R�V\nc���_m�{ ���d���1��J�~�lXb����9�����c�	Dl$��[S���)/���h�ݞ�l��ҙ����c�#
F�kW���'�f�2\�QLuE�����Ȣ/K�ҏ�T�q�l�
,W��g�#�*!@��c1r]9n�W}/4��\�c.���%!E�kf��B��y��XDv̹_u~T#�s�"��s0�{Y�3b��@~�ߘwp�8�:���5?�:q�f_|I��B\��1���¬8N���̓V3��������B���N%��'�>�@��@hZ9�h@i٩=�=�����|"ا��jZ���ʴ2����
�7�^�E�U�܋��#�]�C��ܩ[<#�I=�@CD��MC�bY����-�� 赭S����3�'�@�e��5�5�r^@���^�/��^��,6$6^V<͢�u��8���7�)�����>�������v������m�Ɔ�N]�<Q�XۡikY��r�m��y����2.�(̂2�]@�:��9fW�l�@>�+8��Ӽ�#Ğ8�0��l5�hM��4������&��KE덁��G���/�ϟ-��a�E`/�2G�.������������o���3C�80�O�XEդDPJ���K�=
(�1߅F�f٢X�H,�iM�Hgx��P1\�gC��]Yg��(�P����ҹ����(�>�j�D�Qg*,Wp"�6�������̘W��]��ƃ����.@	���A���b=��b�N�`��g�tޱ?*��L`u_液9O���Y^h� �ދ���zz;���O�'e�.�ӻb��p�5Q�R��xM�곌F6��<��o��M@r�/0�$�w����X���@I罥E����c��ȟ��H��E?0�ϛr���X K
9x]&�A=4;N9�����
4���j�k�^:�Q����K6e�%�`%���Ӣ��å���ޗ����	p0���[ҽ����< ����y��������K{|��b���NX����Q�uqqƞU��$� AY�,>�����a��N9�g��y�N!�$��Ͽ�jw?[�y.6���o_����] U�k	4��
�O���tsc��zew_�p����](���P���e��o�Ӯ���I������Eʾv�<(���U����6�x_��`e�4���v7(�V�-ΝL�܃�~X�g[��'�=��ό=_����E�f�@d���Hu��Ŷ�Q��t�֕�����*J�}�\�M�6��J�կ��D����旣��{G�R�b]J�0H�vj0��4�)��;���V�,�'�aL¶�;����l(e�BE�T��:*��Z���D?��F�WlbqnlU*u,�E�S)��}
z�~�����.^H�><�Gj�|����	G*��a���N3MNE|ew�*��u1���R���yB切��@4����Q���[F�X��+sE�o�N���so1�8?�W�W������(]]	d��C�FQ4��	G��B�����-N��/O�,cW,j� ı % ���=ت���^#�褚�9�^\l(<%��S~�M)-�l3�HX�E���?=������ئ���yB��ͧTR-V��1����4K�����i_�C�Σ�f�k��Qw��j3�Qg�u驆�� �^�>�:�{eW\̢ύ.����s�Jg�8e�"|Yh3�R�����2u�����s2jNXX�cr]��Q�^�;�"�⶙G4��H���4�c��=7�޶Ł@=��$�0A�h�aⵎ��R��=SRz��336��F��DDv���\�m�v��=��w_�kS�/�{ ,j&LΝ;2��,3���{�����[W�35��$qX�_�cS �b-J^Cb�d��l��u#��d���Zr��Gv͒�R��b�C�+�ɾ�+����|��G{�݇�`������O�'����@� ����yk.A3��J���O ��%h�?��������O����?������2���d�:O���l���:������2�=
���񸵫�{{x�hW��۫�<+T��"�7i���h�Np.1{]�y�j���ڄ�$&�
��\ �jD���U#is0�]DG��:&/L�*��a�lEq�Qw�o��z���n��Z�hyB���Gf�0��h��5�A���؛✽��{{��o� �T�\��,�YÎ���I|�L��3-����(��>�i��O,�zoQCI��Z�'��8�����W��B��P������^a=QZ�?��aD�������:���l��ҡ�	2-fiVe>���}�˓=ށS�)��KE�Q�cN4����^�%�a��Q+E*�V3��t��g|ѠF��h�}lX
!�{�xS@��?�����=���eqh;�PPI �,��)H3R=O��#�A�?��O�	�1��F������a0��@L�n�_K����)��y�-x� ;�e�N��jU��zY�����qC��=�����V�Z??/ pM0����Z*q���;q�����2�V�����y_��Ayl��q06Q������WG1�ZC���o8�:���١�%jiad�f(� �[���ʡNO��9U>k�4��?A���we���~�F��ȗ��;+�>P|�G����ig'
 ��v�����Xw�=G���ρ��-f����(�sU���� d�.ΐ�:���o6;;<����`O;�n��+���ʼ���a/��Ǿ �{��lB����Y��H�U�
n���ޞ�>�ݧ_l�xW�=0�Z����D����N+���[��Ƚ���=80�3������hj�k򉧐O�l9��׬�03_�*�"9��7i�ؤS��q�h�;�ڄb�U�J]\��!��WD���eo��8l�L���[77���QCa�*.x�� {���M�
1:lJ=��KFr倀E/9���z�XSެ��C���5����L��5|���;�-Fʉ$����+��Q�@'��eC�"�i�=y�g�{7�o������XE48'����	-i~A�L	|�;(��=�� U�=<T��0�DhW�:^j�*� l��j]^�wN�YC=GW�����d���5s+��ޥ�j�
ifz�О>kx��A�'�3�j���ʡ�s��~�z�,(�Ko��
	D@�	>������wRB֯��@gcl�*���AߠhJK�w���U��4_�s��e�%����v@Vz�,�=���j�j�e���d4╀�_G{�����e�I�s1����G�X���~�M�S�Lfp����w+OT�z��=��UH�{��ެ�X�Ú��mI$}��H9J'��z�s�/$WSc^޾}c�^�b��y(N"�777�78�n"�n�D�L�I���I���<�Κ�a =2��{nl��[�ع("��(��(&�]��j7��j�`c[B~��q{/���2#��߾����o~g�߿�����Uq*^���Л�j �Fm�"��T
�	��i�E�{��sU�>��ǿ��>�},�uP�?�{���<�0�h�,Ξu�3Дn)����{ʖ���ll�b��7K���Y$ԃd����lee��6.��RЊ���b���i��bm�%P�;�.F8QP�+����8�v_���/�xc�_(vad�NVj�1ܿ�D�*s�����������p~$�ݚ��������U,�4��i�N�����7�tS�oI��4��uR��8���[f()YM���N)'=A�;�৵�8�,���E)ۗ���i_���6O��wk�� 
�g�I��`01����JL��5N��{&��l8�F�E͚��u���c���� �x�:c� �[��7��!p	��")c���j�H~���~��(#_�в�̲��'m�y�d����Uq-a+/.ι��S��za��S�L�I�K�k�.$�����>/��~� ��W���F���~�L������_\�~�^M.�/3�9��ᕻ(a?�F?#�������%�R;�]�bUl�+���T�[������9ؙ�7>���T!��>�����Ś�}
#��u�g�L�^�| ����V����r�X#�hN���\��7d������(�#M����.!��`+[�+���\��~n����i٬p���.�,�{y�o5M�1/@;��[�:��C�<T����ϬK����iޠS3CKs���T�1~�9�ݎ������|x2k�xL���k���_�bǥ�uw\и F�zR0��g��� �m�-��H��ev/�
�E��2��3{-�+$�>Y~�fTAV��D
Gh��\h��&@�xeGrU�]bl��V�����A:�`�)��ߢe�����[�lI��X�S�4��d|ȶ��H�o��q��h�	g�|m����c'9��i���h�Ľi�$Ǒ%���q�Y�u@�İ�w��~���v�EvH6I(ԑw�������{d��H�L@���nn��O����W�^%ٺ<;��ޞ;(	�+��f��ߣ�h�����c��P���h�����>`��!1�>74p��v��כ����lK)�Ħ�&����C��%j5��{ �mp����Z���f#Uf)���s�X&�Uj=w,��lﱹ�9Ȳ�IMG��$��pyQ;|_d�K:���Of�@�+?˞��C�m���4Á(��x��������>ᑃJ��7��r�P��ߘ����2v�k^$�{����������op�[���$R<�[S)��Fo�x�m�V��-�<����D�@���_����e�i"P�}uuE1�GDmN�ZR�ȹ}.�D�Y
�܇�������3���,]+H�"J���(�a�0����D���<��m��ٳ�\��ќٟ���V������͗r��<ͤF��#c
$�K��\�31�M�PUź���w���Tv��(:?W��v���\����^6
�������n��>d: ������pj� (K�ۣ��39?{�6�T�'Wuj��\&�����[�yL�:I�5P5#��c� G����P|c])����}w%�7���������u.9o)RԵ��XeЎPH�v'P�:՟��>�z��^�K�cO)ALƆ�\Db鰦�7c�ux�����#00���uWh��
 �J�U� IWC`M�_���ų{�lM|I�l�:�����wv�W'���4܋������%�g:�h!��e�F��)�p]��¶�~�s"���6�w#������:�mP��{���u�C����"mk>�ˋg����re��Q�03C+ d �/�r~<��/�y�~��f��3sJ%�#�V��/��)����ǵ)1{]�V��v��~�P͛(�H�@��~�E������q��uMo�nJ�O9|:�Nd���z�%��o�������\^�|�v�B���lm��"��g�b��|ov��u:��6lP5��M8�sI����o��7��J^������~2E:X��{��&�ڔ�Y��ó/�}��VkIZ�/�]��Js��=.*���%y ~�ś�(j#�� Ȕ�[�s��[Pl��km��=m̃謬�o� �e�*���D�c�&k���(P��k�:.nUg�X������qpMP�ŉ��)�:,&c�3�+N�wڳ�6CY;��QP&l�(�,�OO���ul;Gj�w�F��������Kf��w1���~�끵�F������_���l!q�k�ـ�1�(�s��	q0���`0�V�uW�8��f+����!�D���oE���z��vvq��fr-� DOG�����p���:r�{���XT ]j�Dd��F�q��)-�ߗ����	�Tj��>bcn���r��Zۜ��EX;5�-D.��
��|d�a�3w��#N�k2�.�"� ��^����;�;"y�=@�e�\�4�1Ŏɢ~}.���Ŝ�uȌBw6��a�'P,<"�u�K��>�-�����
�����MWQ�E@����J��̒��� D&��;g%J�<�^g��)�-݄9��!����6ЍF$D�эF��	��JF��n��Q�B��d�K�����	�sz\*�D�m�2�g2��G��T�>>�C��̣��J~��oOĂ2���R��S"�.(i�hO��@�+�%a�y��z,ϲ2|C�f�|=�P���	3���  `�	G	N����m���r�� lCZó�����I����NP	�TE��m�uBCp8�;9]L�w�7v��1�=+�"{@1�BC�2 i*�������o��o��^~��wrq��TI��0Ue�5վ�0 RPk)�[>�2A�$����rr�6G�9�����T�
:�ݒ����z�C`���p��l�ٮ�WB?�>O�Υ]�>8��
4��3e�N�UEFG�Cm���C�fX6vQ&0��0��e�����Cv��Ou��� �n��)��Y�LA����[i4�(MԹ>?;��Z�Xmu�lu\ ��B����~�[}�|Mu�����;��uŃ������x�D��X���"��ސ�k�D��sOz^} @�j^�J����-�OL.[�bj�e���pJ'%��dS��*ad����r����^�&����\��@�*����ĩ��))W��VoY[�C-,)�Y��  J����wo�y�� 6ߞAB��߹٬���������Ec��*��:�u�O4�-��\�>�[nQR����������,@���z����g���k�
���w�.[1+G:���@b^u��
Bp�7d�qM���db{�du�K�RdK&�F�kc��X��}��<�|.��[���, �ǻ."h<@ׄ�Ӱ�Tcu���@��Ĝ�zm���x!o����W���3f����ϫ~��rͺ��~���B��3f[�)��îA�{�i���	��-0^A,6
0v��u������[Ǧ��;�������g��x���A���S�������3LN�D߶�����-�&�[�1�8�lWM�󠓯���x���9��39>��o�%y O�%��v���?��8�[2¼ij�r�ݧ�%�E\�.���K�^����'�%>���������N��(n�Ge�w�}s�e ����2M�T����L��fJ�f=���czk�x2���	��8�'V�qP��bL�Z_kˡx��J����8:O=�o1c*�
R;+�t�d0�7�@�E%��(2�����%x¯8^�h�1_2�g"����ѵ�F k�����[��!��!�	M�n��K�﷚ ,�f@-�C�}wO�շl��~2��g�^��T��4uPجw[Ro��	�o�+�E��(!-��Ų�|we�D��Fq���1ӯǝ9u��JACz�Sn�����;y��J����ͣLԀLhM[DtC^w4|x���
k*@��ln�e�D6-s��BX�1��MF�c�z��ߔ��E��xP��`nts����IΑ+H�g���6�c���ǟ���ÿ��?�P��H���E�o�Io	�0KR/�5GG��}��+��hF����RD;8�9JX���\�Cct��%��SAf�jW�T���:���h$)�z|4G��I�j 4�g
�.//�t�ՑU�=���Ϻ���,�5g��G����a���n�}���k[���`��e�^�qiQ�A�����+Nw��W�/��سVK�Z��^�x.�|�������o����/e�%^���7�VUn�$ҘW��ͥT�dx"��u��� ��:�$5��p�Y-ϳ�;�rM�V��������nyAV�� F��C���{��P�U[s�/�k��>c18T� �'�2i����2�`X�����e��N�� �r���c��
�vP|]8��w�G�>u�oo�����bo����l�\m�B�k(����R�����>n�2�1�|�J��7rt��}?5�R7�hyM�5du+@(���"�{ԯybo��.{�׊�	�n�_����:9=!�g�e��%Z�x���c��A�K`��Vg	���e>*ʳ���|X�����f���i �5B�}��d 歷���S�T*xټ��E5ͳ4����Ц�e�̣�>y3���)&-��T��G&.�}���w �#�k�.O�\DB@����i�,(� �oV�N!Eۓe�QW=E��V���D�	��Z���!��{���9vk6oZ݉Lէ:=�T�����TC�����K����3Y"Fk���Ϭ�Vb��O+
]���Y-Q[�ӎ�m��Kvkw�AD��;3`	a�P"�J��&'�����˗rrvdu�؟�����?BeCۂڬԖy�iO�cN���F>��3�A'G��� ��W
ht�f��ڷ6�S������`bO��8;���S�0&N]��l4��{Xʏo����5�/Ξ�Ź�Ι/&��o��7׷�A���w
�W��� O�B�xi�Ĺ��+�c���o����&Ȃ�������K�m��P\�A!��Ȯ1K�,�g�XK�xO�*��`]�J �SU�r�����{�Oa�(��|���aG���#Wn��u��0���;�E�O0�6���(:��6̈́ XhS�:q���~��&���鶡����%�T�7�������bJ���d'o>~���C_%D{n�-�̔PUT�Svz���ڕQ� ���f�ɕ�
G3��3ySJ���+s�_�@bB��!�%�s��_z�����q��6�mWF�h*f�:S,�L���W�����u_^���H;���UH���,QF߂�m��e����G�	�f�>9�+��є�<C�uN��8�m��M�X���la��0�'�3A/��R(����c���S��R�ޮ���gDR]��>�g�f�Q`Y���X�;{�MZ+�~G�)��{�whY��3��ʳ榢_�Ȃ��d�ź�{���d�ۢ�2���Z�|B�6����<����=�.�>�an���@(��Ħ����1���^~aM��r��d�?����[�{A9���g��<4�E�	�]�-*?c�wd���o��c��Ȧg���pcdOm��bN�}W^�~M��ۛk�kv��{�q}�
�>Wb����uh���������J��l�И�f�i؟�����:@��5��L�����/���W��V��qGcL< BEP�g��IF�rjX��rq��_Ϟ=�"*�T��Y7q���o� ��c9y�3������Ln���n��c���&�#�[�O���F�K�Tߩ=9e؜��K��S�����3�iy��[�H�H�A�K��/eΚc�,(��I:蘹����j����^�*#>@~5W�w�R���z��6�P̎�/���F�����f[��#���J��^ʩt�?f�+��9����>��_L�R�ڬ�b��aPuV�{�=u�T��]�F,UOzfϟ����� &0G�*U!�k��mmW��J��NL��^�d�6p��bYA&h��o�r�8,��b~LP�l�v۳�T2����7Y��٭�ɳ@\8X��Jt�9==�O
]��"(������u���_Ij��޿�A~�A�����o�_��;yyy��A���G��F[�������Z���E�^���_dU@���<���\��Su���+0��	XNtN�����W����N�ߑ��@��?2���i�>a-�1(�"sw����
� �ι��؜�X,�#j��a��/��b1]�x�5Tj��:]ۉ=�`r@�n�o�X�1�bkS��z/tN]��lv�z)V��u�c���^ǚ���՜�r�[��nuN�򷿾�?��o���[����痗���O�X�6r��3-��`�?��?��w���"77w�G/T~���E &���vG&>��V?�g���;��ϟ��߼��|��R���N}�{˝���?��统>���=m ����K��>_+���][�g�_�䃞��?����O����uVx��ߞ���h΀|6Pf�D�fb����~8��}02�� F���
2����[(C���� 	?��@�����I|���-�����0cu���ܡ����bV���~#�O��щ1 J���t�,o�F?d�g`��b�s�FS��҆����v-ّ1ͮD��sMm����4��כ�7�=��B�6���2�Ԗ�)�����X���L9�ޓ�*�~ON7?�Y� U=X�Z�Q��D����� m�ˏ��$�����&!)��\�Ū�ݪ�!ci�GC��uM@Z ���{��b(�0��-JC��<,}�(��Fs�s@��4tnGS��3H}%��O,*)�>4<�5�ݕ��g#1D��t��9
�hz��	��
f�NhtG�]�h�z'u��M���$�����J	��8NI{���c���)�f8]d:YCK�D��&n�[k�I�3�so�-N����Ұhr���T��5d���q�) (���0�|�:J�X�4�#����==ίM�Tw�R����K��2u�F���t��o$0a���aV5bsJE��l)�+�����x3��6�Z&�H�{\Z���8�e7��4t�/..�����X����x�	 q���=2%њ�w�&����h�ڵ�d����!e�=�&3�	���(vъ"��m����b\8�_�_�V^�<�x%�:<�P�\�XMHp(fB�9��a�G3�W�5�����h��Xo����U�@�0e���:&[Y�@�Yy#���ĳ�Ƌ�,6��Ol�z/�խ�ݼ��"�|��d��,2�P��>�v�h4���e��k�6f-kIlc��=iC���B)m͆���iZ�y( ���2�������:�����|A/'�^>�s
;���T�X?�/McBF�	 z����=�S�Ch'J�A����Ϛ�d �쓅%�
xe�	l��7W���:��u<��y�n��h�s�$��6ۈxo�mY�p����n+W�{Y�l�0{�r�X�9�>bvDXGdN%�/���q۽�7X��r[a�i7 ��Ս�n����2���-w|��*�l �ۛ+6굜\��W��R��_����ۗg���	�ط�~#��/୺��@ �`�Qo����f��5*��AYxkl��ԛ͔~���gg:7�(�kzvzB�9�d����K��~�ѳK���GJ����� ��m�^�ޛ,�HD��xf�)�u<��[j~��z����^�����`)�������:�e"P�������f�=Cۉ*��
�o!]���k�ᇟ������5]���)zVQ�#3��5�L���[��w���;��ߟ߬ՆϤ��t���^.�>[�6 �����/|?�a�_�`v��v����B?�R��rus������!���~���ڨ���������Y���~����[2�fj��_}�w?�_����/����>��r�`�����~�G��7��������x�J��9��iY6��[Qc�;�l�j�k�cB���_ğr�N����΃@��y1��f��G��G�2"`~�(�R�3O>@U<�.Hb%O4��d�[z���BL���\��*�޾�""�(<��L�}��n8���P]0)"סq_�q��F[0,��n���&: ���h��ʼN��4�Tn(�P=�7�r��Q�ڍx�A022�rc�[�Sz^D���~������X)�{��>�lR�� `I0.FH:���g Y���O.oOs4 ��(��`�"�d�K�,���#�o�D)H_pp*d���Ⱥ�g:+����ڜ�I;#��N�Ǩ�T����"s#���=�C1mj����$f�=��PV]��fH"k�hױ	���	7�W������3�m����с|+�)�ڍ�\�n�D��g��Š5���� �I"fO��1�H8��8��>��b�o�sf"�S�EO��g��� il���}���mXʟ;��sAy�� z1�S�r����ʱ�a���^:2��:,'�(��#�;8��'n�	:�N�! g-^{���Ŋ����F] ����vl���F�����5��q0�G��cv�����لN"����٪; 	��,ZZ�Z��Ǎ:ڨaM��Q�Ak��@D����>O�� /^�����/�&m��q,:ԉ�Z Z7�)R&:�Rhܳ�E4\�����&#�n���ׂ2�_��UOSR}B��M@EP��=���[�鈢F�amΌr�!�c*a��6
�Y+�f��M��b�����f���78&�9	�# x��Q�(�j�b/���	���'3��%�O �Txb�n9W���{f��1�<�)�b�@�1Q�������a��u��<���3ifǔ�f/\?m�5� Q�B��t	�� ~1 ��2}��jp��=K�NE@O��:1���ӑ]�����l/�xT2�Z���ڧ�NJ�&���݃���:�
�V����=0�ތQ��e�Z�Aq�cmAdc���=�:�&6푳��A�bM�u��G���C�*z��O&�ۨ�B�^���Ă���Y�u6�F�|��k�٘�Su�?�V���<��.uۊe�c���ye�?�?�[D�t��
␵;C�Εs��+��vՒ.v4�5  �s���2O���\A���5��;��i�cq�N��NvF*���{6�}�0K��a�:sh�&3�v�L�꘠���׍����Y�-�Y�}lg���Z0��QAЇ�7����_@�;YL�.*�+��A�B_[���{�S`|�獚)=N�P�VN���-�!���ou>(�����������{-� �Pw~�i>,��F�������Oo�����p}����y�/�	�8�<��c.�
�n�V��:p��o���Gy��f�D�أ�葏hv|%�z-�+a�`{֨cE�����Y�{<�V�ӹ]�zĞ��6��R��X�N��go�S�Am�(J*�`���s䗐���gM��⎽�d#X��"WvN�Q�$|�Bo�"В�3�lGeu�T�M���Y6 5�|��.&����B13���*���O��I������t���_���� UtDPG��	���c�Y����k�<��Y��I����bO�5�9S!�:e}Č����R��v�ӈ��Ud�b�Q }����޼�Y���彦�β?q}ag)��~f�K���FJH>�$Eto��l���z�] ,+ۮ)Y�|�xd��F�UcQH�6Z[��,��[vg�&��9b7EC�b:��%c�U�~S�lM�5r��Xģ߶���b���]��8�ٝ�Hǂ"��vF��a�,����������qer������,8��|�(@_��z8f�G�S��n{�X�~i-A�^���G�'� ���Pה|�6_$��L�ct=����E�R%�a)x�7��� ���:��O��h%����x���Q���w�Ty8���.�{,�Q֙�&[&+��ϻdwE�zw|�:�X.�,V� k�-{�8G��8{Ꙇs�^"��p_z?�o�-G�Ԁێ �Ou���W�I9G��9$#�	?)�CQZk�_=�X�f�+�o>8�>���./������2���u�6����6�d?lvi�5����K������~oJ��ŉ LYdҋ���+Ҳ�P��T�I�)&%BY��rWցY�z4sC��l%�h��T~cC�c6G��֯�y�"��b�ݜ��5�+�`�W֦���:���UZ�އ���G
��Q��I�p�RU������m�g���D�0�֛�9���n�^ nJV���YS�&ݭ�
jhs�v��:��\cQ���7�L��B����L�N/�с����?,1w@{l����K02~`�K
�n��;� �m��,�e�`&�X����p�;_�PnÞo*�����������r+�w+uZ�*���4�޲'
J*�Z��s�19x�o1X�s-G�VH��^�0Ԣf��9]�|��+ڞ����/g8�kТd���72P2L������UmF'o޼�o^���u=B� ����#�:w�����/� �sq�$۟�����yv�5��3 yu����}v�`���v��W�-�v4Ga��Օ,�=�)c>�}�|��n��S�f��duX��ȹ�t�� �n�ю��T#[S�yݺ�jʌA1��G����?�,�'�?��Zbmv�����N�!�Y!���j���A>^��۟?���?���U�(��v�A?���=�2�u'+��d��-�!��<��ɠ���kv�Q߿ޛ(��w:��>����2��ف.�����c��r����<I�k)?��#�-�
֨�_�6s��{��ϯ���F����Q�]}���I��֥�+�{�1�[n��
U�nO�5�Sj_�N��5��;�g���~�{�]Q�+�O��l�W�~����������Q�� ���^�(T̒g���L,�S��;�$��CjLn�f+��OvU)5���5�&�:�9�U 3�2���]�u��L�.z��F�pG.��e��f��'�.
+�*X���&е�X6�;�c
*�t�"�����A�\=�WS���;��c�T���H8p�9���q��� �������OG�CT~����m߄*��Զ���ىC�n~ύ�d|�݊*Zm���`���fۆ¨��_A�"���dk�`p��f7 dZ�C�SL���^P��{Y�ο/��;�h:��1�zF�p��k77���HD���y�bE�!�G��;��@�Fw��>"��a��>�����9�G:*J�r���G��F��Ɣ����Ь�F-���=�
�~Zh�$P���S
�Ƽɇ�*�+����6?Y�nT���<P���{d]�����{��/ H|�}�D�	N]�����c>�o�m�y��f)��I!��x�^����qԮA�Cj"i��M�;�K�3s�v��'6&�_8�������бh�u����8��%�@�ֆ����;�VBr+���z��r�/�Ru�Z�w���[5$�6�c�̦5Z��L�՛7���~'�~�;y�����9�\��M�tќ� #�Q��R$�-ȆO�n[�0�w����:��"m_�\2�l��=�X���j
�܉oO��W3s83j�:�PBl��9'?��CQ���7@C��ޜ?���>��e�f[UcB�溨RY��"?$�y������)��h*�UV/�J� �}A$h�{],-ˊ�\��x�
�m9����ɫ>S卾A��|�j:Ν7nE���{��՟,���bUJp(ؠ⸤�1�~X�ڱ�FF5SmA���1���H�T�5���}����ؘehppE�X��@?<���W�q��װn�-@m+�p*�Қ�F��)�FPC{��F��K���~��Zc�w��Y�9h�G�h��auy����1���}�W���]���i���K~��r�왂�+������0�߼����?�����:���s�@�H���GV"+��v�ڰ�3z��?� �@aE��w�>�����( K
�{�ޅo t�����7[��7�B��D|܁�]|��l�F��N��JA���ѹ[�}`�27(�����~��s���B�QdbQ2 �'36�+�[���ύ�@:(�Ldu��'+=�GT22���,���5�����:a��G3���M�vv ���t4��GׂT]d��D6Q���Ú*�.�@��3�w`'dUu�빬�����%����DK��3$�� ��v�+yo>��dPO�8_1�`f�b1�d�w&wuuM�I9�ڲU_�~%''fM��~r�s�i��Z��(��R���5S���$H�!��9Q�C��r���Ɉa42d�w�_�`.��d�����C&��}I�{Z�5`O�+cʉ��Ԗ���F��~Y{�弛@ebũ1�a�;K�x=�X!�m��rYpdCV,J�g�k�0	e �*�Lc3�\��=�d=�dJ�����RƈJmwK��1�ON&.�zF�f(�ڒՃYKK;v��a��j�!��ۊ�LY}�jA��a&, y'�|���m� U>1@�Ե31�&%�����g�Ao/� ����B]A�.�����Q���t��ې�T�6��s(�q'��-�NF?AmBtOAIB]�~��}~"���L��ɚ�f'u� �{z3w�j�� { T'��S��6sD��b�*�a�(@�ֲŸ��N���C�C*��r�^~ US��{�ʢ�;DsNQץ��H�i���c�@��J%�@���*�N��FG� ���p���g�63˥ǅ�N�L�k��<��D��`�/��PBB�:r #:�`��d�HS��M5�%����SU������{�X����)?a^�p'|�y/�,Eէ`�l|��w��	2��P���g�����f��d��S�رa����U>�
�� ����G��H�J7L��!��2#!�D��?�ƀl(k�`V��=���F����X�B_��ǫ���{yv�����:6]mIc�K�+ 'cn�:�Pm���~gY]8�P"C/���(��/�$4��K����=�
)�h.���@渦`
�q�� �9�X��O/���7��W�7_�N�ϞN��.��\??�{2�B3#�7���P�#�Ia+�~V�N6�^�Q:���^}�-6�I��'���PTL�uH���)����G3^f���&ܔR'�����Ux��5�D��4$*E��$�ToP�:b��L���@qϬvc_��ܟ�7�eM�u���8)QK�F:s�c��\�I�C�}��i��`�@ў���l3˾MY{#,�fM*)��ʐ�����V�sTʺM������z��K�qD��|ff�U'�,���cZMOe�8�(Rע~�^V�9�
:Q[R45�A��z����߭tm.��~�,¶���k=X7{
���2��Fb셨�ڠ�7�ܑ���v$�7m<S��o�[s?7��ڨ�hF�U�~�"�M��y��M�^J�/��?.���7rz^���O����869���$w��<�����L��T
�fd��j�v��o�����rr�V>|x+�߿�s�݁6ӟI���ٻw���?�$W
|����^�B�������������f%�1��(�8�Y� �k[�k�����0�Cp�ǿ�]������g8��v��z�u�5V���^��fB�eB021��펙ί
j�F�E����{��_�.����|��+�NΌ�f���s�-�:Ai�Mf�Ԝd���,XK����j���ro��rEG��\u���O���_�yf�;�S�m���n��`��c�rJiW�#a��^a0 >�����l	0���7�}=7���h�"×B�^�
���?�R��������/��� h���O
�R����;h�ӵD�݊�l�槷�'����:A����냿cA�\2�����X6U��2!���(g"T��.���_�\�Hi��8-���|�=*Vmm�2�jc�UL�ೂ�8�C5�b��d���`�~�٫�7�>�+�ѫj��;�x��!콩'n���Z���:��O��ؗ���HOU{�m��ŲmkEŔYV�f�)�(�}|B�#���q1y\�pEAO��Ȼt�r�;��m����+6�����濇2K��({A�����j`$���'T�z�0�O@i��+n�0��e��r*�N�R��43�	����S9��٬��5́�GO��}��UDy�p�:v4 5-���xPQ'�c����!"�� d��@j��j�vpv��¸t���dzP&u�`~�v��d�xd?zsz8לk�S��h����z<�s4D��Yo�\�#�UY���)$X;�Ao�C����4��3�3fpb���"C�Hbn�1�E�z��c�;��F�����9̬������9�.�,B3q��������22Y���9Rt�{�|R�UѾ3�sT[!����w�Z���ɝ>�;?��`��>Wj�W�௎&���D�{(��]1$�?W!����GA��[���O�']������)��Mp||$/_��'"�2�1C��N�^q�q��2������a���'2����������څvĨG��R��YT��Xe�8���'qY�lx����HmgIS��0�8��)&�lU�ށ�;�����c+
7����B ul�,C#�T$�k�����Y��}db����j+�XЁ�@��� A7���FS�{�`i��{��>�/�i�iɂ���O�U���B��-��N�X7�k��,��\]?��j�:��uF�E?'[#+Lg��)�lÑ�DC���ę%Cso���)�����m
!�bE�Oآ`=�b���E	�9��on����'��񽂬+����vhQ;�������e����Ǻ&�����t�F�����N�?�3�t{s'��_	��զQQQP'�sk�5�������5.,����l�eژ[��0X��F[/�`![��������lۄce���3A
�]�����]p�̔d�"��s��]_��u� �˥<;�Շ�<���;:�''����|��]eԵ�δ��w�U�u��X�@�2kю��`��S@�K^+D��'Z6�=�v��Sj��x��"��ڵ��,Lب�{���Q���9�.���Aإs��/c`Q,����Z�I5W�����]}�Y��o�^��,4�.�f�y�eb8���~�JP��u������r���&&��J^+$C�|�;�eI��5=�����A�0Fe�d����=��JdK��;��Q�,R�'��k���Tn�)J�<�߲y�(,J$7��Q�:9>���F�hr��嘑"5��0*P� �9B5�0�l���SF�F���������f� �#�m��cJ��N��G���8�9��gS��Ig_V�T�C��]�)uZ�֎�ї$��_�o1*b����ǂB�É*4]�d?�s�8?V��T��9�vQ:*��b�sO���Eo�)�ڻ!��P�?sc�Y9ec~<�z
��B�b',NgJ�y��TgF(x�ub�{�@j}T�'J��P�ٴ�T��v����n���SIk� �\$��Rj)zR<t�J�a���@�B��6� ������*�x��ڼ	��OL�Ȟ��I��=cd�/� R�(�������j5��f��O�1/��qX�����aFռ�T&�w���!P�Z���{<_�Bg�B�]�����3���J�����3h�f�\{o�t!0@�����?��< A'���|R<z�l쏕��l�H��e����z��y.�'��*o0�5G��Zӹ��Sy����x�J�Oό[roFKL%���<G7᳓�Ӏ��Ho�mGGx���2*@埯��d͍8Y-Y� ��i�����(�=�iP��XR�*�UrZ��������֜��\ٞӗY5��m��y��;oUE�0G�f5����S:<wD�:���t�P7�g�.Y��b�Ǎ�~�/|��g��� AD]K�e0����1*�y,���� ׷��)��'kI��*��\qP��j@��Y_,q��_�#���P{L'ګS�!y}|Lq
.�|R�kd n�ۖ@J��0Q�9bua^3j�~���7�,�.���w�P�C{������WUims�;�{}�������۝�)����[�С�M�Q&P1klnH?�����Cr�umV�4�j�:[W�����j;���Rʟ�S)1��L��	І���l>���'��;i�;���������|��=���D�T<D��F:땙C�&�~�c�NoeV㵺�	��V�<���g,�r�4j[��J�dL�����S+1_�y��FA��<�Ǭ���Jk		�]�A���f@�'J
&m��8֠~#��Nnt޼�i��������{�������5��t��ŧ������|�,#&2^��|��) +h�n	F.M��}3��J�d8�!��w^{%v>��c�v ��,�xb,0H�H�w�N0K� Pg����+� �ѷ�E�b�J&+2Uv�y �F���d�ƹscݿ��<��xo�J�@�mt��R��6H�Fv��⬲���~�F�=hĊ֪��39N��1��}D��i���'<Z � &�B��=�sj�E�_C���>D�?�8D��W�B��v�����_����H�v�ĸ!�F�4�?�(w�2��<�F�L��Ky��R^>?��g�QPC�^=(���{3�Gt��cr�tgr�8_DTB~�h3we6������sF`Q��"�K
M�*��r�{�6{�O;9�e�S#GN�$6�1���F�N����
�ɀ\�Z�vos*k����"],�Zh��"W40���~�⦌�z11��p��Y!A�h��e�'o�g���q����*�$�:�(�?��9ԸF��'/k ��ѭÏ�'c�&�h��<����R�\ylD���(�8�6�W����2�it(N�eޗ���ʚї�ā�룟N�v�6ꘊ�1u&���9_y�cSg�@E8�qoz�P��`<���7�&[ ���Q�pH-؅���b.'��|)��-�ļ��BW*u~	`�#P���Oaz��d^���gU���5g�#oז��'ҹ��t����ζ���t�^E6Ν_��`���j~M ��'*qu��0G<8d�,�2�)�4	 a�����hӝ����銵G�ASm��%�6ǘa�-�H'5��M:|#�+sK��6�Olߧ����B%ˢq�|r݀%�����k��w�{��]��ku�����^�[�ɂ���ł��F;o(lf�l;���֪T&!MUQ�{hJ���`~@�J���h���\�Wl6�*&q�o��X��.W+�I h��%�U��ĩ&��"8,����&Ң�e��M��N,c��:؛Iσڱ��;��P�N7e��*2��ʢ��@�� �G�sԟ�� ����W��[�xjHJB�1Z�P�̚�5hE�a�
���RT��8���!�0���XV �Y��u�(L�Z2�H��ؒDV�h��k���ƚ�r�d�;g �ֈ�Of�w:^�-��T�\Ȳ�6^�gC�MeZ�:$)�p}T�����[���񄴸�
��,`�D6q���dM�֚��:�>"���&5CS�wײ�>H���NA�Շw:��	ꋝ� Dq��{U�����ܶ��M�9(���� d�+��6ՠ��)Ab��÷�8��� .\6>K�����^|'�d�샯�A5��N�Ć+�Z���j�2�Z���k���+����`��n �e��P[=�i�� g&�Y�K�'BJ�Τ�͙j�X j���w�YW#$l��s�HLdJl���6��gQD�!�.��g��O��F9���)�@��H9�ݨ[��� ��D���߽:[d��C�Q�e�W��[�3���0FN�nU�nf,�6��|*'�
�./���sy��>d�8Sp��fV�>1�f�ƪL]�d�ے��m�N��E$��"��gO�P�"=���)ŴӉ�ӎ`�W պ�<_:s$��@�^zݠd#�z�@�gM� ��Sٝ��$��v��YsKI�n�x�Q��hR[�7_��[6��(�ܡ��d�_?���Lrr㈉��9.�u��?`�/K�L��D� r���UF��b�c��a�?��嫟B��s}q���o�1�r�z��xr�t�W��a��&�6�^�?T_�8�Ӆj�v�r*N�s������)�A4
�D�{��{m� $��#kI�ȊX����o�`x8��a�0Phۢ�p�d��F�	dݡ��3�q�;����7r�N��ٹ���q'9/�F�Jf��k��0�����v5��~0�F(V�?0��"�10]+҄k��u������S�7�=� �^�Rm��D��}o4���.�B��� +�Kq�\�Y�(�:3���bCҜ'��`��y���K�V��qC��V&�K�Dv� ��ug�HR9�k���Zg�ڹ'iCsL�������څ��`BMYz����Hu���5��}/���\�n��f�:��nF!�^|z�Mx+k"�}uh�R\�R���/�_s?&����33"z�������٩<�x��$��g۔)��@��S�5���
zjOH�Ē6���ɦ����nvE�A�*�u	��s��a�.�"��C����h$ h[�`�?C� ��l~�������r͊�BK�о��z�5�4��a}�. �HQ�L��g�S�z�{��}��yd��l�Y��X��g��I�?����@��`B��b`���)��N.�SoIc�2X ��<�~���m�^��QX2��)�ǉ��NP4	��a��;�c~��V<h�%@���d��zݔ�gS�����bf�<K���X��X"���Y��[m���= �V���5�:e�2x�x�����ń�K�^����u���B�t������ +9['��-�	dz�'?��$�}F�(���T��R
⛌r�#�*j��%c���m�{����d�rA�1}n���0�`�al��m�-�pv�#�J2�r,|g+A��9��pP[�{�uq&(, �r݄Q��֋F_�z,�&���dbH�G�����5��O�"�NC��2ZC�Tq��\���p^�/y�������(h�c���7��� B�\y4���r���~ɤ�A��ڙ�E߭%`�FK @�(e���~)5R�sS�Bϗfjz*�5+58�����+�����ͥ�z�L�_��Ѣ6.j�30�@�ʞT��4��"TCAUA��zo��w���x��[L ��B��T;m)�=��و�k����
Z�?������������=���W�t��rw����n������,��[���"�`���H�D8�U��ފOA��2Oe�kK뛃]2[9��yt��ԯQ�>�0l2Dh�؍L�`�"C����_�ȣ5p`2m���K����2X�(�jVl�T-E�s�^d�7u��1IO7���gL����cgѤ!��͛7�6^���m�@���t��~��c�vs������nd{l3l��ʌ2C�XF��jYp*v Zj��1Z��>�)\��Ӳ3���ŉ��g2eVc�"L��X_8
�1�*��6U��˜{\�:�9�-&��\7��Dm"��_��ǐ�q��D�٩95��rΆd<��خSZ��ܛ:�	\@���S���vԛX�~突�����wlO����)*S���(߻�)���@�%鋖�a�kD��dmrA�E'�L=H=&�n	{���]�<IQ������<Ƶ� Ou�f��{�z�
[��b�� h:��j-�7;y\"��ń�$}8�������C�+����;�(AC(���T�e��@ ����2�S�q���5��:�'3*l`.%��P��׆��`�@����ޟh{3��np�IQw+�0�`�N�|\B�tkv8��	�}KY�-?���)�H-��!Qz�F&���'�Ί��Ђ@I4C����=2�[�ǝ�{w�:�T��!����4
JD������A�5Pptg��4�� ����A/�o��Z�������K����!�=�VT�<�����0�=���P$��� [L�X�z�b�u6�Dj�i\R�=�ؤ���o�BR���)�b�Of��Y��8��;~���k�w;S�e[�ɬ􌥤�������΁����,)�������~g>&=���d���]m���Z��[\�VSP�Vp�Z#G���q`Բl�8������)�<�"�Uz�7��Y.�v�Qط�+�ѝ��}��_� �Hd�a��X�[g�����Ye�-wVP�$�zok�r�d�t,� X��vR�ٹ7lpʬ>��1�0�C_��M�i��7)k
������F��dFr�0R�a�2!�:,��R�	��Z��8@i8>f�Q�Ψ&���~2���z3�t�q����hY+���'��Ɐ1�6��z�@c�$�K 7{��<{��Xk���S��=�$2Wh�V�<�5uU�	�&�>nGs9>=���S�|�L^������������Ζ������WflG�.Ԑ����������t"��eX�}���P�Z/�s� ����d�ک��Ŏ�0�6�-$b�Rd�h�������:���S}��>^�����������{y��&X���[����EVѤ�'����5�S���U��ϖE0.�-�쑭�?����__�����������j����{��'t���|x�\V�6%�`P`�x~���̏e��s�s`kT,f#hLk��o_�Eiѕ����6*{
��9W!���_�w�}'_������_*��� ��rY�{NA���A�#Г��}P�2 j|��(ًŬ��)�P�kRoզ.�2o2|C��ğ����͑�+ȺԵqL[ ^{a�I���32XA%��M�M6�'7{�D�.6nryw������ �_1&��Q��RP-���0>�`����y_�}��Ӣ�A݋���֧�7L��p�F�p�[o�s_
��7׮&'p
�@4ή�(:w+�,��R�U�}r�{��izF��5F[4)�$G�a|����9i��v���=$��, ��2�&���v�l������J�˲R���1�mj*嵽:���_D�� �i��f�'��v���`+l|�"d+Wv�mN��L ��n`��C}頝�<F��b���5����"ej��ԇ��2���6��<[v�+�Yo��$���8ǡ���H�mK�r�̄yK��U-��yCt���&�ߥP�B8%X���{P�@�7g!���b'�_<��ť�~�(K��`� K���2+�
~Vbh�=s�{6=F�2^���Wۖ�,z�}��o����^^\���Q��]��C�~>?��T�]�M��f��4V���L��'(6C�B7����F�k�j�h�p���p��ɳFֺF*��Wm>kH}�zޢ��5�&Y�ɥ�;��%8Z֞6�2�m��������4s�Kȸ#���k� �� 6�y�W`�۬t?]�5*vC��Y;Kۯê>n�r��n���\e7y�� ��O�K R<����@����u�yZ�{�� -����$#*�AI�Ƴ��c1��;JM����=C�B�6E-��tn��� ��i�9�zk��X��iwIF�j(�F� gI�ގ��쓰��	�9^.�LG��,�}�P���d�"�z��P�h�'r�fz���a�^�z��\��8�e|����^T�խq����'�b��U��wiR�7�Ɣ��;?��Ǝ�1AdԴ�j�&�eve�]s��w+�۲�0j����kI��g	�ŝXy���DE � ��]�`]�������XNO� ��D�1�(�b���=Z�ǽHn4!��L�n�+k�k@��K��y�^dJ�����1[�I=ؐ�PUj�7Ɵo{S���
GAch��,�nL:��Of�\-���fǼ�����B�B�� ��޵��ot�7�4�<��Μ,-q����~jTxr����a6�Z2�6W�
	�����_c*����3h��?�G���W�Gp�H�%���Xt��ɟ~}�P)�)����H��-�LA��A�����n���R?�*���g��	�.zs�h���6F��o�PO���ꫯ��=�̾4�ޑn�G�/�1��Ӹ�ml�ݎt�	!z^�Ōv6~9�(�Bv�9����W{�%���=�@�e��Jag����q����� �!8*�B��4pt������&���"A��@uY5zXE�3iX��^�Q΢��
WCo<�� 2�5.㜝�Og�v0���11z��\���-ֲ$��,�h�D���,�eMĥ���<�P��Z	q�S���ԧ)Sh�ޒE� ���E�#-�cR�����zd	�Y7w8��sd����0��ڴ�����zP���u����1r����怽q,�l^�*�<���'�G�?Q3�Y��z#�-E�O���f��P�5yo��>�	�Ud��h��&Ԧ�s����3l��Wy ;����S�}� $O�1Z�e�6(���{�K�+�I���2K*�ܒN��qN�O^�\�d�6���D��g�@���n)��*�\9j�'ڞ?�;��k�S����9�{a�e��������Q;������A ��d/k=�>��^��7�+̧�d0QHm��QP%K�]�����W��{��'�@�fK����B����k\����XR�#�Ƽ��X_˸���� 86��̖-����~�vC�5gb� ��l���>֔۷��TD�
b)A����}Q�w�\�1!��Q#�a�ٛ|Qp�ׁURT?c>FK�U�N���E���+��Fq���w�k4�.ZA*y6q��eV�S�'�
�WS9��c��3V��:�&�D����ёay�(����&8�48��h�i���d�� ��ܭi���9d!�y~��|��Z���䄀jqdM�֫�dp�^�x�����a�SA*��U�=BalP sO� �=@�p�^��Z��=*�ҋO�V���S�t���{��A���"�w�@�k��B/���f�d1��Ts>���'�\��W�.���K5�Gl@wt4#�yF�@z+�4("x����:f$d��(�'<�;O��#�-NK�]t�"��?��y�@�!=qo}(��3���.��)r�Z��bX�
Q%Dd���N�r~:�T�^���P!᜚3c��q5�Ĭ��:�]i��hNޣMSP<v�"Υ��y�1Ǹa�C�_(��L`���R:D���)�gr��J���?h�bDu����If�q�Q�_8�/���������{ �(�GT���
�0���ȶW.6`kջ��sP(��� �<b�N�=Dao.//����!DCN���b1���|��˿�����=���T�&ժ䓻�*gSQ��཮�r8v��������W�=g�	g!�n{�g����)%xt���/O������O30����/�Дcr�к�Ao=є�Rr5"��ʵۜ�l|��b׫<�CA	p!�<�M�eHg�����,d������嫫P�uF�;��o�қu��~,�j����	�R��舱�>+�Yf1*�U�$%g1�z4�b`�rY��Z���DFO�Hr�{o(�ZM)�VG�CQPo�j��ۻ� Z�]����S��4p.�Cx�!��R睉 �i=�S=&s�ΡŜ��"`rߡ���>��{��aB��A��m�1�!��KF6E?��Ё٣��s�C�S�{�|���Y��#m��}"��Iu��P���:hGK�ز�q��8��gTM����.k��\ ������s�3��~+���k��%�3h��CD$��%�(��^ d�(K�v���ĸ5#� �;jL̂0�XQY�Ek4��[��u�h��-hL3�l|�IC���
��Z:�FJ&�er���>�ln���.Ȇ�UOќd�2,؍L9�_,�hx�=����Ֆ����9l����t���i_]y�t��q�/�d��QuoT7�p�n>�f���BP��M�V3��,���Ϭ�6�[<�5���ux2����!���ߐ�oĩ�&F��1���fk�>��V�DhUcO��Z�_���13lmc�� �⁒V�B���*���
�r_ф�i8%������ش�o�TeB���X���r̽����x�X(x~��o����^~��+y��� ���E������0��9����/�	�,|�}����8��UR�W���������*Ǹ�W����F���h�&n�������pL.�mT�/~n�,�5AlR��$zb�/G#G
�������K��z}� �RAl�1�3�kQ��i�K��f5�T4&�%��"E���8�p��@g�'1B&�u�^9}��L�R�o˾V�3ņ����� ����@�o�<���":��d��9�R���B�)�\>���#��;�s��0�F}���^�vB*�,J�2L��{mR-���<�WpJ���RVt����&��xf4_/i�����_��t|ί�3@Ir؉<L��H�\���Ύ(��"Bj�A뫽W�Q@"c5P#(�$�(�y*r�~f#� B��;xτ�3����x?���<��T3�"8lY��� }
El����R�����~��)��* �e%���@�I;fq�6����%jZ@F}f��:�|v{^����¢_r�G �7�x5����8Ŀ�G�_�9p�^M>/<CTU�O8)+��|��{�:�J�}tj}_�O���Tl�k?�ʝ^;�{�֓����ǹ���q=ք=�j�G[8`@Q\��3����c�k�(1 �61��&�e`ҩb��;]��<�������� kX�=� H��T�����L��Nq+7w[�x����=배Gt���2���+����)Qƺ��{�+�����K�"�i ����QgǠ��k�I���j��m��Ojy�+(�ݐ�h�j������8!�(�-��!}�Z-�W�WN���K�Y��r��3<X�15�{P��Hk��FM&��K��De�t���,�MK�
��x�XCF�_��J_/(��x!���;�A��:j=S��]�Z �)�4R`uЈ@�sՂ%`3�y0�6\����[�������kvݕS�S
�K)�mLl��0l�T�L�)W�ͱ{a3?���׃U��������=M���.�n��A�z��Ei4䙎%z�e��7�� %3N�h̍���\nv4�5 C����	���b����څT���l�p�LJ�BL�/�%(����n8���fZ��a6u��]�I�d�Q�5�fq>
bJŇj�x�xO��}�
�J��C�AO�ڼ�vM�������Q{���s�'�\Q��]��i �)�K�uJ"}��gA��s:H�Ή�q�
mi f�#y��|��o������V���1)�(����b��J(�pv~�Ƹ�p֧5=�z�L	z:PТ�>0�3R���C�c�cT`j��,%aw:���Lf	�z:���["��a������'Ql���m��DQ�>��}��7�Y�E\,*5��Z�G�Re�(F����[
`��O���X�x�B���|�����%�ƱN��JՐ����F�D���>U`�^�����Z��!1�Mk�{믑<R��ߞ7S�������gl�g��He-���e�FϑvAť�Z�f�('EPP��]v4�8N]�9��P���^7���.�}��5���)V��,����h/��'��N�����/�3�N'��{��E���*��&�@����*�Nݜ�D�,S��@R�*X�ٸ�h;�GEP�g�"���Yէ�~�;�~�jd4R6ޯѱ��J�ZN}1:�s���4٨��e�(��QE�D_9�ö�X�h��@�%͟�o]�-Kp�ms�恹� BvEɚ���7!g�@m�Z�׍Z����S�F�;����qa{�Im��p^�z,�ҙ��%�l�:gK���=k*~-���B��(���_0C��%�O6B/Cg�x�i���B-��"u���Ok�m\K��`��J�P�ˬ�B�z��i���t��e�s��fI��j+��T:d�����a/'^g�Z�c
���WR�kG���ܻ=��a#m[��0��عxĚ�w��N�;r�"�������k���57��Mڼ�ё@�m�K��=�DX�7Y{}8���;d*�;|H?�y��tZd������z����^X'�^�PP�u��cO�֋�unR~��T�v��a|�`fT6�	��������٣tG(k��w���Bx���2}�C6�D��I��q�T��C���	���[����(���z��bq!�f�,�nov�㻝���ɝ�˭�]��y+�L�:+*�� � ��_G���BO5��`M'uM�M��a�̶��S{�#�LxO�9��}�`f��Ǉ5i�WP��	)`���-�hg�x�]�3�T�MIx��Q	���R��:O��l)w�
�օ�����y���9��� o���_C�`π���)�y�7��9�����kA�){aJ:����+f�����wo"�=��{/j{/��C -{NO�..��;Oh�`�t�����Q�m���M�=T4��U�ǼY��?Zb~�KS�������wP���Y����f
��)�[�1Mi����Շ��x#�
����u��Α�H��6�3�̙ ��Dk�	�����癢�}e���S.��7[�M�"К���ն���Tl�V�	�S�h�
�U��#4{k"��Iۑ�|� <_G?Q����#fې�k ��M�`G�j�S�FMkK�*����:����>l���\�k,} �q���s�M�,d�f��],��V�A�ւ�p�Q/���~5�0�� �mG���*�s�}[�mD�30E�b�s�{�����[
V�Pů��h��}���F ��Db���R�=|��5�k�y"p��lq��^690��q4<���t���'�:�OJ�>��A!�*78�T[A=������ȿ�ۿ����
����FH01�����Y�AHi���}##���,聣�N�������fHu&?�X��p<%6��������6�֣�HGz�a�~Y���Bb�]�7H�8x�7��0I��E�������卂-]��-��/)���������J3hn�0N�.�χ%;����d`T�/�XH>m;����r��n+e�l5'}o5�~� ��R�ɮ1��0��8QA��t>[ AY
E� ��Ӄ�5�V�z=>��fw�N�178��k��hO��/�l{Z{J���c�o���f�xO�l���9�enl���=;�~b��"�X �+U��e^����FY������8���N�����A�;�VC�}tM�F�{�N"8�>�A�Fp){�h��~�
�^/�a4�f�o���� uP �~�Ѐ�uww+���rrz�����@�܍�9�T}��2�ޟ�y�iq�}��b�ʜ)D���H��8�)� �]P� �P�@��հwt�Lb"ш������emw%=|��G5�i��z���_K9�R"W��X���B�n���#�WILz�9�ܠ���,�p`��}�+F��Y<B��䔲����8>�=m�B�����*�聞�+ �60G7�:yw�׶ٻ��}�K-��l�x�������ŉg���;�V�6���ۏ�pvˢ��0s߳$%	�dx�?�H�����#�6p�ՠ+u�^ɺ��欗��N��������:��m�5 �>�_�2&������C�@������a����-����Q��#sn�fv���>������xG��g�B��x!���N�c�3 ���/2뫕��1�e�.��$(�^��vg}Jf��?ko��H�$	��; �W\�Y���N�������0��U�W�<@pw[UsgdVU�~���d� �n�����(� J{��Be��&E��`�i��@�z�M>ߔ��Z��f&څ�c�޺ ��Y��)UQn��.l�k�Y(������Fr�͡�$�ڎ�~@2@�x-D�����f��30�P(D�������^ �@�[��������s��7h�����X^��/�K)ͽ�UL\�f�A�K�K�2�5��f?{�ˉ���=(o���XWK?����BbE� F�@��i����`����]يZ�e7���m(��VV8�w�8U��w�a-Rzl7�g~^W����
ۉ2 ��(!т�<���#�x�p�R�� b�|�c;<8&h�����U�M?��c�l���Z�n|r�Mu���5�n��(0�U{�A�s�W����v$@p���L���|�3����_b5��K�������6��`@��fގ�S��ZK�G��i@9	��ݷ�ٟ��*�"���N(kE�q(A��g���px�I�D4� �Q8?[������������֦L��T|7�����Yp�k�P"�C3�����(M�۴A�TS̃2�g'\=+@�=yrn�'l�G� ����B`b�Pix[��/ �h�T-"*����HQ�EB�)x���J���R��O�]G��x!aJ��=GJ1ZS[✆\�[���46o�-�8j�nnnY���;�`�l൬V]ٸ�<��m�7���Fs�
	g�-A� d�-��4H�J�@�jK��H���-�<����w�uU͝'�.��7�^_��6��:�zg�e���nr����7wG�Ȃ�T�_����Q/�{K��Wiګ3g����!���ݍ䒋SB�pR=��=�����,(:5�t� ,��E�=�1������vv^n�`9X�(g!��sm�f"��'͵�j� �I�#mԪ�Hۨ�)#ޭ��Fe*$��&��C�b���I�詊G�^}�U��aZO^c;VZ���/.6���٣��lbs�����w��{��&
�׉�N����^g!�Ng�wت�"�(R (��G���а����N��<;b���Ș�?8�eu^�ߞ��f��j���kF�!�}{sm�W��sO .���z�*t̄�j\�x�L�X��A�F2㌨�R<D�zo�$�Q�36��b���_���LϏ���p���b���j=�|�?��,��-Z���-������v}�a8� X��:xZhȌ5NK[�+~K:�Uëj��
��H4�>I$	��6̗�k�����{�-��R��q����f����o����@=�4�O-W-�<�j^X���a�#\�������!H���œ'2��ˌʍ�D��¥�׫Z�W���D�W�s<���{�����l�l����;{��--�����Y 2�����괰����s�Ө��vP���|(��fJ�}�����&Z�9I_�Z ��f��t���tY��\ǆBF;f�v����"UY�g�����#k�s=��|��
ڵb����_h��?@ufY����
��@��i�@z~�<� UZ�"P��Ulb�,�`�n2����/�!�Gk"��ֳl��n��V����lpMkt�"��D-�	�$~r�2�ծU�<��D�s����
��{\����5P}���̀��vY�~}}Wƽw@�x��.�&���)�_�0z�\�~$*g�͂�a���#c�kC�`{����I��sC��'UR���O� <R ,�H1tcY�ɣ
M:��Y��v��w������Eqz�����Y�����P�� %2�L76d4�T���T,��c&�R�2��&�����|�f��i{�M�&�Ҳ��:�Q(�:c�	h�a�u
�8W_`�RP"���9���|����c{��ܞ���&i�@a�~wg���E9������ȼ|����{�Ĺ^n�P!��hMm2����r�G��a�����,�7�\6��J3�Q�x�@��[�^��3�2��4[*���)y8���wtzك�:(�{n��vG����2(<���Ég=X/'Z�0�$N�(E�e���[��X뎄;1_9��߉��l5��+b�+���s��b�#���0��;��:�4et�b�ړ�Z*N�������~Ĳ����@�z:Y�JLNt�NO�@�:C��(kH�na͌%���Xv�ӏ^k�&�Y�S#n�ͺ���j������+�{}��>~�`Ϟ?�gO����"{1��:��r>�~L
o��`2q[4*���'i���!*ۨ!x�����@B��};���[�m�>(`t-!���a�co������袏C�գ�Ms�w�mfVE�+E{��j��/�������Ri�[y�[㸡_Ϯ�L?�(�F���>5_<ynO���ӳ��P�����ߣ�3?cq@��3 qó}J�.������������/l]}�X��'[�ݖ��*R����I�d$h-�B�6NOi����<�ݚ��DӺQ���Ȫ��05 b����Y߿�d}*ʮ���b� d�����UX����*N��Y�vD�l��-5"P��T�NM���r��6ov�M�8��}���k.��%����0(w_ ѡ"�pj��{��) ����!���O�5����H!���l�΢W��B�^�X#���E�-�A��s`�6�W��G����=~Hm:U�����Ÿb\�4��o��*�ߺ���?�Ͽ���~���}�Pl����A�0��� d)��������2��*���o�l��|Χ���/?�/�����NG�����EǌU,�{,8���א�G}؆A�Č�8sB�s�[0��ځ�
(�[dJ�L���T��Ӑ�̪�%�Y���� �-�a(Q�8)�������!t�Y��-�FqM⼄)����#K>I�l��P�����8z���>O�ϙ_;�3_�uEDe���:- 봀-H�/�;�ڹ�BC��8���Y V�� Y��!����aK�RF{t/�sa�%������Xp%ʼ0�=0x�0/��`�hĢ�;��yՈ��}[~�kt�v�H�|�շ�'U3WJ+�j�@�!Q牡K��������1����4�t��݂O_6���1r���<0K�ȡ&��by��M*HkB�!E�g�*�wG#:dW��YU����>h������ �	@5��	di��$B����,6NPds��\�wOS��<AE�@�:=A��R���i�����ȳoe�$���Hj2F{�W��gd�s���!vFidf���j#xǃ��39�E#�Q���M#E�Dհ��[W�����g!��B�ԁuv=��w�f��Ȳ:t��[D�*������fӲ�&~Q �����H��fd��f�m:��霈�����5Q��IT�����4��+Kkk�7Z�#�̦�(w��DC_��u]�x�_=�?�ƪ���*�I�=����x��ִ�o���Zi�d����Ve_�H����ý�Iu�Lɷ�o��eNwqW��c��s��!**��s5P���s[W尺g�Y����<­@�����&kv��#)�b��l|a��(#��J4��X�]�`@�zJ5�H�Z�����bc�W�����n����B��A��ض".>v����ү��U��W�	hW��f�;��a]�7������=\�����[��4��" �FV��*�gAv9�Ϟ<��/^�7/��Ͽ���3�k���2���k��)�?�]Sq����ഫ#�?>���/P���}.��Çwp�����m�o����%[���M`�ؒ�^˃(|B���6�7�Y_[:#/u�;�� Z�|�o;ӿ1�>?���)Ş֩6�.&/���*��DV�8������Kd��v���/�&��"�o� ����c������T:�Q�2�qvF��a����<$G�FwF��I�����A k}Z:D&�@/�[P�V�۠RM��:V+ 5�Z9XU=��;f�$T��ڕjF�-��[ڬ����r⅝_\�m���ϗ�Ŀ}����Ȩ��cM�-s�@�rF܉d�`9�$�Y��|���T����՗��>ڛw��4��p0��x
�3�Pm�ZȦ�}A�۩=.�J{<�vW���w;���؟�t^���d�	��,��r}t�N�s�.b�TEՃ�L}/�d�a�ŀh������^|��N�d�3,��T5�iK�E��a�1��g?K"��%�"���Q{�����8?!��Y�HL��\�l$�����)���/��n�[�k��?)j��+��%`{�Q�Y��=�[B���}0n�t��}`)������ٹSx����������Z6�N
 {���R=���@���5�dr���M�����w��ly���5ۥХ�y��x��3߲j��<2��P�{HA�ՑA�@�o��(��%�!m�kPK�'���W���|*���Q7����Z�jĦ�F��Ii�jT69ؒ�hn��qʩ���׃�ajD\3v3�4ٯ�"�@���Ӕ�E���������8d�,�f6��+@�ķ�6�^��f���h��%�V�@���`���6/�u����s������pѝ�l��C�z�;(�y�Q��GI�e8�x�~T4��~Bo@M
���Y�Fo�W��f�jM8＿~�Z������2�Mj�`��H&Xo���f���1��@<"^��N��`�����:E��su>�����C������A�nΉ03[QV;��:Kq�%/��W�zn<iV����Rp =J�������b�~�LӿF��E_?\U������xD�x2,�?�}�}�R5\����U�1�ìoͶR벃��師|v���5C\�x�P�P����8�TC+d��N�^1�蹂5�P-�Q��|��q�|�˄%w08'�M<�Gg(KEɱ�v�ݖ8j�5$%�}W�h�cZ�AX?]��/��w#��8m�>=8���=��[nK]Z:2a>���n��E@��湀���}�5pY��T�d�0DG!���=}�<}^~��x�����N,}x���GK�3@_=���)`�WC��G�ٷ�?�g�_\���ݐFxE*����p���Rs�*�V<�������v���YX��4���NN�o�#K�4u��g	x�{tPJ�)/���Uk�*���͎��_n��{��.!�5��Al�&(�`�Q�4���:F��~'{�z���s=-���jlF��Y�s�1G �Β�����9%�����}�^S��/_��������ʀj]㙙e���R9$��vD����#�t��{�c��-�����s���������=��vrT���)�����޽}�L��?7��1�!
YUq�2�ȋu$J�@U�'P!�1,��PK��=k�n�X�6�.6����f�j]p:��w��m
vDH�{���;�Ug����޾}k�߼�?|{nϟ]賲�� ���X�3e�:g��)EY'ґ�W�{���_��W�SrM��6���S���gg*�؃4c��3�&�GU�@V쬺e��p�+P1?,�^Ma��@8k M��z1J�����w)��E�������k��d}G��{�S��VK�\5m�-�\��X��8<� �Z8��~������"�M�^�1���3U���ey�z�)~�,�\�8EYL��ϙ����=亟$W߸/2�d�l�WZ��G�����p^�s�Q��f�-=��[sA��Mnlռ�����������Ϭ���qrz�%$���%2��]��M�lѸ$��S""Vu��)���2��A�D��p�v�W?�Q��\�T��8�z��"�6(���Q�F�c�����d�~(Q4j�Bμ��ES �,����e͛�����	-�� ��R3>Po�A:�]��G��=�Lc�%uqgĹ�^�W�_��%�L�IIJg;�Ħ׹׵�x��igY��T����Q/��UT��(��(M��墍֭"S#�*�.W�_��r)���#���Y�肭+��	3�`PXm��N����Ѥ�F��~D�������\te8�xd��A����гWU\�ѓ���t��Z��gl��_=&��!��k�Ș���V�&���Ĳ߮F$��#�Ը���a�BXƬf�߯ֈj�+����꫆��}��8<:b!.F=�n��Y8���?k�C�7�A!	 �  s��j;��u;[�ذQN��a&���>_�����!���?ޒe��q��V?���[π��G�ۺ��9���?�l��y�Fj��t��	�f������d��:w4SG���HP��b�b����{�������Y���EZ{H���� ���p�ͭ�^�W�5��$9;TC-c���,�r��vsxlGG�t} ����;:mm���:��g^dޮQ����r>^G丼�QY/;����\��:�qM1�Z?_�������ǯ�&�]�ֈ�׍Gv���?\ۧˏ���s*wv{�)�®|?���f�m�s��^�j[�M�ST�A�a��M�n(�2S084�'�j4��8̢TA��/w::�1~Q/A��/��/ol�&���~�����/���[�]�1X;I�e�W���Ds�>�I(��O�Eq�N�Ȯ_�\�1�e@��NO����L�B���v�ǔ��qd�uQ?~$l����w�Ȋ�����+!�(����Y{�)׵w ��ױGT9��l�ckV��vk�E�Og�b����.	Z��xi��׫��HZ.h��������5�z6 �]�.Z�=���}D؋��.ݳɊ#��9����w�v�Ȉ	ug��I�u�}Q�zڢ8wG�� r�_H��.�?��uָ/�=@Oq�$���uM��u�wſA[���JUTmR�������o��#;�l�(�9���A� K�L�g׾Xo
���@6��/�.�r\�� <�� >�� ڨ�1Ȅ�;���S|�|�<�*XCW�����俟J6��a7���,�K�S�q�'
3�;~�_�`���Q��"0TY�踢�2(J�a�C����Trʩ^~~}}m���ŀ\�۷���Sa|c/_�,��E���䣅��/��P�n<S���I�4����ੈl>��(��@k�gg�������-��  ��IDATن�N�7�%?��q\ üw'3��Y+OsGCJ>^�JE����N��I1�����.��(����yd�tR#��T��Yn]�]�����Y��ӑ#�s4�78u�j����;�N1�8��N���D��d�׉XHd�����V��<�����kAg�Q����(�NJr���,�  ��?���#�=�'-dp��c"�z�,�'f#��jV� @�8��]�-��ot������5�S�6�*�sd�`�7����8H�s�KR�`����4�)�����<0&��=����~f,�{���fA�S�}RK�ov�BɁLv
k?=E�<�&A����~z�NTDi���ňrb���Q�w�pO���<T�P��"���C0�C�$*)I�q�H�Mi:�飂��ѣh�˖<S][j�|��Ȟ�հ���X���~uc�_��m��w�3"����ow<���^?���C�9���5�h�3�� �LMN��&�=�@'2M���V�S�k��:�	RP���<,��������dA�b��(fg�{+:N��M �0��!��5e;&$�Y��/2��ST�2�l�~G��+P��i!��� �Y,�F-�8^�K�#]��謌Eq@��X�I��c݀:�<05CI���=@+T��c�Q���� ��.`곽{��޼}ko�}�O��է;��B��(׾C���O�l�=RY��P	
Pύ�X�a�Pٍ)�Su�ӋX������Z���Q=�����K��޼}g�����!�^���/?����#�Y�1c��j�S�m.�E��*T�q�؇�8��@���T]�1�u{s[ �'���(���������y�'l5�A��ةo^�F�^u�府mW���;�K�֊;��F5��O~���<F�Z� ��7{T����}$�V�@��=��(��u\!�L���-̮��}��C�Y�cٶ�N��V���~Z�l��Nʞ:?=�C�sI�����'����jA�52W-?�_�>�DP2X��g&��ND����J۪��ln��R���C�y�'�Y�J�����-�Y,ή�B5�M�}�cxPe&,�<��z��)��2�����ƃÍ���>mi���޹�mxx���#���VNr�s*�w�H�rɒ��r��=�qP��k6��1�E�+�����g�L%~ό��rew��z�R�ErQ� ��,��d�3윲U�3"�k�-K�U.3A3�P|l�^ ��c'��i���8�AF -����a�@���td'��!�=�L��Q2_���o�����8������D��(,W�t�!Ít-h3w�"B'�)b�v��H�if((g��e/)�R	#3?=~����G�����4�)z̍�'�E�G��h��aZ��h�ֳhgq'�eۗTsY��%��ϟhA�"	*���s��c{�\�����Ɲ�l�yZl��.��K��7��C�p;2��Pn��mT=����c��,P���d�_���є��|$5&;�K�JϨى�{�?s�YQcI�vrL {�B���;��B�׊�^���ih4����a�.���4*F�6��RmP�����ܸa1�3V9F����1]���Ӛ����$Rw�h���&�"%���]�Cjd	��3�U�	���#&�����d@�F�3^T
I]��Dh!۴v=��?���R4z�Z �i������ak�j`Q�9��g�M�/��G5��"2Ĳx��JBU[_-"�leR:d_#ԇB�d%M�1��&y�J�j朐�mj��s5x�xmD4�;��՘��`1R�� ��Ԅ�A���5\7�w���[����V@���r�F����s����+���1s���n�V��2� @uelFo:	I�+C��QȪw�|���A�j�V ���[N`Ȑ}|�셽�������vr��ش�*Z��Ӝ����oK�P�Yv�����{
���p��,*�.j't�b����0��{����X�RQ [u[����{\��iq2O�_i��N|v�}�V�vG�sJo�h�ߩ�?��;������EZ�������~��^�~eo_������g6k�k	rɐ�+`0�3P����� d�˾@6�
���}��|^��!�x#�
~�z9p(���ZfO:9��������Ȃx����YK���{��ǟ���^�B]sZ^�t���C�b\p!��jd\��j���^��ؖ�����uxؗ�~��٨�.����s���C��j�� ��6�sf��MA�ƴ��c��ټӎg!���@y.���� �6�^����x�!28zQ�R�P5eدN5U�w�`��U�=�Ծ{�� �S[��7�M=����iy�mͲ�Y�j�;��Ծ��c�B�d���썳T`k�2�ۇ���J��}oJ�������Cv�;f��S� �����,�����.ɼ�ٙ�,����c`�M5MȂ���`
2�G���כg���lV�*=
Y|�c�d�Vm�#�k��['���i�P�Q����E�`�X�:���X�-�#���L��2�\�(05��@�-{p��̶��^[����!�&�����ƿ�^�#1��S�V �ᭃ�ks/I!kR8h�>P&�,(�1Rh}T����(э>�P���㏅�4!������V�(��=|�s#��Ae�h�H��*�7��h�{Ñ��fl*��Ǎg�׸<Oo���;)O�C�<\�G�q��ʣH,x߹*I�H_e��B�U�)��w�� |�gO���gO�:��i�k���Q0 4��B]�t`���^-�4t���0��f�0�_�~�u���/���R�=���^_7��T{���rlկU?��,�z�@K�Գy��):�H`#��L�s�	{x,E;X���}��{䭼h�3LEW@Xo��_����4���Z�6ƀ��T��@ktJ�#����a�R�6��b�[����2�0��s��n��fT1+ȳ��S։k-���_�k��^�7�N�Q�Eu�����M{b����S049��g�4��4���l�	�j�7nX1o��}Fh�hh�4N���~�%R�.F�����{j��A)FǷ�C�9(�=��|t�u/#����.dg���)yѬK�GP*9�m�Q� �kѦ�i9�Q����7��س�-�l��D��� �bAO��qk?���~��G��o�����j|3P[��+G����V�_����k���dKe3F/���=��-6j�(�4r�/�ZFe@���T��1I�4`���]\؋o^��w��ol�wd���8�hD���ty�<zT�"�l�o�n��~��S2�ɮۄ�/�% �*g���U�7�we���8��]���2�
�lяgT?����������u�>'W}��3�K��@YzN@7@�#7�?|d����t� �!Btk�?�����۷�������d��u#��$�U�A�V���<TЏZE06�N��]/�5������h8F޹|~��"��.��?T���"�FY$��p/�?]���}x�6��>����8[+I�3C���i����,¤�|x(*��	UR�@pgŠ����^BL��պ�*�-Q���o�^O�xZ����e��Kڰ(����l�ϗQ��Q�:8fծB���e�w_ب������w��
�C��I��D�y�CR ��d����Y�{zd���Ջ�l(����Q��H~��[;+~2:=�v��k��I���e� Ɩ5��!8܋߱d��� 1�Dm�2Y�'�3��\���R�!�E�`a���� �G?k��ym�,m�$����=z���23� �ԧf҇���K�b���<{��lAӘ�ݗ��3(<kbD���c q���x�3���YF{����:[� 7���<�1yRK_��-Z�Lg4�Rd~1��Q�\��* �DOP`�NvO6֛g����j	�Y3�'�of|�ZH � a�h�B����.u���@2#A�.���P?�4�����}8��GP��߳��'|\(��(.�R˸������R��;fPc�M1?������������O�@<�A1g]@(;���=�@�A�܆j����wr���̬��.E��W%{���� CS�����tL�	�^�`�*�N��6z6`2�;�;M(e�pO�2j�c��&��)�m[�v��#ݣ�[Iݫ�S�@�M��!y��V�o����Ҟ�۳�3{r
�R�RJ��po��-�	W�\$;B�,����lS�+PE�Ӹ*�}\�c˞,�@��QƁ�Nʲ�vDp�����'i��Q>CW���H�P< ���F;(�oN�(�$�4Z ��V\�46^�,g<u��4K� +
�*�*�c�0DB���/�_���ɡ-����۳� �%
��@�=�6����/#j�'��:��?PC��k[��
-G[�Pk��E��e������L� @~��Ɗ!��.�2�Zk��YM1���j��h�V�:)Z��oD�7C[)4 l�_�ܹ� 杸bvu�	���f�2)�J��������(�n�����H��~���\�0] d/�T��9��Q��:�ܳ
��je�KI}�ާ�w.�$
����_��.��;��X�k��>��Q����lp����r_rg�.��
�.=���0}�lqf-�^������2ZWO��A��]~�{f����Z6"�Z�7�}x�����/��'ggR�G��px��#2ۆ��j&AR'P�O����]U�
g*��G�[��L�����{�}�ꢌj�>���a@
x�s͖����HA�u��������������ٟl��ت�jCb�M
�~�g�|R����/&2���拎�8Q�gB�{�0����G�vQ �}gc;���b?6�d�	�.��:|�L���l^Y*��EYH''��M(����$a��6{�N���<k���c������	�ݪ�����C�*��T���Go�|��~����_�7��ا�;[o��vdcY��bgo�q��%����m?��. \rx�2v �}R��	^�."��H���U�J���`�=y��ƒM^w��(2Y�r�ޜ��k��}��v]��Ns�;T�j٭�ǘ��T��\�bgl��@�l�^���:l��$6���d� �pQ;x���Gv~^��n�
��^�/�i�Z�r� jg�gŖ��#e_����R�I'�����u�F���"���hw����A��nC�H��~�Ζ{j���!�������#�C���l���FH�/��ŷ ��ߣ�q�c��4��m�\�F���P��dĖ�<��Szd��{�Z���Y9ǋyX+P�}C����kY �_�7A�5yV�*�&X��U�a�xŞ��b�c����Qm� ]��CG �\ � y@�$���g�|�n��3,���HQ�5���� W��������b�qG�#�A=��ݗ��=�^'�U�mP�i������`(�)`�C�&M�+��a4�Zta�	邋��^+�9�Y��7�S��]زD����� �t!%H�P
�K��7/���Ӷ%�?�*�)�Є��ф;;:��[٩�9N�IQ���i��%W̜;쮦�Q �|��7��ݹSǛ�!Y,D.����FO����	�r5�^͆E۟��z�x������P>�"gg'��s�B	 �����������C4�Y:k
�?����7yt�N���O
���5�U��LL$O���*��9������g��,L���)���8<��4:�[�ʆ+����9G\���)�Iէ�ye!D�LS6�W�cH:|���o�m�)ÊHS�\������y��=@��F�ۙE���(��Wr�a�d!��k����^a�q�A�y�|$�bT4�Dz�s O���ne{���7|]�B���R�k�Ғ��3�tP�3��4 �r�  �]P����A##mf]B6��:i	�G8�8P�F$oi��
�m�x�;�ʙ]����x[X,�i�Ǿʳ=��ٔͳ��5�g����-2�UD�� ^��� /�q�k�h�����n���a��NC���ŋ�ݷ�����|> ��2��a��{ō�u{O�h��4Mu�s�*���?��~4r��Ơ�+�(��$j����G�4�G<@P�A,��8??��ھ}��}��wv������G�m��h�t�7��j�,��!��cY�l��G��ܦy�Қ�X��$ŉ�AaFe%Y:�^]~�/W_l�2U�k]����R��G��O˽>{��]\<��rf�Q�^o��vv���$��"����,P��g��@,�A��b�����)!��_(�~���y�R����7�:�Ἱ�b�߿-��%�DP���ڑS�ۺ�T{�}�R(���S՚2���HJN�m��=j�{�5� �B>|m?������?؏?�*g�'�����ub�n�}��}D�6��3ڧ��P��g)�Q��|�6��dK���� !U�>YQ��nG�k%��� ;�T:v��͠�����\[�&�/��R(�m��WPo�vVS��|���g�i�?�	�@y{(��̠�^��3j$^\<)�����->����==	���E(D��x�J9u&�#V�(������l
���.�칽�!���;知 r������@3�1�j��Qu�u(�8Q�BvA{`������h}�I��:c�rjw���yVF�a�c��a{��,Z���A=2�^������ �h/;µ�Ju8���V�l[��A������W�ѧe�$C�~����R�{���i[����ȿ��,J1�%k��(6�� �Nf5ٴ�	�mVǄ��L�X�S�R~��ɏ�Đ�E��a����C��������J �Sm��65�� >��D��[C��a&�x���Y̉p,�.̄yr��N5YsGĿ��d-�K��S�_�0�]PΪ��e^������ʢ*���9Ⱥ[�1S���H�i�g����0�I���,��\]^���}E>�oO�<q�/��ۛ�}Yh��K��"��<�.9|
� �Mj:���?T�o��q[p�%�`n���8E�q$�1L�#���̹��kF*�����/N'8�PBm���A1���~Ǿ, �w�Y覭�l�$�s�{��w,���`�#��)?[� �q�	ZF���w΁�37�d�	��4>-�Hzì���㙙ȯ����/�J��*��|,��|��''Vف8�[f �^��%�b��	��]o�n���Cd"���ѧ�9�k����	�������E!���΄�/&ﵒz�7�2:����4PJ�B��^BF){�hf��n��=Tu{���wx��Q*��Y���"������!�� RV�����j���kN�W'o\��PڒQ���T�yis����y-��r;F��-"Ţa@��O�>�Z�y���E���@R�hc:�Z� YS�a�{�~�y��F0��X��Y���rH� �]`�ŗL����- ��/o��?����=�����h!ۜ&�W����um������s�DGI�����9�8�#r�M� �'���
��re����|I��\��9^��AIi6\���b�g����o^~[��Y���{��^DG�o���������|��֚z���`������8߷vw}e�����bs^�cγ�c(�U�_�,X�v^�:����}�f�s�@O�4Vw�{i�g��Z[/���涊��b?��F��
�����=�~�����������~��}Xwv���c� ��N`	���KT���6YB
\uކ��ƙ��i��JM�YD����1w���8-���]��Mݧ0�R#՞�az�}�a�	!�r�u��+�r�?v�>}V �{um�C�y���sz�f�O�����#���N��������;�u4���\xeGg_fG�R/3I�C�q'�bd�s�lsߓ�4fe�K��^�w�!�"�n3Jq-5A�_�͛k��A�� �}��oR�Fo�n�	8WHm���5P��)�:����9�d`V������b-� 0������z-x_X����*X��p����4%��F�T1;�b���� k��$3� ���'h�#�������ۖ�!7�YM���wam��ӄ�[���Tk��y�=?V��(7�x�r#�LV��c(f���h�T)�\�� hV�bj��:�nk���f>�|�O�\�����󨟘8us����k�����IeC�v[�2Ыby����]8��7�ɜ]�;�������Xp�#��N�e#�P��Z�(���f�@V���1���l9�#߫w�f �e'�&���n�X���5��jp���Z�h��u��f��h����o>�W�O�D�_B���z����!���P<���gei�\�(�O��3:F- �J�u��[��Rnf�ʸ���6�@E��X�8�o=32Ff���R�̞!J6-(8(HO�6��M�qlaE3��<7�����Jʟ'�i� �Pʿ��j�nȲ���]��C��f�@�F��Le&�Ff����͏smr9�T�q��b���n��m���'?��1�3�JCh<J�	n*TK}���uy
\�b�7k�"� +���<�R,��.��ll�xX���R�f��k"��O�-�5��w��`�Sf*n[��՟����qjn"hR�\�O��+��&�8#?�4ٮ��eQ�5Eۂ����6����:"�>V��(Y-y�X��1M�}��_����J��EI�OI7�w��v�G/�D_ldo�?������h�|�������
�t!��GQ�QFd�������*�f��ˎ�q���L��
4��F�G�����#���IC�f��^�H�޼���Fx;��B��qt{���>�>(%d�O����^~�{��%U�J��^��T'�Ҵ�x��l#$�;���z>=��ی���ջ���Iq���k�.Dx�7^�0e5��-$�m�2���k?+v��d,�,N�!E~@1�@blc�>��� 4���6Ω?M�ę[\ܢ	[���<���n�ݻW���/����������+�aݰ�۶o��4�����]8&PYR1�8ݖ���A������B:s�3��ZJUq��>�����_�z�o�!�ɦ����6{q]N�(��Yؕ���̓mP[�J�l��|����oL�gu�;�n�Г+�Z��u�v�{�<yʨ:�7���k8�+����8V@%���}+q�V�g�s�:�~���#���ur�;��b�p�Z�feҽH=�έg(T�p�ނM�#&!���,Lv����\;vtT5�!pr���Gl�=�[߳i-j�@ido/��К��ᒨ�۠Ə&�U=�\�k�v	���asg�q������-�fwY��j�5H��"[v�z/�;����Z��:�J�Mm��.ZQSY��F�#@�{�*�=��6�i;?s���ؔlh* S=�=<-�ypb���uMs�3:�JcQ���ls�p�gv��-J�"�}y#\�R���1�x��b97�=|"87ѓ��9i2�2�ϥ�VI�����4��FO^�B���y�mrS� j%��T;H�9��f�<�l�GU�PNQ`/p&��:- Q�Ѹc�&���� ��8\���P��Kvy����R��EF�h�<�د=..�>��_����W_9���4��6X�h.�F?�x�d�RЊ4:�rIψ�G���Ԏ���عս#3�1{(�j��?,����EcW��cn��spJ�x�*lW���lV�.EN�b���V٪{���]�n8��٫V.���z��Q��;n��F���6��k�c�=�΋�uvA?9Mʾ�B��Ǟ���C�LE�P+�F��XDfA�Uu��$WC2<yV���7�I�چ˟�4�Iƕ sT3�����tD�v-	��g��N?��H͡�Ө����V6����Wd������^�%���P>�P�[�
M*ڨ��&�ا�T�}�LgtKg��#c���S7I��dw||�y�AR� ��؍��<\�Z,�?��|��
Խ�݁����*��<�F1j�1x�U�=6e�F��ym�O�U4"t)M?�:���Y������6� ��������H$��A+S,!�����y��g{z��N���6P
`�W�X7Sp��@���'�A�O�bo5+o�h8���Q �Ӣ����eA�����w���O���[^��r��7���9�Pr_vX������o�����ٳo����%�Oza�j�y���*d����/=�����q<HN��O.s`�����Ϯ�
P��B���3
~r�3�����A���o�|�(#�IA�r蟜n��肵ip\�^��ш;�f�h���Sq��u�1�R��v������<���P��������ؿ���`}�˫��5qc^r�07R�-gh�Y��V��_.����8v8K�m`�ˠf�
L��"L�1�oD��0�xK�#8�����:�3�V�?�����uh:�` ,Z����J�=�F|f�^�:��8@	�\��с�x�ܾ��=yza�{���0���?茲���Z�ܿy��ӧ�T�E�R�s-�LB����,Đ����pD��[�@�
 g|��q �|ouĚ"��n�4@�h��L[�\��	���n��;��v�L� !j�F�;	eJ�g?/�B�$� ���@��R������݇�������7<��L��MP������?��<B ~ ���#H��B��YS|d� W4��z���� ��;P��e>�w�<c�r�+6�����>g4F�=�{�7&��!�^z�$��QB��k}LWg����?TJb�A����2�J/@�ϳo^K��%�C� 6o��*`�jp �ɡb�3	����\H�a&FC��2�+pw5�e9�/^���<��9���PP��k�+������3e_��X���>�0�c�a�T�9�䈯{$�;{�௒�J�;�7n�dx� �-��4^�"�e��r���r"���e퍵E+u|n�h0NeB��g�^�@,n�E�v�6�9�2Zy��J��G�����<~M�-�T�*(v���P�Uax`�Cs�ٗ�-P5G�C�L� s
!E/��x���NOY8�Y���H���,�D\
ih#z�F��o}q��z���a��i�W�Q�,8�Z���-G �-aT}�EW�P~(���gG�Co�="�� #eNQ�����I�Bi0��;�	IhR��m6G��=����6�pC�(�������ĔF!��O*~U�L�a�Z��&���]��֛E�(`���7��s�����+d��m����4}��.��9�����87�f��cW��E9 �xb�E"r�ό�%�ɉ�VA�lX�y���Ճ���:��.�:��юզ����-'8HӷN�͡~Zi��^O�*��P�m]?�Y��˫+6�<<:�-B�x_� ̒�zf�<�.�E����)0���:ɽ�{rꃚ=�^ x՗=�����(�����e���w:�X-)����rug?���؈�����9(t����ȑL]S&AǓ+BUpY1j�%�"J�}�[W��,�� ���� �S��A�ݚj���ho^��8�?�������=�����]�Kp��8��^G�{���<�T���:�F�f�E�7��H�qЧ��9x��4���Ζ��V9��+�Y-�K
�::~b��g�^����p^���0��6TR����@��'!`�~p��{;+?G�t��{E��B&�8F�ѢY)G�q59��8͑� :/ь]T��{������������?�'��uq|�r}��Vl�-)W�c��g�?'��e���p�@�c�e/��|b�;��J��}�����&����Wi��e��iKEǑ��%؁��s;�H���V�T5�}9���pJ�p�+Ky߅��j�쐪w'T���o���}���vq~��+΄g��7�*& )l����'v\ V�?�܃���g�aA0[������O)�t�g�̉m� у�9�sS�4��˕�@�zݝi����8��{���H�#��H_N���'`]gʏ�Ǔ����h�gƮ��n�����@�v� ���nm//��\�~��2.{���<�!���|ֆ���
i�d�X�~[�O�\����h���Z)k9u��!��Z)i`0o��6�۰���3*g�강�Av|t�^�Nv+K lo��]����ŏ�_�Tv��i��Ɍg����%	�%����q��F�y'��H��zL������@ ꛏ�����p���q�o�-R@k_��0i�ɕ��Y>)U��+�5x��M�8W�߹�A1��1ƚ�G�<{��}~����(S�bW��o�};:Q��5�r�E.����Drw\Тs��若�U�b�u5.8��s���E�,F��4)�!j��":�>����i�M���p�7���|L�Y
GؿFS��'m=M=�����k-�HAm&:z�q�Ɵ����0m��wA{�(��{�N8*���p�6;�25ۈϼbi���"�cl6�w8��#�B�ϬR�`��;�u��r�&���͆Y�q[^W@W�{ftɉ�*C5-0DH-�Cmy�y5s�0��0ʱ̤bk]0k7�� )�;�4\�����׸�H㙬E�H),���>�P����H��RX�����7	�ǘ2ۋf�Y]٥:����6lnl��6�P���� +S��uY��t��F�X�ѯ"�-)=3ŉ��4d�!L� )|��w�:� e���lj�Z��y�*43}��ɹ&/���d��Y6z�/�3՛l������ ��a�b�=Hn�54��1�� �f[�D�)�'r�O�>+��;(�����,E�ōOR}q{#�vs�����L@S�����ÆEml��̻���6r�K�9VtD�^6�5$^S�!y��o>�C�}��������3hV��LC��*��%�m�w�k�0*��+��J�Ͱ�>�{(���z��޽��~����׿�����E8P|��7��SمU��'�v~񼀲',��el)UŤ�Up��}|��������C���c�s�C���T_�X�aX���g�w�����HP��5�r�:�ץzeϾ������=���>�K{{���\p��,u:]7����Ϙ4W���صZ�8_ ���ӥ�y��~����ǟ�~���?�}t_�jf����17�}>�u�d�W �����a�e۹2���̨�-_삄(��;�6��̐E� Y���N����G �WML�~��m��RM�ӓ�᝗�ӳ{R�����T�>+ ��Bz���Ӹ�
B�V"W)�̇��z���?�\���#|���+�7D5�>`�{�e��랳�_0��)��NڶR�0h�)�����׉�H~����ħ��������"�S�Yr0��xQq�6 ��/7��/�����I�m]|����aC��l`� ���Yʆ�U�(���!��<Q��5).��!���r�O����b��@�fV(M߫�<�����x�M�PA� ���b^�Z��3a��TV\�a�s�"L��DX�51/�Pm_��S�!�E�1?��ኴB=�&{��?�K��G����1�鹝���"`����K�\T�h�1#5�^Wگ'2s>w� ��h�<�G�W�~m߳�ǯ����"U�3�2���ģ�,JԼ��su�jݔ#Su`�: �&�B���[��*����gԷ�̨����p���L�YM �۝g����5E��ʯA����`HS49��>��yf0(M�W�e��j��	�ՕUu9S���Ǵ���N�Q��Z�X�B��L�Q���������],����yF��w�X�׈%��;.���ž2�~�2���D�1��d���l Le���{v��
o�a�,xآ��ݶ*��,��e�	b�u*`F�fl���PS�Ց��F/���؋󝼁7�ư�ik�����D�@-����pȷ�Ln��8�~%���'VF40"8�	U��1V�@+�}&7��6�T�"�;d�����Wř"�Bam_�u��8#��AԘ%:/u}����N�! ��Q��t��|��eߟ���;Ags����~�Cc�s�yF7�P��<�~'��82@�=���Ɏ8=��a�=h�9<���"�
��������MY_ʓj���E�*~�J;�c��G���L�s��〞�d����6�B�@�.�����%����XעL��,6%��WH�\���`��vrp���o�۳�OHQb�)f�4�����+�rq�*і��Ziͥx���&��QL.�`O�n3<0{w�,��`�{��_�~����6d'{
��߄b�ԥ:�I@������?6	]�N����8��&���Q�]���)����鰯t�dU9ϼ�)��`���Ξ�����O���Y�fe�7p_ýB;d�������*3�%NR$վ��{�Gv�9���c*�l�n��@j;������um&S�������Njgpb��v��K���/o�ܽ�ׯ������>�xC=5����iOG'z�,r���?��eAܱw"�q�,��7ʆ��Qk�=�Deт�ڭ׃�pףb}�4k�����´5�jf���1ih��A���QU��J �2���/�O��=,��O�(���/YWEb���'�UȰ�Ai�r��q�,$��%e>WS�f�n�%Q����+��;���ٲ�t0R�ވ����ΠP�@�fB|,g��F`3z͜�ɳ߫ڱ�j{�x3���f��P>{��<�U�/�������1�9�8���`nG��H �5��5���$;WmI���M��T|aw���]�ud��*clc_`t�DI~�������$�u�z���p�9���O�F��l*g�����P�M�P;��5QW�:�����G_s���5�q���L�K-ٓ�I <��!+Č�d�A�3^�'�P���,���S�ɡ�=�≁*�����;��m��yf���ĭ���*�E�����^DLn��_�"��h	d-���� ��Pka����߹�fT#���K��y��N4::�m[3@�P�����d�o"�c�m�N����/G�um��?���u������B�� h�G���jYq�9���=�*�Z�&�=�	�
:1��참��r�J�Qŵ�����k���h�S�7%R��'O���Ϧ8o*�[��-�0�_�����v ��E�;8x��� 6�8�ᱫL%��"�թ$Q�'*I9X�"[nJ`��a�4��_� �]½��΢J�8�c�G���<F70�	��I>�Ѡ6ꦘ�tǚ�-���i����P��Y'tyw���E��\)��'��ِ���Î� U���nK�,8C�P�aO�\��=�JFm���BL#ϝS�s�SM���qGd
��,V -��jъTh�(�K�I%j��)#A�Y&��9��,9 ��g�ٽ��.�� KR��K�&���9�Ƴ���SDu�%�*E`f�oEz�X���Lt�Q4�e�Q[�5�@�
-	��Fs��pp�.�0@h�ۇ5)^l�q��8l꒠�6�hт6�ý�ݖzPI�dz����}k|����e�������T��j�7��f��o(�rx���bSx�X�(a��YJy�=���yx�h�))�p45 ��,πTg������4�z�ǹP1s���2(۰`�j�����N��~S�:��@�|C�1���A]��T�|�%vU@���5A���s	ʆ���s|e3�����S�`�-� ���Zn�!@F�wo?T}|_�_���e�a�٢�Y8���o���tSY��Z!Fi	�:��[���5��Nٳ��=�.�b����f�ևl�r�v��ӨT����(X#?G�!;��O��4������q1���j�y�;��-����˿������_���gvv|jG�9�X����i�)` 
3k�������5p<�P�s@��aK�iO^�9_�\�k9`c���W���l��hN<����M���R��.��J�yP~Lu<8�$J�A�l5�� j��,�p
��2�4`K)�R������r/O/���tL��%����ؗ
�����߉��I���	�6�Ԥ���8��X�$E�ӊmn � @� �Jo����k��)�^�Ǡ\�����%�cH�o�,A�Ze1��QC���gw
�o�?�T�i�P�bL,ȳs��fY�G��>�TT�,{ے��A�Bf�O!��,�}��u�:����`���b�(QR�`��.���k��v>J�~�rO�4�����&�Ī���ۚ�x�*Ț��X����	�6�qg~�I����Z��y���(w��G�ٍ$���N�"7����G�(^�j�'>�8@_<a��{{V�ItmU7�+�ő7�@���Y�M��������W�{��e�r5��N��`�D��9�6շ�oL��\��yt�Ύ�Yz�f�|& ah:���%�1����/SG�V�0	8�v�T�~Ÿ�3���� ᣎF���д��g�:+q�� ��R)OP��T���V��K.A�0X��p���*/��Q�''���
T���f����'���04<nz?��f��"�U#@F�#+c�@>Ei��C�kŧ&$tE/�� �=n�g/,�Υp%��u]Q>����|%����mևFz�e.��m��V����5{�")]�D�� 壝�(������j�0]�����y^3����Ʀg�4�S�m̳Ϫ��p���-%�ю��E�vtH�ǜ����� q��L�I�^��Uv��̃0��k
�4B�N��p��2��8��-�������6���Ͽ����:�{���Ğ��z�� 
��0��:�=N_�lyԐ�/����hf�p�����&�[_*��/�Q��޽�Ѯ�|��D���#4B_��N�z���ꢰ���Dߙ���N���j&��I��!�S���i���z|t��3��x���<����Xk&;��"8�h�
[z�^IG\gh�=xsz�=��м޺�c��7%�c$x��8fF[�������iI><,`� -d����ʳ��={iU[��P��z9�]]})���]޽�X��'���l���[A�t���w0w��
�nT#v4�D��n9�O�/`��� ��[�xϴ&M���:.�oT��3�M���	���F�~x��"��0r(�|�����"KȬ�܁��9��Θ�������_���jO���>d����a���Ng9 ֧O����L|b]"|��͈7N�.{xkg �tؑ�</{d��,��u[ j�;�9|��-w��k+����2W@3�b-A�bf����Z�2����?��i���H晬�2 �{���8f����s�Job&2|`S���7b�:,�ϙV��5fQ��y�F"l ʴ��a�t �j� �Ã2�`[��_��G,�+�lPɷIdX�q?��g�[�a_3���P�T833]D�������|�v�~������2�f^��k�Z����/�6|�<L�5���Q'�惺k�k���dej��`C��P4?�i����B�,սl�it7�]X[g�������v6J�`����������$s�U�4�ޙͯګs��x&J�w���S-/֋�,558�''gvtxB:��z�Ft�(�׶�t�;pACG!�N ";��n�{����C����)4��)�/ X��죧�)j��u���
QV�n��uy��P�*5#�@�T+�$Y[d^Ɩ�9�;}K~��1� �0�j�m���f.m��M���E�������:[oS�(�?#�����f��4�i\���bT��Mq`���s�}��~N�JJ)�a��˞�2w^�Q���&�I�*th���)�~��@ϽÅ�;$
j #�d�Iz��=��qG�wXct�x�9
�q�k���c�n�1ͨ�6�To$�M�X4�ふ-�8mq$�ŸGr5�r/QH`;x��8�m��y@�el�X�F��o�Q3D�
�)�.��@�k��}�#i�I��Y|g�<��$ygsQ����yW�몼�e��5�},�Δ�(�����#3�N�@d<�k�����|���"(���>u.+c �CH�')!+P��rkAM`sb����%�A�d�W�}FʃM�mr�������{�P$���h��E��]#j)֍2�[�N#r:�t���)B�@H�+/R���؇RDE���u�M�Y$�ث��N e��s�UC2���4D���M��<�pP0���p_W��"1P0r��Xd:�J8��]Yð��sgc(Ԧ�x{��|�ܶ#Z <)o��쉥-�!*�gjv�1�z%+?��M�i�ç�L�&�$�6��k���`W�?������W��û���tV���u<SD����W�����{������vx|dmqp��kWIHS hP���i!G+@~�lo����<�C��qFUK�c��z鷲�؛m�g�~�h6@�����L6.�+�w�����)�ݙ@�AЙ+���{)��<����N����~�R��g�у�c�,�i�QC��gP
F-
8�6m���<�u���WP��. �mq�/�㾶����e���=����swU�DG���)�z�F�b�+ KH��r衈���[9oQ9:������1.��50|��
����΄L����6z\C-6��zq�bV#h��=3��W�K��?}�G����_��_�/�}4��l� ��~|Y�^�Čӫ_~����_�B�y��s��i�e^���X�/'|O���e��ľ����-������_��>��/�mݣ��������X�>_�'k(�Ul�e��x���{ C���8�
d��wY�m��}Y��wf�oD�\0]�k��jc���5�c�L��澜�T	\�ն��E�r��?��{*���������ɳZ)���/�v�J`�����>9�?~��}��;9�gF���Ž�D���1��?�����W�P矇��/e�������|s�&�8,���?{N�VWE� z�%0~����y�Ɔ�7�u�)�`o�g�H�t��H�8����5�
�U�9yi�����l��TDn(�#Ptq�&p�J�o���z�%o&?l&( C�� �r�/�m��2�+x��b=�c~[�9��]"]���`}]1�\�\۪�R����p0e�,��&l�Tc�*CA���Ju�l�����,�I= 4�9yQ*_�
��������j�q�@��T�6k\:�u�Ɩ���!���999��ϟ�_����_�b/�yIP��.����G%�=����4�0���|�y��f�Y����-�T��0 �ׁ�G��f8�)���/�Lq��C:?�g�u5�R�q������şe��@���A���u1 ����O$Yxw`���+�wV9*	j�-�U1$�\ۺ
��!D��Z�<j�j�EˢLd�vu-��t!�ov��'PW����Ŧ��  c��AdH���C�;PcDE������#��#�/W���jc�ē��\�qǆa�*�ߌ�S��2��LX5�\0`�eM���/��3�8�kb�N�jP�,Y�9(����i<"7��"��+˙�����$���[��\/�8 � ����,{�T��;i��{�l�Hn��#��Q���p��Vi��@�+E�B�^�er�m]J6E�#��˲�g/V��ֵ��i��h�v�h"B�&�h`�U�-L.��ȱ#@��WF=�jyf�T^诋ڜINI� et�.��E���+����q�Ü�\Ch@��4��{������]g������`A=�v��y�N��̺L�<F/�����m��ތ�����i�,�q$h�Y����.��p�����+#��Cr@� ؍~g�y���j���I`F8ْ]���2�p�CMM�*�O%8�T����v[����O�/��Ц��oُ�EH�gr�Q�7�R"U����'�&�fV�	b��A��y1��dfC�s���e���{Eb�A���lq-fRN�H�X����Ѥ��V�0�m(PR�������P�:��^�wd"�k%�����{-�FJ�ӮnKP��#���1�����޾�T��{{��ܻh>>���y]�k��z	���8t��8%��Lte�x�

�B�9w���jy2 �U�w�uQ�q{7���R��;1)j�3ұ����Ei��	�r=D�=��`�q�W��RZF�z������W���c�۾�ց����v��RػL? �Jp��������}���g����,���|����7o4H���+�XKW%����u	���������c���?�z�>�^�	j�D�~��SU��^_�=�����]�g��Ӥv"����r�=����eѪѿ�:;�_lC)�i\�W���/6�\�JR�f���3�!@wVl�l�˚�@f~�9���{�:���H�����k��_�����������r�.������H�����ÇO��:��/��}kߖ$��b�Y[L� z�t{g?�}g?�Xl^�;�k_�$�/��7�|���:O�3�紐7������?������'��M�4�B�$�}m+FG"Lj���_�<2�Isu������-ڒ������Ka/#���x�á�F��49 ��o��شsE��m�{�T�4t����b{p�A{��-i)T�ԱQ��ʰ�v|y^��% ��"I�}>aq�ې��KX�laZ�v��-�T/`k����b�VN%�d�
ڏV�̧J��S<�qJz��K���+���#_�J�_|���������_�_��w���"l0��E��6��M��AG�B�Hfe#����r��p�p�^�����?�9����ǫ*��J5�lK~36�z� hpx(�]Y�w%�z�duR�3(ں,o���/ɔ��-���f����L5�a�|>D���:�#ɂ������b��i(�4J�'�sW����]H%J�M�|ù���,��(F��ࡥ�oKQ*[�� �}���l�����ɦz!&&W�0(�5�e�l1�t������lt��[`Y�ާ$'��'h��D�7�"��}VhOB�"ј"��K�Rxc���#�T��T��T�������)n��+���>��@z�:A��.k�Qm̚�1N���P'UN�c�&���Ƨ�!kMN�VlO� I0B�0�9Y�g�Jr͡�/��r�<oq�ϩ�tYlӹ�!���;!�*~����,���4���Jn���(�A��=�f5%84��ա���*�Qoz%Ul8/��������ݝ=�o�����7o^Q:���Y�oM�4�ٳ��x>��G�Ul����={�v�3��g�"8����G;��:�J0���x���9�*��hsK�<�_2��J�WM�"c�|�ƩtP�dc�t¡��x�����5Z\�S���C!�x]�_T@��tp��xo??�H�Q�s����FT%�W)OVXi.w��YQ�dW|��:+��]R?���rl��|��;��T��a{���������چ�\sЌ�h��u8ND�Մ����X�4�9�u# �dP{�{��$��������؂���=8�֫]�@0R��\W={Vz&ZMV���x6ח��$�>�*z1꼾��9hQo C#q?���{���z�#���J���G�0x�J���nP�92��n��ܿ{��>~�H���{ݝ�Za�Ƹ��)p���o�|,����v�1��K<�;;C2T�/^ٳ��v����vT�#=4��֒�bh^Z/N���u�S��[XY�!�Cߪ�ۑ`;ŗƣ��$���w��q�8�m��*��P���>���W/�7�YiZ�6���wϟ]��gWv}ya��������A��OY{�:��U9���6�}�勒\������U��]����)Ƒ����$Z_;�H:�q,���/���,�5N�P��L���>}�a�XCW%�yU��/���./.w�����]�8/I�{��Y>���w��?����'uqX�`��я֦�WK����;��N!�lF��۴�C0��D�)�}�($�.�k�y�8޷o��7��yسH�[KD+�N�b����R���s ��{��@��Ɏ�ۮRk�֘��b����4�3,��`��6
"�o�������}�f�}��.�W�����S���|�������Sy���H��4�"��$KA������9���,�����7����b���/�ׯ��}1g���ǽ���(�I_��d�}ˀo�7��-Yܜ�w�]��}�ga�;�%�Y��MM|g,"Ӭ�L��*�"�fd�P�@�{���=ޕ �|%eT�:"m�kh��E��
��Sr������5�g��S�Z�w3H�����bMҥ�	 ϵe|J��BAɡt�l��J�qNךO�����B��s��F�@G��|�r�ðRo�䌃3s��5�|r/S���U�{��c����!):<�A=Y֌$�i����g�y:_�u�{4Ҋ�vZ�b�ŔlL� �5<ȱ�NX��fx*�-i��A��dsY��ɑd�5Fw�
�OU�b��bo|�W�u>ߍ��5�A��4,����R}/�������CT�8́-k
켴/f��ǧ�i:�eqXd�]ƹ�z�y�}�]Ea�T�1N�i>�H���:�=�A?�~�%`�H;�-$��:��{��XPC�u��cB����w��!邤��W/��Kя�.�Tv��'�A�i3)�SS�5Ռ��%y�Ǉ�Tݕ��m�Iw�yϾ�4jt ���V�K���8��4W�؋PC�K�U�aw���JфQsΚ�������s��׸/=0��ќ����Y;4fKJ `�c�T�dr@�\�i�7��]/;��_x������\<+B��pYw=z�=�*��k��ɲ#�J�E�)+�U��Ц:���D_ktV�����GOZ�7\�Wk��-����6��Ȓ�F���@{�@������A:�Up{X�[bS�С'�I�Z����6��k�x+�Q˄2ư�u���&Ő��I l�3�Aa��z����ުL�z�!�w�wD�on>����E���#}<�p*gb' �.o�+	��@vW���KVw��v�
<@"P� R_]�����Tyn�������c&�<QP#C§�m�,#������IJ���d�R�L��+))���b$LĀ�����J��$�_}�I�*G���/�__R.�͛�%Ayn7��m���`�1{<!�y}	�3���S_b϶��g��/�����}��m�D����ˋ�6�UI����kG=V���ϻ�|�D���E�����$`���o���Q��rm�7�א))<R�<���y~a�O��m��
�7�e��㶘̂F�f׫K�'�W��FL��:/m�����Q����m;�5�84ۤ(b�Ҋ��Ǐ�X5������VG�X��(rM��9J���� �"]�q�B]�w�ӬT=�<���K?�C�������#�7�sh��U���L���桮��
D�r��*,,)���ԓg�͒��#XL6�!4L+)����t����п��_�����d_�1�����x��}R+6���4������)��c,��j`���O� �����\t�����E
�k`Y���kN�*͟�OQ#�~Du&�K�����D�v;p�rm��d!��m�H����eeu?��D H����+�m�6Tf��V��<S�sZ %��GU<瓳��|E(�/D�B�sE����39�Mg1�[����'JC(�H����朐��_x�R°9��ۙ��^��t�71Q�&�xjR}�=Iф-it6Kz��tU-QNL��Zx�Y=QّB"9���/��+�2���#��+w�`��BNZ��@�Z��i�_�� �"�m�xN��õ.�tnѐ������.�?
Z�`�ڭړΫI���1UE�yV\�̉��7>��f����y�z2|j$Yp��o����a(�ׯ���A�:N�>j�H�#��]F��2­'YN�׊����g�6h�N�=����Ɗ0�J<�@%��._Q� h�kW6xmj{j�h�)u}���?���%�z����7�_���H��Y�Pו��H	D�d��2؛��(�rmQ��>(�BE�?l�O�kr�j}ԀW2�\��nNJU2�٫�LS����s�>`�9Yc3P�Te֟�?������(��"b����_�@ ��m��
{Y�
����>�h���T�ڋD�Bэ��HZA.��5�L�b@b|�~̬�`���T~�{���v(�ck�>>�$�h�]S��Fc�	�0�\K�#�q�s� �*X�h����v�R�&�v̶BE	<D=�VZP�.	����SV�ň �?�gE_����ږ ~`�T���^��#�\����Y��Ľ��.��zH�7��v[���N	m��QF�LP��l=<>h<Nε�3����=-�+@ԡ,�T�D1�&pw�=�*�/����|��[d�Y��'E"�J��;�F_6y5�ڤ'��, ����FI���\��tɪv�E����#�1�d�X�
)��.z���k?�;�!�)��Y��T���l�1�M����uc�^���zUl����"s�*���!A/�����|~��K{��\�؃��R�e�F)��n�9�4���6�]�6�ݞ�k�m��V��)R���m���b�^������5�}�w1�a�S�m8���ʸC���>��E�=��Z�͐��WVa����\��	�
P�N�<*�����G�X�wk�)�r�����>II�wޫ�A�X�>�Z��sa����/����9U��磏s��q?�D?��oh*�{���� \�2���5�����
��2�y	t-����s�C��>.���$�A���e���h�E�5�j&��P'�^���H]K9�1�}H~���H�>�gi�} ���`��AJ���P-�Ct|��hr�����1�ƹ�"s�`>��ԇ�)�I>!=IJD�.�
�.$YؼX Hv(���/͎.�f�~\9����MMx�3}BYO�#Z�Zo@�3���$h�J����bO7�SH0h�m����U0�n`��5�HT�t�CI��[p�18�H�D�UU!^�fE�LЏP-���P:����E��<��_�P�V�{�]͋���9%��	CrNl�7������p��d��ڌ���`Adk>(�3�����b���_~.��e��b��@�iE�-��*8�5�Uh��II�Bռv����r(?�4˾G�h���«�@��xߕLBhr4C�o�ᗷlF&-�)'U�L�"L\K:9rGtN3��3�r��ƚ�ӨX��s�t!ҳ\(��9�uN]Zu�����b�ڗ���e��݇{���(��uI�^�xn��v�H8�2���a_��VL�@B�$*0@��#��B�P���8�!�q��1��C?FseN��Α��L��=lg�����'&%fD��%Y�_
_pʎX�>�5���Ҹ��f�a����UU<�T��TJ�,@v|�^�́}r`�D��>�V}�j�l2�NW�1o�=�tj��>�<�������̞�+V�O9�*����K��L	�9��[�b�,�)��sg�)H�|�>�wo��j{:��G����5 ��T9k{���[y�s%I�f	��:�{�@Q<<�
ź�a���j.?[w>ǭe�	���n�$���S�I�@���J}OA�?���Z�
�'�g�扉��~�k�i��]��������}��r�@�+Yn��f��XE�ZIG_��>� `F��S�ɜ}d�	��7Jtɞɲ!�-e� \	�X�b`�D���B�:��b�6牽V�le"�����-jB�J�rϲ��s�b��4�zT�M�jg��U9tT��0w���"�5(  ��j�!�ױ��7�������j��+,���S���d��+=�$�J#j�T�������3��H��,c`�Ѫj��(=��-��<��Lʑ �G�⌒�˫�
<D�5:%�w5���Ƚ,�}�j����
�b�x��q�+ioT�?�ǦS��̌��K�7V�sL�x���s�Z���m�N(b��|rU�0r���w
X�x�p#�����z�ǅ�t�hJ[-�c�AA)���WvU.>�$4z
z ����R�}/���lL�	�E9s�8��0��h�����k���=��X�~�Ͼ�<8e~A��b���ԡX'�F��͘۩�ß�zuB���fBӱ���D�}���^����㠜.��Cg;:����͝/@cu������Z�gϐ^��CRw�2w	��s#,�m�Q��e��v�`@�ٓ)yo��pJW�2��d.�*���X���}�0��dMD<[�5� U�5�H�t�f�%_�3�1/7'w���/=[�l�i���z�z"ae�A}-Yi�wSe���Rg��d�v&4�O�z*���<�⽈M�C�Q ST�~nAk���L�"���Y�!�3���y˜|� K�Y*\N��`A������E?�^��.�$��>$7�ϘYk�{O_׊c͞ǇGr�� c�g}F�X�N����������S:ۂ�?����3Xq��5�1�a�z&1&tTVJ��|(s��V��xzI5��z�dw��%���w�?���+��Ϯ�)7�^	<Wp�P�$̂�u�Y��d��(�9��3��Ȳ;|%X�A�#N<�ʺƓ�CP�ܹ�+��E��Չ���g!j��-��{z�[Lh�,���� ����A�V{cs�ոOȩ��x�.��P	���4w�4L�͞s�bhy[�ѱܮ}ɒ����ۻ����h�nvv���Cy��%ۖ���!�٫�Q�G����RP���ʮ�f�����ӫoʴXI� �lu3"`�U����@���1&��S��9`��E�DET-�9	�
ɡ����,��8yTQQ�0���j-Zo?���ݶ<wd� G��b��*T�"�V�7Uf(ZquI�ľm��zvZ�����p�*hxҎ�����R����}�޶O�o��#B6�i}-�5�k ~[���I�@�fԟ3V�(9�"�#<��8��"y
5Į�q$\S�����z0�֠>[�9����P�u�1)H^�}\� (sV��Y[���)���y�<A̵���/�������/������ߙ(��=� p�w���=��W%�{f�e����nZn��ٞ =_��|����+WWW��w��{ZI�a�ۻ���������m���ߗc+ɋ!>�t �$HJ�'dɩ�c��dM����|����yr�����6��V�2V��_�?��:<<{P̙�
Q�f0^�4��3���Bܿ�t��ڬ�[�B��?8S$D��_�����[�K&I-x�I�o#�YwCpJr'o9�R{�R5�~��V8�&��>_ W�i4ohH��Y�䡨*P������>TsY���+��/�9X�5P�,�~����'{zP���
�W�7A�o���N/j$��iy�e�#����u���L�8r�C��'@i��Wj�1#t�V�ߍ[��P�Qu η	5�ƃO�ZG�(�L	�+�h`��F�4�U�Pjik#=&U��Wl���᰹):QS��%��9jC��Z�Z�D{UCyWD�h�VJ�hnJ�y��(�	�+�h����//�����P�Lp�G4pA�A]��4xڶۡ�%�z *qdU+�Jd}�;�
��"�r�¸���m����s��i�NE�9-s���ρz��8Eo�S��!�-��H����UP$i�0�@��a�j�g����3{�d���4��O0�F��H�-�S�P�؋$a˚�^���P��I�cA_0��Y���h!���q��vH�v���+�[6�f{��G�1����9Ӹ,G�ݨ���DЁ�\t鳯9���&:P�(v�3dt]�9!�[���go��ԩsu�_�9o^���>9}������>���y_C��LI�����A�*��-� �Z}f6U�T��4г�9+��Dob)0��J��4�=Q�G��"xA�o����3��tN�j_�_�%������(� [x{�?_&^��c��M΍���[�;PUܕ7WB����i�i�@��$�$��+��#f�T���T,��=�@��ng77�om��P�$+�#��N�Ց����=�{Zl�ٯZ1%x�`���o��跈S�Yp$|8�5��ht*�D��p=�B��
��6���.������/��";�1ɴt�M����Ԥ8�!���J�P��q$�G�E!�����ݸ����X� u����'�*�	V<@��]��Jlt~>̓W�(P(�����ފ�LG�X���޽[����[̘�S�I�.��w<C�Cٮ�~I+���#�/Oζ*�	�G���XU����uwJLuL��J#S:��+��P����F&��䊩
Z>�xQ'ˇ�?�-9��<<���=�E��5��V����_ �;�R�����vG%?>�?���?��ٺě�DEk�I�$��a@��|��ۛ{�m�ނ��-]�e9֎�,����@E�ۻ{����ǭ��!|���˲W�{��k���=|�no���7������?��?�$�w��v׫rB+-Y��·��iܺ��R�%�p#ɚ�S��>�Q� (�����qLӸ]#� kP��h�'1���T-�q����h�x.Q}ӚW� �	��1�r�4���ȿ�"BYT���k9��m�X��&��˂B��ndꖨ�\����ճgvqy�����A��0B[�c�M�9b׆"�J��0"R:�_�~���_�5)��&O+%h����w��7���}������gW��7��˒h�kbIv��ټ@%��5�u�\V/��;�!w��������S_;����e)�iF��8.,����!��� 1�f�)� PuASn�e�ת���+�(�O$mT)�B��[+��|@06h�1T��6$���^jQT�����uħJQ����T/���y.u#e��ͅ=�z�����hI�@3X�"!U6�u(���:�}:��į=�k�˨�Ugp���,ɇ�Q�B���N��m=��O,M�=
�͊}�W1�Z�]t"źNf��
Q\��� ��0���:�����MQY$w�T�^�r_���E��<����QF�ؤ�� m��"�P�r�J$Zu��!l�T�=���	U�^A�b"�W�B�_�����
\asb�%��:
�6���{�t���#�	�T6�M�쪊S�+�SՅS��X�ð�� ]��0)�c�'��T)��@#S�y�O�AI���@��e	����Y�ݕ�sa�7o�G�P08�$YϮ6%x\��kE��n$��ʜ�U�����7I ��q��������|�^��,!�f���X9� �CD��0�����z��U���G "ڬ��γMX1B�E�ۚu�P�n�����4L�E �h�sZ��R$�#�Jl,��9���@�iߖ �g@x��+�Uo�e��Ŧ��UyO���=������Gv�h������vk%WY`��e��w ��ze���k@�5&Y��O+���3�d/G8�u��Ril�_��V��XM����&�M���A&W�X�Nր.�����,�l=�>/6i���G&X��F"L��	��&���&D]d�R�>+�������n+��۫�J
l�{�ۧ���w;���M� �t]4��}��x���/�uM���A�J��b>R�+��
VL��	�6�M�{}X%��wicG���*��|��E�PH���� ���̌]����'{�ᓽ�xc7���t�̭��+Qܚ�.����I����h�����S<g�Գ+ Kڬ;(?��`?���=����oH�~���cI꾼}a�g��r���P�+�����������ĳ_~Yb�{�VԾԉ��������?�?��`����)&���6J�{�+DŃ
����+�!ƍ�����3��er ��6���8�$9ɋ�!�;���LiĞ�Z��r$p9���N��)����G��1�hG�5��-cV�\���A�z) e�"�Il3W�'p��������~ޢ�s=E���L��������(�pv�U�����rT���G�lc1u(4*h�~���
^���/8���S6s6d~���n�����%��#�_��[.�c�K�]��j�h�Ŝ�$2Y;͛~&0����S,��B��N�s��w�w?��{_�M:>� ��Bua Q����#�.��uQ�Ҝ�\�sسӪQvIT�p ����n\�K����A�A�����S�
�}OZ_vIqI��N���<b�IE�jUI,����-�캬���8��J�s����s���i���H��f��%�������<Hb��̫<�s5�+�
����J��ɋE�iH���P���h�W����C5�n�iei�~?M���G���:���ߴ��_�ڞ,5���\�s�&ҫ���c
�>w��狅PG�>M};Ic�=���X�Ó���Q���Tq���q)Ho��HaЇ��;w��]?{a�%�����'��k`�'��6�<�{�u��d��Y��b�;�X�H�%0pF��!�Bꝑ�o�A$�m�]��g�!!E�*?�U�͑�[{ڨ�L��׷/_W�*tOg]�%0�q�.ig�$�bn����ޣ�����Z?F���1��2&����F��$4�J1~���1p��[;y��Λŝ���:�l�%h��?��p{_�TT�6?�l�-~��^��P��TY �=-��(��W�@�B�� 0�w���#a��Y�B����!�P�ê���=@D	���
V� ��l� a;2�RҤ$+�G*ub0�N�]�sU-S��0z��4W2�]��B�D
a+Y�5���H`���ֳG�ߟ ���_�k�N�
T�K:�|�T��!�5\P�Ӽ"�IAՄ�U$س��8�b�0���"�����C�{̞����zx�� h��|��0V0[J��c�W��{L�u���}�_�5�����@�G^O�����#���N3¢�"�$T���˅$uɽ�#�ڴl3��&_ۤ%�}a����J���k3is�`o"��� ���h01Xp Գ�7w��ۏ���O�⪵��{�QICRÙn�>���ǒԜ��� �&$�It<�X��Yqm���׿����my�g��9��LRߗ�}_�������P����߽/��'{��3%Y�Σr�
ֻ����{����7o^ٷ���^�|M|d���n��{��},���}Y3�;&�+��2tS+є�ḡْ��j����q]��p����§�%Ks�t��F�W��Պ}o4>֧��Eg9�+O��uJJ�7��c�0y_�>���A	�^�{
)2���*-������z��&�bv��	-*k�]���xѦ�t1niY�\�uY�kf�O(��ް��UD7V����E��ɛ��l4�[=LD0!�
�����ꬼ��]]^��.��a�`���-�H�����_�uy~,��|���_Ѹz�f3�/dGw1|�rzG��f!0��r�����'=���*�����܉z���R����8�&M�;5tͪ$)�D(�i���h1��ԋӤ^T$8
����M�ͦ\����bHR	Q�z������ ���V0X�ZJb#�>_��'HTdbeR�������_O�=���I��\0"��b��3	���ԛu&�[@�ҕuF����R�s���ٮ80��^\��W/^���35�&%ssoU�xE+��$�X��}��������n��+��P���k�4��#�A�^X@��gս(����Y	(פR��@JCM;���^���fN��2�I皽�j����3��=���Ҟ@�(褔D�X�v"��M�Ӹ���c&T�Pm)Ze�p�"�z=���HZkge��=wA��k3�Ř����}(���m����@�1`,ǋ`ώz�5f�A�򿛖_��Ć�}�h��>�����bn�s=F�E5��؏�6]��J�P��2g�I�kO���?�_~i/0+���Z/�3JgO��Ӯ6`���g�q�7��5�JP�5Q��OgYh�D�3KN�����<�E�6���.d��'��e5�s�U��:���e�
R�
LI= &�Ȭ�#�#�m	��&��I'{�<ۛ��Oӎ��5P�h�o�O���~]8�+j�IK{�=ĹE#P̑ 	@���@�e�a�
����Sqp�O�v���j#����m�nۦ촥e��;�-ؽt����4�u&_�r+$���ԦM
���|���k��Gp���=�D	m˪*�fR9�_E����@���n�a�xKd�@�uThͰ�����C���cI��%��m��(l�S���rm���	�ֲB�*w���T.�qz ���56���8U��F���+���� �6�J���z;�?
���o�U[��;/��Y����������ǚD�؏>�8K4�TpM]���L�ő{䘕�I9�qPE��MY�w�Ͽ��r,��������z���C�k���'Q܏S�G�>E�MJn�}|���������I�g�]�Y�Cyi7ڍ]<S�cT1��V��%�9�MM�G�L���A��35o*Qp�(T��,D����Ѥ�fC�3�aC����;�h bX���mGUC�;^�HYGO�5����'{�߾����د������3���v?ڧےh����ͧ[�eגh���,�{�-c@��A ��p��?�Ὕ�[��9*�w%�ٕ��2��y�>�����ݑ�3bVK�I@m+6��� ��'�H����o��h�JC��l��)rq'���xƊ?�Pq13Qe%���Ϛ�F��W��q��D������C˭�p�(ێUjީ�� ������%��}��\�{� "Q̾��ڷ�H̱:?�L���`^�yc�roY�4�9,�h�J��fu��(�4ξ����%�d��ӳ�.U�M�9��0x[��8�r����Pދ��9x��|�x�{�t�&[�hƆ�ųf����ؓ��S�D�	s�j�,\Ļ'H��~�����r���j�\�s���x�V��
�c���b8���Z��Q��_ͧ��5����H��ԁ���\U�N;iN>·�F#�TǙO��X�+Έ�����¥#�U�ȗ��KM�=LҠs�Z��x�J������f��@���jt�F(��Ђ�V�4�nI�Z��U�9�GU������3Pi��zf�̠�U��M�Iz�ʪ6J���-|�클���QwG׹�a��V5"�_\���Sݨ���bqmf)�6�`Ԇ�X�0o��״����u� �8�.Z��5��V�M� �jX|}-�荎qM�vV�n��Rԉ����9�ܧX����,��!����J� 0��� 4*��F �+�<Sb��u��y��vȞ�I����g(a��`P!k�ʮ%G�f�{\��.�<���no�YT���)@�k��}�TɉD��{_3�� !�)ze�\bn5E��X�y=3���e��$���ߡ�e]~�u�����#����Q��4�֮.�Hz�ɚ 7�ހ*��1%M��q�4���BeM:��fZ�K{cF�S9�[N{k��2����C�k$��uZ|�|$�ه��K�O�ѻAX.��>�Og)�\#=����>��}c�p%���^��o'�AA��@l��t������r�w����z �CI���$�k:?ht��M	��G�2u`-W�8Zp������i��d�$��@.�g,�xSC�*\�6��Q�4�p��ٌ3=y��'	��\��I�*����'Η��ʢo#$�}?���HC�[Y��(E��������~�C���ߗ`�g%��Ą0�9f��_���D� Xߓ_f�
�W�Φצ)��%�~� ������Vϋ���6��#]�.ꓒ��LV�EF�C{��$I�K�u��Yr�h����T��]�nv�8Ġ&�2_���8b �������CID��g��H�F�������('+1)�Q��vg�U���jP���P����[��0�����Re��}�ߔX�`1Il@�; g���˖��
p����qxm���$�����jI�o�3�܏����7��}]�/���Y����ا�ظ ����#u�Ŏ�1��SK^�ef��cV��o�9c5ݫq&�+╶i�����q{��,��kz��Yu�G�qD����;��l��I�y�/�ym��	f�Bu=}M9�{�È���,�uSPE��߫��_���
/�03���YM�q�#ъ�R��Q_�f�I*C�ʅ�Ñ�(��M�����7����?ۻ���vG#��y�u5ˀ6y�9;�S�6����j���#K����E ��q��L���:�YZ�j�Cc�xf6s�"������gV�������p���+wrS�a���]\��-���g,�F�&G��l�T2e���&@0��v`@��s~~i��T]�t��A`̃@/��E�)�� �Y��B1�m���}tn��J�x���5�<�j��h�O.��4Lx�FϔU�п�6S��H�9��g^Mf!�t2I�&O�\�̓ٚ�EP�@��n;y����<E��ԣ�tJt����J��h�Ϧz�*��`u��T��]O�����;=�4"��(���9U�$:N-���X	@�K7�ιVe9�����7���Y�n��;M���e����嚞� Μ��z'5�UѺ��=���^��s���!��7��U�/^�7�9;�=������xF���1���Sɑ,��d���YM㬪�i��\?�)�w�y��T�`gx��V����\����d����{I��ػ(��S�N�A�9�1�1��l3�fV�H�g}�.+�u���m�{7��%4.7�5�ƞ�]�/��<A���$@[!����7�jR�s�k8>�I�����N�@O4�������������\�Q��A�?q��V=Y�E�p%Y瘏��:�b�{��GV/ʽ*f�i�K�5��.�򀤵�쁊�נ�	VR�����5C�]N����5�B�2�G}cc���ێ��U�*:{5�Pg� �˯}=����$�>�c�7�kB��n�i������<	(��H�e춗�b��5����&�Ydy����8�~c��_� ��~�W3��p�_�&u��ҶB�G�� ����UYPT���W}CP��r������5Ջ2��Pl��%դL��E�*8����/��j����$f0y�W��� ��Xb�Uy=ڭ0�zeV�FңWI�@�>�A���N�NTGQ�V�~� ��r<�^���bu.�]&��\�F8�r��i�Y��)r��m��B��p퇱
&���*'�s"*[oT$C�.$�1�m~r�.��{+�3�����9����~Y�sܿ|��:�YV�A�}U�̵�E�w��x��M
���豦�ʳH�2�K�A�˩-���z�^}�~�h��D�瘍�

��Z>onU�q�]8�ѝ?(X�U�6��ۑz �0
�����\� ���e�y�܂�ո�*�E	ābbQn��D�����������?��nn�e�(j ynj\�O���X^�j�"0�`8���<�7�7���Y�<->/R΋�>7>2P����t�]��&?�]Y��`,�J�t�V���7���^����7�}I�(�ɏ9�=��8��3���c�jz�^����3�|�L�8�R��U��p�k��r��S�JV<���Qe�x��Q}ZV�.Εd�\��M�X�&^�i�)�r��ǯ�ʹ��l�e��v�<�i���[7�bx5!g5;N�R�s�|��W9�\������<VJg6�έ-Ϧ;+F�D�-����)�
Fe�^̓�x��GJ�w
�5�	�e���?^�|�</���I��e�B�a�d��w�w)v�����-[�i���+��6E=���=1�u�[Tskp�	mT|lMrH��*���}%�9�4�e��d_~�ey~Q�ҵ�WTo(��+�I�W�68��n?����st���=���p��k�����x}�M�HB\����73��޺����}�ّ�Ɲz;��)A9�8�v����v{ovqі���������)�6;�P��'�ɃU3l����I��
X����Z�D��K��PاQ��4j����ρ����Tf7Q/��_��\}N����Ɏ��d�zM�v�������$ԩ��=gZc
�(�3H���j��R��+ORA��� ASB�@�6Q�Ǧ|&�V~���H� g=LRl��H�Ӛ��R���f �Y����NŋA�����a�@cG\���=
 +���$����v��׸-V�dU F_!����R��\�m���8��J��nc�J0�n�4����6I";i��W����[4\����!�хq�E��Ȩr#PSs��&��_T[���8Ԫy�#(�$򘏓�:l%�;b��Ĝ��s�3#�տ�������_'�����`�hf�Rv)/�!��k�j��A|s*#7�lr�>��Y⒲"/JV����^?���󕝕u�A��A�X��$] u3��`�#���=�ĵL�u-[�+���#�U�O�f��x�qCd�� �FL�D�ԓ{�^��+29�73_/�����1�jխlY�Z��{���D�������/_O|8��y����Q���mT�4�N�&G1`N��Y��L�B!5x�������^7�N���)���H�,\�w6��#�E����q�K"��x�55���>��x�D��B�J`���H�������pV�2���?�{��<u��p���g*8���\�^�u�ux�Ç��g�ށ�!�����T�{� |.?�T�O��e�k��lqq?W�K�h����Yq����������v[��	�S����:��,�3}��B(�H��TR�,�L.�q8X�H"*�2H����(IŜ�Mc�^��i뉍�O���Q�����ɍ=��bI΃�	|Ŭ��M4j`�Qʖ��׶C�J�~0����q���'�D8����h�(��)��a!S4*0��p��(�
[o�־P��o%X�P�I*KU�[<��� U�ܑ1���!ʄd����MwQ~�/�R���	 ��&EZ�6V�ղ\���D��588îc��Y]Y�����u%�J���k��cB�a>�Tۯl�"�2G��3o���M��/@��wU�;�R՜樕}�����,:1�Ċ��������4�̓�&M�U����Ы
�/ߏTm��FU�ZW Ȫ�'YQ�i���|�D���x:9r��x��s��B96�؊���U��	U�����E��!q���b:I<�A��~]�Y1�\�Z^���$���V�Gۜ5%�Zsp��gk{�lU���I�Ht�/@��o�Jx@4'NI��J8�c�������i��=������Oc���s�[��5�"qת�{Ī���T��?�����t� D�_�N��8MU&�_C/�����UK�pΙZ�����@ *V#+���c��a[8�<T�C���v�}��C��j�a��)�/���좊e�D7��RV�j���)� �T���m�ʬ�ͼާ���0﹪�6�W�'9(��cd��yo
���wX\v�r��.�4zrP✨�$)�(��(Z��j�ZT�1��&Z�O��&! G"F
���Qb�F�y�q85
��Ǖ$��P��NX��B��#��Mv6)�jҞp��lS��d����E����R���dSl0�n%rš���95FdOE��]ISd�$)Q�c���8B�c�#���� �2ډ.�EA)�ұ��l/��ٷ_���-6�$Z��v+z/7k{~ynW�p�'�
Ed�ˏ�U�!��>+>oC�4��`������cP/Y�N�z_u���jN��c4Y�A6��b�
��NL���)�s\�H =NYq����W�C�f2�� �ǈ�Lyͤ]�V���y2�?��f�����-�@��&Gm�4�_S0Q��*�y��ì�Bx���4	�yuk�	����M�7UZ#??S.z��S�~��0��_E�uB韃ﱎk���r\$������8��q�b�d������pcIߡk���e(��Y�g9R�p���gW��_�7_˯ϟ�`U�$W�y��<<��}���no>QA��]�ɔ����8��9�����̩�g�e����%X��r�&��A&�9Y��Pa���~��8�lG�%�>�:i�ա��/��7��Q��F2$�"�=tN5�k��P%0y?���ʚx$�j/�2P>pߚ���5`r��ZD�Jq���I�x�3I��E��u�p�E)Zb������4��H�p&���v�0���|6�ϖ�[�N#{9���c�q�{PaC5i�o��,�[�	����Jq�͹�=%�cu��c�/<)�aP�ZD��b����*Y�KK���>�0Go���ᐬ6M��j��5�=�2F�����٦$Yg/lu��ߣ7�4ˬF��)"R�rU��b�̕�Y$;�#nxV�3ٜE3^�֝Gג>��|�UU�A��g�'49Җ��?�w�{���H2XTX$�Չ]lZ >���� f\ê�w�I͂7�ȕF�T�MZ^�]4_V�ܚйV�e6��=�#-�#?���`b�i>��^�#		�@���!�f� g�y d67BO��k�8E�չ�G5� ��׮8�u�G��b��}����ʞoK����..6�Eƌ<T�2�3 P�}�3F����?.\S����Z�� g�'����$Z�vv~mW��n�#�� �`�uqA�zU<q�����sR�yShD��s������߅�������=<�1@��#��[�RX���;��hJ�㠹A��0�b�x���H�~vh����H��I�BC�o<"�j��$	���}��F�dOn���O�j�v�M�_�^>��Dple�ެ;/���='�ö{��b.�t��?q���Y0$lGN.��b�@͚3�`O�b���  ���t'��Ddn�ʡ'# 2�w�=ˢ�b�A=���{e�U��.ضs�_��`�@�z{��?��u��k�h��ׯ_3����n>}*k�A�*@%J+M��a�sB?:�Vv�\.^=����R�eeh8��&�.����\�9g�z�����Sh�g��T D���b�f,�}�����k��|m_�~n_|��dN(D�j���u��M���Nvy,�&,X[I���FO�_׊Z?�O�mra�#�| ���|� W�l,�K4Z0\�(�p��z��r�[�G1Ɖ;B�vOT�}�=C����89� m�SEI��^�����G�ۚA-b�������ʒ����β'�����<' )�T���k�d�ƞ�v��$�qU� NJ'~�j$�����Y�0?��ad'�V����.�r��ɼR�0��qQud�+�k�ٴIyP�~�v�W��9W�(���B�#ΰR3\F�:{�c%��p��eS|�����x_6�H����m��dh��IV�"��4Zm�g�X�,��0�3��o8�xO�P��"���\��z�0�`�����J���*n�E_LM�j�>�H�@��(%&b`i-�����o�=�r'��D`�rn�]��X�^�� ��aY���2"p� �j;�S�D,̘5��$%�y�Ì$�%�f��\���Z�wTŒ�Y�R� '�a1��wP�9�=%�>�>E<(<.�01HeCI[�J5�N�6��4�{�TS=��>ֵ*Z�f��I�h�,����U1�gdO�ɒ�G�^��J��Xe5�Oh�f0��8�6B���T�]I��t�
�Aa�'*~2'��>3���/3�����r?�)H��%�������0 .�ڄ��^�1#^���`�l�b '��)��]��#�����/_���qss� �i�fkȳ�P�cN%���	�U�#�r�|\�\��c�J:ڷ�F�U+s��𻹣��|(����-�y�W+rjF��^�UH�k��= ���DU�Z�G3)XĠӾ��P^5§}O���m����.���o����_7tJ9��@�D�o���%M�ЪJ�=�ў��n���we_*�.kZ�`VI�
Rc�y=]�3���{�z�+V3<�,R���pQ#g%��ߐ�~�C�9P]t�>�^�I�
�XׇQ#VCId'��z8�b��d�T�b��je�`�R5.X���|��4y?OC���X��lʑ`LޏmNǔ�nZ�SJz �����Z�X ���`�X7��ͼ����[�6��p�������5�h+��6�� 襜|<A�-��K'k��� qs����DY;ǸC	b�����DŅ�#�ׯ�p�g%�����C�w~���ەD�ű=��J�~ſ���o�֌��wmC?_�HM���9��Q	��)/�V~��B�>���x��&�+��*hF�s^��\��&��^D�0|,���V�'���6)*P�$�NX�H&�2�ZM^U���Ǖ�0���08��ᩭJ�tq~nis���-�K��X��r��:S��Ĥ��Zڳg�낂*�����޻��%��gc=&��ɖ)�N�Fk�(O��z��ั� �ñ��[T��;V��)��Ii^���T�]��_�� �5��i��ϔ�$�)3����6��IeExm��-����1-�\�d����=�by���Ώ%�L�R����=�(�.S�^Ʌ�w��jP@D<=�T�"U��{��^�;���ٯ7k��I���90�CI�,�/^�D�����(��-�^�u�­$��I֜c�x�$�=�j'�ƞ��D�?����H�����5�E-�jP�b���.�����z')�%
���[�L%G�`b~�f8�4��򩫵1Cv:*���0e�5~�#�z>*u��%0 1�(7�U�J�QR�=�4�}G�İk}�US7�d�s�R��Z�`�ltJQ���>�[� ���i� ���TP'sP؋u����ÖO�ZXu������4��
i$�Z/��]^��w	A�I=x)�G�N���Vy�5���8H��l^�z3xb���0��fL
$(���F��ע�֠9#����F�z�$p�II���QmJ�U�f}Q��ܶ�j8n4)�ӭaj\�s꥽U� ����Z"Jh����a�N�r`�Z�a�񡁈�j�����H��:q���PSc��8u\��7���ݽ=�=� ��=<>J��P^Z�َ�"M�Z1�L�"�X˲J/�1��6UR��Q��k��<-Z�dW�gZ� C�����+)9ܬ�?hr��U��ع���V�X��t�ChAU�-�÷S	n ��K�����3���$\g.�O�A<2��e�}�.A�㑕��d��f����Y�~�F{-h��p�p�sR�zs��+����=2����P����c����>я�*���V�F�%
!!�X�Q��SI���z�K�z�-�U5�*>v;��82�H�`��}0���qD�i�l�U���ڪ� J�Ԁ�K��㘃�	�|&H�tqNe�W�\V<�T���`��Q҆j�<9ť웥�h��G�^9�8y�[&j�VV��U� ��#��G� �
���}�v0�+6B�]����L�`�Q}&�A��>A�Ǿ��+�?�_���t��$Z�%Y~�Y >G�Da]����� ��f���{�����f^0�j�-��9�k�+{��`��O�So�*%����X6Vt����
�s�(T����k�=�!�CJ���bD�H��t ��{u�̙RP|���&zꑜ@��������1�j�.	����d�8ʄi�2��o$@����fNp��M�w=����!�S���?�Q$Y٫���O`�뗂}`5<��h����x�o���^2�q�$�r�t��'��Sw���ż�F�}�a�RX����XmJ��
����ǮLG�K6Y$e����:�����y0�� �-A���C���L����.h�i��#�� � �  &���Gu�p0��Hk���^ӢY��H��\����Q�͛y�ɫ���@��ig��ű^ISޒ7���7o��o~Q���>~x�_qSY�j�ioqSue�dM�|��!�
��~~g���<��<��On�E�5��g��[�H���)��T�E�M�!Z1�K!q<R��&Y}���64Tt
k��j04.0���u�3jٔٴ>�Q(�ʛ3p6�s�JcG:/�G�dX�䰋~�󔇹"�iD%G�}.�7���>�&���+�����	�'���i��ZP�|z�q���3�z:��j"u��B �D�ZZ�e�U��D�>s�#�<�+���d�+;�f��D�T1ȳ�Umm.%����lg��{Q�����=����/�'�����������%�ыE1S�H"]Z�u��_��c�����Ϙ'�� d�ׇA���wt�^C<&�{
�"��9���uF�b��m N>ӣ�'��/^<'2;�u
)`������a�����?��r��*��'�.�o;ՙ!'�~M]+���8`�+�Ӹ�k�(!�	��O���s��O^o� ���I��[�|}�ad@0Vw7Zh���Dj�S�:^$c4x�P�z��,A��$V�k���(�`�$��+ϕ�c���RO>�6TӴ�$ơ�Nܗw��R�=���K�F�Q��E�埜�	9��߿�'��c�������6��ugw�����c	�o	*^���s�ZB �j�P���X��0��r�%ɺߖD�f�$ι:�!-\�Ŕ�LJ�8%5�x+pcP؎5Y�~�R�"O�<�]�+�L9��z@0H��;%�JrZ���|60������1E޹5��t�BO[
���脃7ֈ����4��/M�#]�R3�6�:��%_��X ��,c��j~�C|� ��+JV��U���gʈ8�1,�!�g��:��bC����=�$����/~���{�$�NM�H`�?f_�D����ߓ�dV�2��s�^3V�ث��i��z�Ђr	{��H�ZV����F�,~�Z����-Js��UK��v�������U���mQ�w�b!x�6!3�[��յ�_]��⌉�6�oT��2�m%��fQ19�3K�O&����+�H���p�5s�Ig X��S��y�u��cG��q�C[aō�z!�l�a��K>h�M����񡽓'BK���D?R$�ɓfO�L �*��\���N$�6,ՅUA�f�[1�0
!K
Გg�H��I�ϊ�u�"�����?����at��<�)����K1d�9���l���n���v1��%J\Njh�f� xѫWF��y�����0��?S�@�k ��<2x$YOO[���#s_i������s6����PB~�;��2y�zX��[^�zS�0�SM�8�gƶ�9���$F�O���|�hE��Y�LDR������J3M|.�v�|<5k�)� ��j�Y5ҨfJ�"��w��40�k�x�B�f�����6�������W4�md���h�g���;5�s'�+����������pF�g�{�~�{]OG�Щ�JΛ��:�t�'ݳ������s�U�aƇ��?>B�y��|��B%��@���R3쇱�(i'*��5s�t�M�H�["B����W�T��V"|���$NH���+6�#Q>(��+���8�}H���������_�ʿ�p��/��\<�%�i�S�H��C -qbQ�["]��kp�اJ�t_�4{֌�y�	�-&�M����%�����e��K	W���b�Pɺ��"==XgǕ�6��P!E�*�{`�y˦�-FuZ+K����N���b5Q�N
��	<�WX�������K ���6�he����O�Tuo�� d��V�$Փ+qŐo�@�'�g�I,��!tP�[J�c�ñ$Y ��2{�B�+�/6vu��ͪe@�YOL�6k�33ӈ� {�u��m	N.J�|�ެ�ؚ�k �S����\*<����b2��?}��Y+���u�/�mҧ���GQyx�>��hk/E� f��<m�����0��ӓ(�H��5�CȂb%�;���>d�/㬩,�E�3�}���[�mM�D7���OE�@��G���U�U&m�՚������ ���T�Hh��=�6�Ώk����4���*q�N�k;W'"���S9�����z���J�B��b��x�����k��_'9��i�Z�=���#�m�;诺,�@�ׯ^��7/9������[�{��{���<$e�Ϯ��>��*���g�G��'��u�G��<�*��i�H�d���k|���������y�Ǆ��sP� �%���I�Jk��!EbtMWT���y}��)]�D�x? ���v�$� %�42.T��h�R�l� 	@bV#m�94�`it��뼔�_��bdm�IM��|�&9=ܯ=(�c ������^�
*-/�0��T�0�]U[�GG�� �����yq�hR�5'2�)����~?*��'|M}������r���|����R\��,c����f�=�gv9��xm�Y��~��xa�W��2��:!��愋��n��2�'tlz�����D:��-	e���iVFme�f���L� o:l�79��	%y��<�=�?���u��H�n������P"���_}Y��%(���h�/J�]+��L�yI,n��Y<nd���$�)�}U�uocK�-�*��]�`�T+l��*߸G��wj�G5Ys���_��L��~��0Q������+?[��ʣ:{�z���tnIX2�T� !�$�{;�>��⴯��F���I�B3�4���ڣ�SSw%E�V�=H�`����c��5���A���#m=;B}�|��n(��\��U���n  ���RL3j���yk EzO�$k4��Ve��lU�u���Zh*�Ȇ}9�����������]�u�T����{�/����>|z��{��/I�.�����2H�u��Qť�P`p�A{ b�l�ΦA�m��/�*��<6h��l��}�|P��)~		��� �6�q��j�K��N���GS�d$�=e��N��]qR�Pa�a���J�s� =U�t�ܡ*d5������=��L�>�=$vs`#�C�����)�ή����ި�zp*K�y(oƵU����%A�Hz@��L��ޥ�M{S��eYG�fA�Zs0P}���7vw��|>(�O.�5�Ep�'4�8��cr�G��
*�;DgR�'JT��M�f!zC��U�R :����$��k *p�h�B��2��I����
��� �^k*Z�wDy
�gJ�RPSE�Dg�JV���J��XN�6y_M%�� MلwiO��leW�%h�:#]Փ�s���DU������.Re��d���ʱ�-ǵ������^�Y�ť*��Z��$0άJ��WPp�V%�$�k�3bI�~�MO�^d�8�h��g�~o7�����޾�D�����Æs�XQ/��aa���Th����Y�x����b��g��}߸z�D+h�a�(��yЊ��!�y�(b㪦J��c�k��.����QxdI �Vt�>��Q�IT9R���1B��yyi���oʞ�\/��!%�E@�+�LtQ$/��T �6�����uyn4��Q�$���M����l7�ʞd\�F��\g�����{�D���GrUޫk�! ��\��Ij_��H�������P�g��%�(�7%�zc�^~�$�u��Q�J���?�ճL̞�|�jaG��g�+,P�&N#R���Ŷ\O�Wi�Ť�0b��{��f}F�%.hx]I��.�Hy����%�: z�Ʋ�'X(�A׀��1���¹P��Wn�-�;&A�S��ց5l%b�Q�-A�Q[t��'� �)�dmg��U����?DÎ���w�{�o����R�XC���d��a���_h���b9&�[�$G�fb$J��,�ţػ� �I�X-=�F h�����\��F�UYˈ���ѫ;S��~��K�S��`[b��r^O��@5lOM�5Ɋ���D<bf{H]X�Ka��d�nF	��b�����)�:X?�M��QY��9�#k�=�(UH?o�UU��l�6WJ}���� �׶�EB?�����T��9�\�/1uog`�$�NW�-k�&��C� 	2Ÿ�Һ�;�%D�y�ՓY���0�x0e�Hİ0a (���%��HА�V�hdY�4�oQ
|����=E9x	3��٬��� �WP "K|1~m��6�Ϳճ�Z��?_�gv�@R��� �XX��/�Q+�F3�`b(���pP9���Po�����2��1�����}	�MF9���F�7-Мg��y�J��	�d��Xц��O�_�s�Ƥ)�\@�v%}�h��D�H�d�g6dU����M�ڸ�QTW����R�,^�)�|(��	־%���l|���;��-[W��h]��d��]1p�G�tw����=n�0~���7B��Q��qt^詚i׼gc�m,�Z!�5���90\�,*9Ut2g:�p���<g@b%�Nmq���.-�Kb�8��Ԩ*��I��Ps��c{Nj��{@]��%_�Ag��Q	Z�HK[qb��'%���j�@��G6��q�Z���d�}��@����=x��v:�	L+;����*-
��v��|6�1;(1� �/����^�ib.�	IľB�9�\�S�UF�OQEa�Ͽ16�.���wamb��_.<�j��i6W����S0y��q,�ۂ�(=��"WU��p���:j>3����HO��;��9f�K�_�� ��Lj/*7 �`[.1�ƕ�Pт:>��$�!,C�S���9&��]�΄�Nޙ����M̫�9�ꂑ����_,���b;�P٨�j�05?�;��z��G����Ƿ���7�=f�(=��ơru�c%��đ?����ڠz��#�$�:ۊ�!k�U�ݑ�<ߋ��k���t�Fw�k�L���䪧Gk��R���cXQèҞԟѱ�j�cP0����9����{�ȑdI�@
jVuW�u��}{���̾�3ӣZw)�$3��03� ��gϲ'�,2�����\�/�����&
:�8�N�G�S�^�}�g���'��G��*�-R[��CN�|��}?NE���#�h�f����y��c��z`�v�G���y�g/���?��/_�/$�>��y��k��@�w��A�7�|C��ӯ��Q��e����q[�C��(.�0gc����@��MQG�s�[);e �N?T'��1G��������	x�N�V���y��Ǖg�&�����;�2#�-K�+���jթ�[��
�)Qe�6a-PH�@��k `��r����5���u 2�
� .�S����'ZaJR�,G��ǣ�y9�E 	{��,z�"� ��,��I�1��,p��������A���/�~�wp��^4N҆9yYB$1�n���y�I�R�6i� �{���!o�%�	�s��E?Jl��Is��H�aN�c��糤m���}j{q>S#8:�,ξd��ZO��0����z�� ��Dj�| C����P"���S�PӾ��{D��q�EmN��O�תY�������u�:Q(v=?[���9#���w&��Ņ�%�n���?*�F/(	��Z#�80�˱ZS�J~�O_Q�Ҍ�����Wѻ�$]�,eJ���x��Mtx٣g���hM��<9<�RNU!1%v�B��6w����vy��=���)��m�>�?��`� %XP�����:�A��� ��!�k�*��������|�)�ytІ�mra���^�*�i�H��z�t�Ǻ>�v\������_����~����� d�m[�_��t^�b���hwh}x<�g��#�?��t�k����?���iN�@d�_>����ش���V&ֱˡR�.�#�ЗQQN���]Q�2X�3��}	9W�Fk�&�e�=�z���A-]�	��ER���!/���� �ж����X�t\�T�,P����f08�8�g��x��������.�a�\O����,�q�&"{-dzdM�=�̗����mH;Yy7�hr��P]`���b���>u�c�~싒b�����th�P��k������pN)��@�J��џ�M])���d
�P8�_��/;� �5�+�`�b'�a�8� @�bZ���9 ���-��������E��G���,�,`p��;b�vl�G��><��&���n_�:m|�-m�7/��vPf" ���:�$���`[�`��X���9�:��u��(X���az"����������|k�}�����-)�����#��L$�$̪�V��E!�x�q0"��y�u5����u����</��N��+g5�-F�,���JC6X=�|8Z�R��<{����91+r�XȞe�jSZ\6p���Qm?ʬ���ܹ�7�>�BQ��>R���u:K/,��~ó�x���
��N�[԰h+��/g;�}�� ���é�#��DlL_kc0��'�a��V��㏢^_]���� ����o9��;�P���Q�V����6�&����ڻ�'?��FVhH `���h:K�ʔW�������#��H��w)��3�8��^�땉��S�_�L�P��q�l��cO��f-�{��'���pW��Ș-�	������ k�H,H*�y�D�3a-V%��
�p�R��k�UǞX���:R��(�^�gt	0f�=�[���
�JL�8������A`�=2�GMo�-t��N"P�T��-h)��e��{\��X���q�=4v��'"E�n��L��lW0\ȹ�$�)�FР*:#3���X���b :C�����acۮ�]wb���[�'�h|^����::R��59����W��wzm�Je����y��<|E��y�lQ���lnFdy#1x-�q���xD'�D�q�����=�zPCߔ�_ܲX7C�S=Ϊ����߯l[w���_c�\|ضVH��A�3Y�x������D�Nj#�(��L�����l����Jrw�����@	Ϻa+�AǙ�Ӭ�X"0�d��J"sb��E&���:gvu�B�Mu�� g��\Yó:�+/�W�Sdo}f��Ac��<wrpdFԛ��>J�P���Pg�>޿Gu�2s�S8I��P���└�	��;�����{�����z�,����q��H���7�>��\�� ~W((6;HH?��N�< FG�D�p��3��x�. 0֏�)���L���]�>�[I�¢���"N@���~��f��6ƒ�F��#GR�@s7�#`cM���Eq�a��k.1M��'�ſ����x�4���}�nM��k.��Ȥ5 k��z>P[؃��yD�T"��ش
��V۩L���1�Q#S���k��<WQ�j���1e6w0�n%j�r��Ң���.�7�x���ܥ$w�X~[�m=o��Ɂrd�X3�@ک�*e��͑���5��P�����1����-���r�7��M���������#ꅽ�A}����+TQF���:/ê��jW�7���a.!jS��S��
����Ƚ���R�,Tj�B"^U��I��0�3c�c���T}�ǶvA?�z�p��~��;��o�ڷ���:�?ػ�(���,%F8�P�&Iգ��� ��D�!֕��{e�x��� ���5d��z�p[��*W�#�Q ��n�ˣ9�ʔ�^�k��9�J���+:�E5�,gbψp���8�Q�� ��q�@I'�tD�1^� ��A���g]l/*��3�
���F�w��	��#���T���1ꘊox�c���/ڞ�~H��,��(�Y:��"@��/��}���ֿHr����?��*��p�~���.��P��G2Zp����(�]�m?ӎf��R�	��+��N�=�K%b�O�h)<�x����I����w�&��T�Kz���T�<�^*y��E��*�xwg��{[����^�ֵt�����}�g��
F�;{��j�^��A�{t*q��� ��o��ds�>y0��)�U�R�'W9����Y��9�������U�O�s+��m顶:&��Igt��OI�{��w�)۫f�#�:RGf��!�`�00� �#z���8z�z�s-�%J[���k�g/A�����T]P�W��LX~�k���b$'�D�r�d!�`�?9c~�'�/��Kw%�;W�iރ5[�&�
uaZQX#�=�F�b��"�x��>I����4r��:���J��_��tnQ��%��f����|M�sO��K��������u4ޅ2����׆H������͟�k�6��f�"/�b8�X�1������.%��������h��i2�>V��C��	:t�N0��BՇN�܀��}�&�I���	�#��>T���4�u���>֔5]������[$.��ʃs�D������)�4�G���Ϥ����r�1;-D��ȑ�Ʉ�Ի1d�;U�ծ�N�;�B;����ݱ>����T����_ޠ����@���� ����,P�z�H�CJ�0��� j���s�8��P�H���s|���\H��U �o��8�����{Z�A�1�rP�:7l(N��,Ce$�Yi CJ����{�K�0���6�I�`iFJ����]�ߒ6|����� �å�����Q������­`5�m��'�붙��;5��J� ���Q���wT���}�||PB
�9�%v��j�9"�Ǳe�� aNy^^��r��mk����X��ř��Y>rY������7T9��(�Ny�>U
.,�)�I��.f6��T�TDL3�P�S�
�;.ګPf�Q��e���z7�Q����H��bO�l���ڋbw��
�w���d/���n^����K��֐R(U1�����`���KZ>�ؓ�w�Gm������?��?�������_��W��?�I����Q���68�#���d֕A2ֵe���&������{��to�g�B������1����M�M(!6B�CV6�p�NWd�=����I|�՞��Z�!��v���KP�t��Y��Cj~�0K�*��� 0=x���z���l�1�n�޴/̙���ո�䈂��y���m��U��v4���������>@0���j������ATH�����v{s[A����� k_�d���+��^���֞��&kʠS��&��19	-�O+��V�tD f�>�3XC�8�N�R ��L%e�/�g	�p=Իl����Uy��y� R�a|�w ��ٛ���8��{��I)����~��*w�F��*ɤ!�߉%��F[7��KZ����Sv��2g%P�Ne�h@^
}��e?��:�O�^���u����x��H�ĹI&�#�^W�	5��T�s'6�h�AMԃ��*���T�gZ����t�:7uBE4�?���;P~_*|q.�(0���Z���C�Z 8!f'>�ir�����J���3�@#x�3�#�p��Bai,�Pq{��K�N}a� +�(c��h@}E��Q�E��m���max�kv\� ks����~6��ۍݾ@?��`:|�:g*��۟N'�4|��?� @i�����]<��(e	����h���==F��yv�i4d�@pe{���:����C� �Y콼���,OU�r�����#��z['�|�!� ��lʃ��f��M�ұֵF\<��0Nx�h064��A�#@��|MJ�f�8�O�i���08U����Ƅ�y��(��T�V�=U�$Äz���z����'DP��Y�Q)��s��1χ�چ���,Fg�4ydCJ�"�+�R�`��# F�k�e��
���+$ o�e5x֖.C��.wl[P��H���8�a��;�!��^Y��k���8��+���˃�[9/��;'@�������J�ЅhF3�NIi
E��tՌ�!�[��/v�H�>6Q�s�G}��s#�H8�cO��3�w�.����{cMYb�	�E�=-Ԋ�F?�}-a�w��W��(f^\���m8ԋ,��S�u��`>z��q���� �^)'�3��Cę�H��\ҧ0.�Xd�ln�j�6 �~ꮅZ~��:�:��S�&�*��3�ڇ����qy�{[�ŀ�g��V�lw��}x8T�����HN�������\__9u�7'�^��(���#T��(���4<(D=���=���3Z������?�Ο��QⲔ�Ы�����7T�)�B��:��z���υ��}�(��i^r8>!b������E�Ȩ���a���Y�u'Wq��w��g)d(�'sa.lo�}-`2[X�m���t�ȡ�}��s�f����!������E(�_�:����5��x'f���s�$p�PAYߖD2M�V#��Vi��|�T����� @g�Ƴ�
QS�җ��8?g#]8w��`�b��-���Ai�̅R����FA���%�cm�#�Ի�K5X��^����E}ĸ�+O2[�F��Ȗ������M�����88b?M%�sMc]=?�����*�� ����*	RMb�A�]����W�o�Igų�%�Z�<�����KJ�	L�-��4Q�Is��s�T�@�S	t���ߌ����͗��ī&��}@�up���Ț7�o�^��$��`U'���HG68g�܁��� 5�G�u���j�)�t�����(�$���S��&j�f�lGP<����7�7�m�ƒ�m���.X���o���1E����;|�%+�o~{@�~}z�5�]� )P�{��8�k�Ω*�#	���kyt�?}ɡ�%2\���J���o�(N�|������{�{���^�O�խiC�9{X'4
a�&�E�s	z��rBfV�5��y�T�]b+�o��:��/����{�`:1ߦH��p]�i��i�(CV]Uز���p����A]�����Æ*@�gv}���+��H�h1��MF:�N2g-��i��8�2�f`r�!+.��z�'�Z�i,(Z�HdϬ�)�h��C��� y��"�zT(��45FF���uXPמʚ�2O�K> �)��h(�wF�
��8��<��Y���
��
2�*�� �4�~��-��X��h-����,�X%�7a.S�i�1L>o�|�v(d���j_8�y��E�Ii�7�kq ����%���%��/��>)�:=�����Ȅ���X�1R� �d9L}P[8��܍={T9(ˤ-�M�X���ߠ�Urʂ��g�`�*|/^/���͈��<"<�a#��� ���]�����P�|�dы���fl<�:�`����b���@A:��Y���}�	p�`���v��tə���ǯ�ޏR�INH웈�R�i��� ���>��h�];��,�Q*�o�+�z� ho�_^�3�nV���^\]?�����l���Ȱ�J�T?�}� ^�SS?��3����`?����y�`���ZG�GzY:f�rRmU�Y��E0%�Tu�(X�;����
�3�������hw���gm�W<�Bgi�\`�X�3^MŊ�o����#�*�O�&њH���:jf��S�P�4�a��<X����Q��e.VT������?�^���k�����6��"R��g�!�X(B���ym�s�|�䎲7ԆC��ϫ��zV_1����[��vd�����ͭ������wl�Φ�!0q؏���]��T�@����if��8�j��Σ�m:s���e����Z�N��(t�PD4v����QBb����2;��� RGR��AA?�r�({�z{1a���UG�	p
i�U��M���fmW+�������:D���h�Sh`���ʨj�R���ˊ+�!1�I���ͣ�Wֹ�)��ɛ�gǺԀ��I�}*�]˪X)'���EW�lS������X����.|ΤzG�桔 e:dA�
O��R\NC�R��/��c���R�ز���*	E�~��PA�qRfUBk��&��9P�A4����Y�[ ̧�	�e�,N�v��x��5�������1yb�_�|?��_��
�!��R:��tV/Y����  Q;�tz�,����ݶ��r�θ�����I)Q�#=�Y �6-
�A��-WHwN�`��"ʒ�>����)t�T(�tl�
��� D����%
�N��?�}�����%�K�b�G��������� �2$8'<֊����;��G32�N4�T��z���{=0�5�m5�8XQ<�Z-Pd�#Be��̩f�}�oʙ6H�����5���ӻ�U�O�'�qr��=�9�$Ox����F��;�.�KL'���NB�Y튑�z?�{4�0`�(2Y���J��\xx-t�I�.X(�>�ы>"!��A	�_+
�M��ŗ�ظ
dk��螱�	s٫�\X��B
�<nCnB�h�Gsr��X�� ���t�0'����T�Q�+ҶȤ�Pc���R�&}��,��9:�����j��q��h+*��>+1��@�c:�,�c޶���~�u�Ad�d��;���.X�{G]����]^^گ@�Ț�IA����*|��,#k%��4�L�8ˑJ�׋J(y���`^G�}%�5��g"��yM����2���� X����ܤ񶔼֨x�I�&�����Ί�8�6.�:��N�L�Ank�����{��#�gu�tf�9����5�h�ժ��K��5/wtnQ{��v��V��2��A���|A�@�B�.�?|����~� ʁ��s��y���أ�q;YJ�O�F�WD�J�zY���,m[�"�e^��A	�����<߹�`�@G	Я�cJԜv�����ŉ�_�<l�W%+�!���_C��rP�M*dw�u�ʹ�(pތ�����f�{d,�|t�zխ�%��% ����=�h��2:��k�����5,�渻�1�t ��I���@RV|�5"ť��&�hɢ^.�P�һ�� !�/����@�ݽ'�z���%2XW`������?XB�u�P�.����9����?�����S�b�M�z@qے>��+�4M�I�4�+P������cggkR	�H��lv�5�1�70f��(:T8�S֎{;�G���`l/��V�������Y�mn��������Ϭ۬��s@�ݣ�:�N����
��a;�sL�	5I��s���8zVG=���	:�6���h�.��٩5��z�~���~�J;�l�+�[�9�~\�g����OV�r�:6+��0o�1_��m _��z��
�����;,��˯T��c`H��w���{?��Gj�u�\?�a��_�s ��i�xU�۷H_vA?+�� �R�����kɸ[�&�Y���g?���~��ꘃ��V�f�8l������~ �����2�V��qO�3�:�:D/QgD��N4]�<Ç�Y"�9��Hc�p��?�Hm`����(Y�V�q�������Z�w��a�T�ܠ�P�Y�by$�/��M�q%�U�r�X���D��>��I>q �	�.
�+kv=����y�hEg>{�$�kv/�����l��~�g��*z�C)�8����)�߉s	S4߽���c{a�ދũ�A)է�F�x�����y�{��&��au�LC5��
��#ڋ��$J���5.ku�_)s@�����C� .Lj��jH�H]�k�y�c"�F�V�4��/�I�ʞ�g�T��#�D1��ܘQ�=h< Up���%���<��A-Z��!;}�h�h� ���z��"5��\uA�?����t?��3�S�JM��m1���+�]O��Զ�ɺ�4�5|�?|ۅ5Cѯe�h�)��
�r���z4F�&E���Zfp�����#����=�h-�^?�!h;�͚�6y�D�_�|a/n_��	�e�Zu.�zbb��CJ��j�N���k��ʝG3U��=��ن%Zp���������H�k4~`j��6��s̳Ys�)���UHW�p���ǁ�5*�}�=�Ӝ{����]�3Ǐl1)�����NL6���Yzd��(z%������Ov��"'��vκ����Xo����=�W�N�8���Ǉ�����W{��]�����_�㍽}sG@7"S����{m$kC�2�4�.5�m���`��4���i��h��9+[�Ϩ��7E?��*|e�0O��e�ݮX���{�̩X�u79�����z�ǵjv�@ո���A{�Ƥ��!�qžc��{��q���n�Yt8�k̏��P<�:���u��c�6
5�nl$���%T
9�^�I�Y�t�����:@&����^��54��b�X���i�w>�Cؕ�������?p�!����:-����8�=�_}i�_�F���`�ԍb~_V�t[���Mu �q�Zd��$�|8�t�<��iGS�ef�4�o�(*&�zgda7�#k�>?=��K�q -XG[�_��y"�:	��SU�<�Z}ꢺ�n�ɥO .��;y������}VA'������/h�T찬�Ӱ��H,����T�:\Q�y*�uՀ UX9�B������!ұ���`�����E�o')BX?�5E��������.L4�&�x��+�䄢v��lm09�6�%K��d�1��hA���kA_> \P���.��/(�����Z&�7�	[��|Wk���3�k���I!���dL6�j�TFo�������Z�1��{
�I�+ڑ�
�X;��܅Gg&���`��S;_sk�lb��s�>����~� �x=Ԉ��S�>(���N��@�*�����f���Zr˞U�OR������i�
��0�!����l����m}�ȚgU:W�46yJ2��+���E�/�OG�xl��ӯ��¿����3��0��o�L-"H�s"jPz:�}��	N�(�<�TQL]�� ����9x�B�c���������{:�ח��t!�����F^i�˦"��ă��|rzD���/@X)�٢����N�ODw,r���YEA�86��&f6ʤ�P�
�\d��)g�o���w�[ׁN��ƕ�Z��|�؎��{dL��Ŧ?<�#\�='�X'�vf�<S�莝PO�N��;wz����%��G���X3ɍ�P�ͳpY.�Pr�v-eϰ5�x(I��&wV=�Q��={=�Z��\�����.�wCۇ~�i�i�|}*PP�dWZ�x��~;�nM�hs<�}�����i�����y�0�����@��Qd�u``����}��� ]
�z�L�����Fd��O�p���p�EcݯV�Դ�/�c��X~��v�Ĳ�!�Y��'H�x����@WPʲI2u��Zn�6����?�Q��h s0�0�ޘl�񙋚.F�Sq1�� ՘�����>���V���������%��6*ۏژ�]W���� ����I�~`��gڐǇG{��d�˯�ڛ���ݣ�ywo��=�ã�AR�2PA�� ��2�����,kNYL˓8�z����9�_�� Y�I! ���Ͳ<�L���t���=���Z� �B��P4S�9���c��lp?�6��O\GV��`ˬ6�[�/���06�!�4+��ﴧ��}�m�K� JG����3z>	4��l��Ǭ\G��a8#�<Q�a�}��L�ڒ��A�أ�y)Q�d!�$a�9���N(�#��Z�h(~��״+�������ի���_��_0z����ۿQE>��� `�Pl���'����M)�̞�>�����3o�^{2KU�:�Ϋ��۳sC�ʚ�Y{PI����p?#AȞr��z�U�̌g��?��m]�k���05UY��U݋��v]��z'>�*�ҙ�����cT`��J�-�uoCS���T�E5������k�����}���>���{W�B��(e�� ?F���l7{�&֕!��N�ulW�K�� ���2)�e?$yAJ\�9j����p�k��'�����{�����?���~���qow�~��ZFm}<���2q�ꁃJ�2D�-$����D��H(�#C��-�P�,ԜI6����}]d�yR��<������Zz�~�H�W�+��؟��g�TX ��@f�-��Q�$SȲ;�c�	N�D�5o��dſ�E3]8�}N����"b��vVZ&����^��p�qPm*z><�z�����?���������^��NJ���fW7�H?'�teW��^�Jy8�:��m2��t�gD���|T��qÍ��;�ӿ��F��_����N��<�g*���
*������f?4�"�֪<�3��]��a3#=]�gx�/b���h�%��^�18O�$Y��]E��������1��1�{,��~�Nēm���`�{t]D��z#rv��Ԝ0F}�b�d��5V��L�5����~��x.���'fWێ�y>����+{uemN�n
��Cp���[oJ]7���Xg(/A�w����� ��5Z�f�}v(�f?�����W��bww�U�rT�zi��Pb���ƿ>�Q�d]Ry�S��}�cvG�Qw�h��cƚ1Q�"�g	w�F�ճ���8F�Tɹ��F��,>:�	��jW�Htc�Qs������`���G�9������乹���>ze�y*H5f�	�s�FG���k���tCp��s%M^�B������or��S�����} �L�mD��u/����'i>�<���7Q6� ��yn���!�P���!����G*p�Qkx�&�`8�`
9�]�?s���<�th�-� ub(�9u%���s;{w��_�g�~-HM�AJ}w��j���P��V����p���$\��(I�:ⅉ6�s��ɋ��{��9�Z���t8��w������8ںC#�l����Ѡ���WЅ�x�������ir}�h�������rя�~�d� t�#{��龋2>U[Bm��^��6{4�+^�"#yA�r�V�[F���1���5�D�pda;�bD��=��
��*��o/� l�� Jm�\Qo���B��/�'
I�rI-B�̋joǃ��s�
��.��d�l�)���~��+�=��T&eE���NR��yo�V�� ��g �R�u�/W�v}��9����M\�Ϙ���L�2��M�� H=ltvj�Si<�ieI��|�=f�ʥ�E؛�b��*\�5�����^�������믿��*�ze�W�T����/����O?�_~I`�����Agn�L|�~�A�ы�H�ݛ�L���^�Ȝx�z��n�  3��4s5W����۫[����m�kvX;��]�k���>�pF)0Q\d4�=m~N�빑 �P����R{�>�3i�G־U���go���xl]��ǹ�5mn�g���8Q`����vOϤ�n�S��^�����&OG���N�GCo5�Q�=�j�y]����%�8?�+�H�1��뭮ɱ������� s+��́�ȴ����_d޶���+=%�0��v��ڢ:�%�4{����H?R�R�L��#������cpQ�����gվ��<W����K{y������uvk��{������ݽ��8@,�����i�
�Nt�Z&��8����H�1'�Ua����w�1�{��hMD)5ԟ�t��P#���j��̼X���5��XEy����D�T2�&_���Q��@/������Ͼ��/?���6W�x����#�f����[�ҙ:>ն%�.~`LοV=Hߎ�8��"b�NDA��J-(�E�=���&�w�@z��8�~������������ڼ���"����<�a�1��$�ы9�p�Nn������l�,K�g&7���ema�9j>o	�3�;�7ώ�Ö��i�֧TC���r'����#(Y�R����=��j lA�M|!O}~���m��C���=W��8�!��ʧjh.e~Fu*���3���N�[Og��b�s��A��Δ��:��j@�Q4xuyE^5c�Y��F4&�?$�	��e�A��0y:.:&���;�V�5���z$GO�5*ʊ߳k@z|�Co�ڪ�,�LJ
�4�[�>N�0]P�N�ƈ�D̼���'��ia�;�B
�(�۲��#���OWvjo�+��bs|���G?���b�&Ч���?yA��D�`M	p8��ָ�Q�?.�\��sԂ���SZ^Q���]l�:�ie��em4������0�?��!}Ǧݼ�zȦ1lC���t��@�{��������9��Nt��F��,���
o��d�<�����:�͖��t��)%��s9�̓��9��A�g_N>���X��;�o���+H������9�S��t����xØyeH�:Y��Gl���s���w "���:) Z���I����=*��xdO�jk��6��aD�3W̨O̬�2g�b/�q�47S�řs1d�`9���;��f;Ìt��ɦ��˹�(x.8d;GQ��ښ�m�$%:W<#p'�]M�Ao�M\;
x��]���W�P���iGq+\ "�S�6	�S�U�B��,eyB��׌Z��.{��ގNw�5��65��9x;�����-ȳX]�K����� Y�-5�țϕ�u�CI�F(���=�\T���?���Ud�^��_�b@��￷���o������ݿ(�0��77/(UԜ�\�2:c㚂T���T�|�uq��M��ո�J6��tLC��#h�(M�&��/˱���{S�p��9�9e�,��l*,�D���A��9����ωV	�G(�>���@�t����9�B�Mc����G
@���g��Y&��!F�"�#O�27@E��d$�!~�����1�`N��A�.t�
�=6=���:�w�����p�+(U\g���g��z����_�����a������Q~v�fF,j��6;�\�[�W�O2U�V�zT2���4�'�0s�2q��}��ȞΆ�����`��-�-.��>N�k7j��PV*�
��D����ƩI�îPճ����zm�|�MR�d�<=Nd+�������c�#�#�A絆f(���' t���"��+	�%ݤ��Ο�x���j,znD��B�)c,���}�R�_UC�N��o7R�d��>$�o����� W.J��N��󍿰+�G-h@'����K��������b3}В(�+�_`#��|��FqT���y��*���6?���Z-f"�#��n��K(�I��"��ڃ���P�S~�NDVE�����#
��F��g����7k��U�a=|]PE醑D,bn����ée�SE����qx"��Z<�u��˳3x���#3�N�Z)ӎe�� �H�_d(�����? ����{O������3�KS[�vpY̧�ԪXf'ˁ�VWyY�P�Ru��vf�HE�[0���ЍT�%��������7_����(�ĸ��YjN9�ָ�F$te�ۇ����pX!�0���u�GNN���l,3[�c�'��^�.����s���ͮ��޽{�h�n�Uat-,f8`�ԅ����D/�I�+�ܱv獁�>�r�;Ϫ�R;?�������k�,i�!�߆~pz��-'���o`�?��P�>��M�uY�ȞX[�Qo5o�dK���7Dy���Ś���� M��m���1��?�����T�P�P�'�X��l�'����L�=�&���L}�`%G��1�O\�-�
����/� l����ӑ�1n#�������p���i���+Q;k��f���Tg�v�Vj +��jñ˝@h|�r���|8��5A����ݪ�\��'��GGϲH�P`.��}�F_3�ƥ�y�u���튎P߯:��#�Pa�rS����Ҝ-�D.*Η��[�Śk��>��J6�ZmZ	 �����曯x���@���~��~��'���o���{�M�^��z����L񀀋����:	6�e�H� 2���M��N3(ի�5x�=��Ǆ5�ZEM����L��1��D���m���q���N�f9 j�x�GƵ����^�>������숆�R���^��ܫ���u�+׼�
k����8�Aჰ��S���;�&=���H��@�JTY��Y�g+{��TU��������=�ƴ3� g+���\_��� v��+H�c�Y�gAV�s���A�+���	�'6����(1�X���A{{��W�;c@�����wo߰�6��k�b�L��T��tOe��lmQ L�ț/�=�J��@�|He�p���u�(��C�w��y��sۛ,�=�7:T��K~�*eR_�`.3��w�qײ���_BX������/�S@������2� ������jI��J~��j��&x�f'QX�v~�@�n>�/2�˯�쩿�p����Щe� s �q|�Ru�� Y�n��1Q�eI�)Ü���Sy6 yV���Ym�h;��4e�df�������E� Vs���Z\AʿX�T�ꬂ������t6n[�f��Q�%4<�b��F�F�u#���T?q@�z��S�=�����:kP@�DT�~�:��<��t,n�L��c�cOu�K�TC�J \3�B�o���7��}M�V��A���2��A�2���y;ؚ�N@��(5ؔ�3�i�v z��㨂��(e���=�8�e�I\�"��e4�fܣ���Ve���=� �Wsd*r��KFj^�3���\����@k�s�
<�|�~h>��＾c}�9����[�Bc�v��y�<v���;���}�_3�*-�a�p
T�P-�?�S�)p®;�W���OZT}�M5��lzڟ��#�_�����Iʆ�i,1��ciҶ=#�S.'7�b���)m �e�SjM��B��	�DDpP0Gm�%�k��Sv�S �.������Z2/�$��(��Pe0r_��XiT���u��n~���dKP�7��sv�K`���M:��ɦ�)f���`2��)����z�v���"@?N�IO.^��+���M���j�)���Z��$����nw���Cۘ�?��64=�{ `�|�3�0��l�z��MjlYN/�O�� ��R#�	m.D�F�N}���
d�&	m�F�K �PG5����3ۼY8��U��p{�s������B�,�\���jR�_��(�#j��&�4� a�U�m�*(�����tLN�E�.����L��΃�8������H����嗯�swU��
V=>�l��H �����~��5Y�o�����s޽{'I����I�!-�pZ\�"��~o��<�ػq��Mr���l4�!�j�6�͊�� s��q��e� 3�����?0C�׭L4g��<��}w�hv-q	x�8�7�D|vkW7�Y��������m{�Q?����/��9k�}�{�==�F�h�R�u��k[_��_���g��!{�I��puy�u��=�!��w�G�٦��Uw��5�g��:����`Ί=Mq�@�uy����E@��i� APjWk��Ӹ�:�k�n^���-�
�λ�m��6�`�[�hb}}}cW�q}��n�%�J�~v����K.*D������֐��P��3��C2V
���<��@vD3ݫ�uFYR�Ȃ8����j�ԟt5�2��=f^������W	�����1܋N�\���J٨���sy�⥽�:����Y� ����h��J!��s���d� e%>4��9p
�D�0
-���Ha��a:o�	dš�4��\pH��Q���_R�TE�ձ�wj���j�V�Cu�w�>ѱY�
9����S�yz� �v��/��ً�I�����Yi -�~z���'�*����s����-W0ֱN��>Fә���A�Z7sO� (JA������t@D�]s<EZ!m�2��@TA�XTs�O�I(f�u�t��jK���&q�	��5��{�����
��]G�)*��3�.�ݵݜ3* c p���\�d��Y�J'�/]yZQ-0E8T�:���+������A��X�w�?d�ң�Zx�fD�\�GȫQ  ��IDAT�U�m����)*
fm��
��x���qm��Ώ��Ӻ [8�s�>b�/?�by.|��*x-EPJ��627m���K|���>�~݁�>r8�#����N��S!����Ji5e�wP����\��D��ųw�I�M�ԝg�s��T\%�k��0��Cj�y�f�g�G �X��H�L<�WM��J.���#�U,5
�.h�$���[)��t>
�jr�̞Y|`���WV8��?S��R�iw�'}Ʊ;�~k%��&�6<\<s>�'�|�>րI[;� @�F&	�Do^0����	�R�/f����=�����ɰp��W�����"����d�W~�p��K{CkQ���uJ�A +��#}��N�+��i���:_�sd��:@���QP�*�B�/<�.�Q��ʅ�k�����+TE�4:�?z�B5OF�?�/�P��	���i��+zܡA1��М.���W�Uv�[1���;(������J �b֬c�E�;��K��Cf*� ���� a3v����Pw�3c�|��0�ב����E�A���I�鷞��|�ff��9�� +����f��������D\]_�zAgx�'�z��W�\�+$�1�o޾��?�GB�,8�:#��@�%�s��a��Ѭ:��(�a�ȄPDv+�G��B$ �R�4J��Ÿ��N.T�Ybֽ����`����3s�l�1X����;�>�T����~m�3PMuF�7�� _۫/^�׿{M���B6��GR	?���]_\������>P5���T�ַ Eg���W�! ���i��Y�Sÿ����=�0 J�[����֘��4�?y�������=���T}�g�(�|���k T#Yqssc7/lU�����3{��������7��o~��
.!�t^�����_����g����r7��ͯ�5��?�k�ɷ,�����
ؾ>H�sQ�hV��Br�ɳɫ��qT�/6G#c̒��k�db(�.VS�����\{5���g�]
�N.*��P`���X#��y��czu{�q�\��\=�[&d��2��^���g�]���G�,���o��2G����90�^}t7��L[D'=����}E㫺�_�^1��:�X�0,�rvF�9S�����.�g*μx������XZ.�@���ZK}��'Οi�;ev����I~h���%m�a�-��>|y'K+̫���K}���b~8Xݠ�]	��?_�oο5)<ɰ:��N&�rR���%�l�T��g��="wu�7��}���Ohe;RcDI�
d���1K9��>� �Ų���,]J�R���ep�|�mJr���U�*�f�Y�E�Rۓ������|) 623�=
�	�(�	��K�N��:]�(�()�!��W=r����oK�ْ� �������I��E��X�]�Axע�Y��x�`8��|��I�_bJ?�Ii�FEך��3h���=x���}I/E3��S"�9o���~�t��������E\o�r�D{�Q���C�����\>֫���E�("\�����V��&hn�;��p0�����a��f':�d����W�L��z�CF ��N� Y%WBa�P�x���2k���&��<X5C�b��8'�L��xve�Ȓ���fό�)ئ��y�����g���&o�9v˟g�(a�Y�$����Sc�0+j�s�M���L�Y����iQ7��~R�
��Ȉ࿩�(D[�.;\|.�0zD�u����}��XW.46�S����)%
���Y�@�����:�WC1��q��+sI���E�b�Y�F��u�+@A��\�FO�&J���Vq��(2�3�������)���<cRfp���|z�i�H7�����\(b�V ���$ˢL��e``rr��2�iT��ُ��Mo�q�'
��O%�S@�<��=fFǛ�����}�Џ���l�d-'Ϻ[�N���;R'j?[�=hF�L:��h�
�v�?� �%�X�	2�Gd<����ٷ�{q�/Jd��U>޴xYq@����A��݇�
����Q	�EF�)�M�낚"�����R'O0�KA���#SU!Y��G��ȹ���w?�l���_�}�R��p��/*H���_b�*�����9�gk���L�B��˫��(_R�����l��݇�""g`��&<��د X��AkP���z�����w��ෂ��;�/{?�N������g�}f_~�_��
Q�������]g����k���>3���*To���`� ���������:+��cM}��k���G7�����*�������a����ٻb���@���S���nQ�ԓ��,�S} ���it� K���i��f���GI�c�!�߇/��{"�L��f��k=-�B�6ê��=$��}Pq��_^\�+�Z�o�g����u�d7(���qS����g\������z0�$�2;F�� K�ϊ�9��_'tq��6�pj�k�Ι޲��;������_~��c�h���7��.������gM��E&�qe9sͩ�$3U��i���<30���5���s�ݘ,��v}�ʮe��=و��_p1�����ģp�"
\F�L���
䎃(��ߌ�}0�`l�P@0
�A�Bʃ�!2�R�R�GU/�\>=�l� z{����.����X�a�H�����&���Z��?"�R<�.�  .��;�$�i!�׫�WP���GF'���M>����(Dl0)aI�Q
O=h(��yݼ��E�	�.{�[8��:�y��=�'JP���7�l�m��+�t�,��;��atmʍ\����Y������"������:o���e�ۿ�����s\��$QFR{�OԊ��@��ԌP���=�v>�|hH"p2��ų��6E���`�>�g�&��g'�\�\�ԗU��|1o$=9 �󹟅\¤ՕekR�:S{�C��8D����1)��qb�GF0�����ի�w�>�8�0�<�v�%�Qs3��&Wdj��^�HC�XS$ZX�%��h!���O���ۜ�^{�S�.��mR�é�_�/:Bɴ�ԀU���Lz?�뮋����$��[dƊ�nd����{qߣm5�%*b��T�|`��V�\k�J;����UO�Ea�v��Ing�|ꎻ�R�lĝek��0=kkO���w�@g8�A��:��Ӥ��S�t<�26"�ڣk�5� c~�w��x _�g����52x	Ze��ڎS$�ޛ�"j�p ��k��},��YQ��Yʼƾ��Ђ�yź�[�b]\����L�`��������=_���苅��Rezru��)��cuΑ�]�!�_/ao͜	�ʃ '٭�$ϔ{mԪ�Xb� ����v;����0�$� cc뤳Qªhr0��B����a�������5w��~� �����E�oms~&�WuG�n/���
z�^��]Rj)��'f��N�A&j���Q�v���{���`��/.�f�������A�
�6��?�{�fl�N��W/�B�{ׇXS�B���������~�_2�vy}a_��U�;���ŕ�z�+2/�j"hq`6xW�wn�@>~�P}�=?��8d��+( �t
}�I���*s��;Llv�z�=�?�>���t���sȩv��nᧂ�o{(z�E�7�C�AV{��s-y�	���[�3g�l(�cѶ�Gf{��8(�S�"������5�'���8���yH[[_��jui�����v~� �l�Q���o��r�Û���x�QN��2��4F�h����J���c�YE����x�»)�E~�־��_����?۷�^�YG��>o�e�nj;�r8-��,�2���/��O|�v�����A8�1���v�~����3r�V̠ ���FG'P���:'.Ħ�A��H�ޅ}�1��Ը��#�>��l%⤿���a��>k�NGQ��T������*�fo�W����b��7i4xLZE�)^�f��G<��:�V�^� �X=k��^��=�q������Qubl�L�_f��-%zElٜ�Yf��Y�I]J���
zQ����[�!����N����?�ę��tB s=~���	�Y��t�׶(���K?2K�[~���L�/���2oƓ���� �*�����"Ŷ�8Ӎ�ԍ�z�9j���|���,ƛ h@���ZjY;�@ȉ��+�0��3�p�Lү'�N��Sú��5�������D9p��}���9\���:��4���托<�.`&��l��G��b1/�y�DA}�gu;E����6'��<Cw���u�uj���v���e�;6�Q�����J�m+b-�Ż�/w��c�׷����@����A����2�|/�h��\�k�,�b��95[�ki�GN�m��wek2�y7 ���lkxo�{�es=z���в��_�u'kj�_cL\�M���:L�nJ`�<;ш((I)�5\��bh �ʻ��cv� �����I�^�Yτ��%��!MV�P'
�ћ�[�Jx��J�R����n���O��Ȅ\UG���}��k:�8�ޔ�>5=�X#V��a��7̄(`�s�@1{�����?��gގJ��7N��,s�!jZKҡL�k��5+?���j�I�I�= V[pa�|�y&�ȶ5
$3r�%'z��@�������ϫ�g�3K�P��Ɏ����\C�4Տ@��3{a�W۶gއT��p�W_"1p��Ძ_:^���e�ΞuRP�z������iL����`[F[ԣ�χ���H�������}w�:�k��o���_}V��3K&�JPڑ�½�����fd��h`=������F�Z��qQ��$&�S�|��j��5�3w�G�����?@gU�+W�t;@�h�Zy?4�J�;(�۽S�����0���vF`{�s��:'֘�˘���!�d�,��O����\�z�=d�w+W4�����^/���՗��⊦P^W������W���B(WQ�;�q]+� !�!6�� �ȋ;�֡D� ��*�{�w'�e�hA��i�f��>���A����
���������ۿ���������;������,(]��٢V$���wo�ǚu�V��^�=��1wp"���p��i��_���9�#��P�� ����<���M�yƶ@��� �C�H�s�����1�����CʊBNǬz%D��q?Qͯ��ۂ�}V����=�_]N���p]^<s��ںぜ���`j\O�;U��R�Q�#2Pj��cN�������)^}����0z��$f?xp�{�O�N��p #� �����L]��\�Q��*\���c�!]:m�1��kS1q�5-�U,� "i�|��lY���Xe���+���o��@�lC+�c|���e�����'{UW,�Z�ՅF�lv�S���[�1ڙ�����65���:f��*]S��� ҵ^`�>�Y�Hk"91�E24�Xc,�:�r��v�����Τ~1�-J�`1;�9��a�#�dН�L�|v ��3藓�+[����4۩��g9T���s���4��X8�9vk�� �/��N϶�}���SN_T:[�t���]�(����C*��/lu��H���@sR�M�ۜ���u^#@� �y���.z�]�:Π�f��� �b�'?r"�פ({g���8/�ח��f��[����縈��!�,����5�I_G]���;g�����7���2HW�ѷ�qD.B��t͡@e�ܗ)���U�!�]���lSb�ND̢EMl���G9*3"��t��?��;�gǎ*�Т�l�H#�k��E�ۀ���^�~EV�mvՙE���>d���Çw�����c�-���ō�W������X��Շ��X���f��ғӐ���TÞ7Ɩ'NV��U5=�.%�i�×�}�y3W�s ۅ�K�q�ݙ<���5�>F��U2��}�*�\mΘM��ϛ��u��b�T7�@s�@�a]X\���X,��C��v=�X��᪔O�3"y�V\���!D�gk�+��@8;Ә���m?�����i�6J�{��n�Qwg������ �;[k�F�ώi'mofz�p�
w�X��1�k>����c�E�]������v�L�+f��-E= �{���m�x՟ @���>�+���v��f{;/uȹ��`��>oV����L����>�/��$G���7�{9���|\��Q�
`��@�'�W$���}G=&2�����e}����X�e'�$�������J��A�Yf4����Y��4#�N�8 f�B�ΕŁ*W�*CA��ݽ�������������e���?���7��%�[q]:��^��4S��2Y�xv�=��vD�g�������8g�.扟��a����<$s�`rQ����{	Oj��!J>�Sԫ�k�"��.�*V�F�8)d�IԎ�}3�`S�$�qh�{>�O>PB�]ls��뻧� ����a��zP<�?չ|d�_��c5��Z�,���u:���EFZ��R���N46o�� {�T��G�5"|{D/C���u����|m��Q�ByEF�0�V��hݰX?K�5�{q�e��.����'�C�2.C�i���&
�Ǻ��3��n�����?�Ϝ��c�u��s��=t�[�������)�~�G��H(�G�#SS%Au�9�@����a�{�y`��r�UA����C�p�`�����Y�C���@�x����ί�75@��Jd�"��xhqK[V>�a.��q�Y>'�H�s7�	U���e��@��M��`��.���rI�.Ϭ�g��@�&�c1_� a���)��7�ש��7qMq�KV=|9����|�ӬkP����SW�	K���u˪9�Y�y�m�Kr/��9�W\�%3h����y:�O-��PI�۵D���[����Ѱ;ʅ���9H�e泼�����s(�����}��PQA:./��;o3
@d}�I��A	~��ft�rd��^ԛj�F�9��Sqg_�=)(No����fMY��'��}�M�k�ּ�
���� XN���1̚���~d�3��=��9��~�R�)��#�)���������T\�Tc'cB%����O��������s�Q./\cR~?N!���6L�=�jc�dE-%��7�E4�l}�0Ł�Ȣϙu4�Y��~Q3g^�Z�G���3L��>6���S{�g�/.o��]��%��Ա�?U��+����{�O͞��|��x 0[}�����^R�+� i����9�$��р����,?輞���̙�ԩ�6ADn���!SAR�p>���2��%�Z�2�Ǳ�-(��|
�l	�j��Y����H�p�h��5V=X<�� C���z˺��>�\u�G��d�Ba`�><>خ� '��9j�����lE�==�")����x$XIQ�}���F�B?����z�{{x�<� a�~b
J�	��]���=�W�����tm�� i�/hAQ�������K���3���!�S���5�(���)��\�N$	_h:zm@�+X�8��ar�+-Ξ�H�����M��6Ӣ�=���7]�TD�9�������h���=G*
�y�޾�����KFj6�s�d�wh�(��$o5���4R8U�S(~4Q-\�$�^�+��O�-�x�ɅJ8�ij ���XD�c�YּB|�8L�����NŎ9oI��M ���?K���+�<� 9�ڔq�`�+�̰w	 o��N8��$Qm-�b���:��?#��h�v����BO�Q�=���l7[J�tS����
��T��۠^)|C��]����ٓ����GI�����%F�/��*��rNt5��=���Sݔ��/�<h`(�D.�:X��%xa��Ҏ�K�=������9s��=Za
5�\����)px���;��0S!�d�,	�=�XƼ֊~^k�ז�D�+��?7�*��&]8���&HZ᪆Kw�e���C�/\��zcV�Y3��U�t/3��nam�`WJx��M�C�n��KG:z��iX�u(��e���.w"��Z�Y�8$���z��̼"J;T#Ki���z��� Y�e��z����0��ay`��} �O_����	���T}�gw�Rs�5�8�׍rЯE*.�wm��.�����7ާ���7���Ӟt�pee�P��]����LkQ"2)]�͞���g.ʁA|A grbT�E6,Q�N�1j]�b]�5�(QS$����T��Ia`ռ��5c��n�y�"�~�ژt"����rb蜪���j ��k�uEhU�Jk��w�� �w�<���|��,���Q0�ΐ-?�o�Ν6:�A�4�}$2���QY�Qv�裸���N���m�F��ʷ��$=��$(��bN�A;d���#p�h�a� ������(�pzo���:t+2k:"�Śܺ��`��	<)��Z/8�I������G���ƃi�m��y 32��������>�5X�Q�(�Pԛ���
���R�R�A��� 06#?'K�)+�K-8]X3�3�WU�=��#�z�I��B0�51c�,��)j��U���慿?]�M�);�59/o^U�p`m�9R�����u��{��u�Ի�YW�$��W�P_�D:�<�hS$r�� �������}T��z�S�{��j&�eɡ)�W�����f�si_�&*����+؄��{���l���t^�Bo���>�'�{��/_���[mW�K�]FO{���d���E6�:�)ؖm���k�����5N"c�2�R?F��N�A-�&���1�@�*(s���=xבŅW8���F��B)԰����S��d��#yy����q��8�+�s'�'@�+|�|�%��^�ʽ����3����_�utA���
��z��	�p6>��X)���3���,wa������ɳ�%�Ea� �5�
p�0N�b�Ա^M+�����fC�;��v�.��X*`�J�ս�'ݏ=
�\ُ�YE��d�mS(~^�U�5�#Vb�E�,�p�?!2��ak���G�#l�0<P��,��bć��Ϊ�~{�fФ�Nk�̂���I�PQ�?ԁ����O�"ÌR���f��ƿ��
�6X\��Ц�W�T�W��fd�G$�|N����K�|�ǯ�^������s����l�"���ұ�X&>��6
q!�kZ��^�R�N	���I�y�:��u�8�4��yu^܏�i���sĪ��;�s�9w�J�69o_�R_$3ϣ��G2���� MIuɮ*8����bo��k��H���?��>�I�v;��=�V���O��v�]]���Ņ6`��aw���r��̲	�B�^%��~�H�bP�f��q��A�N�䄗��\2�4���rJ�o�'K��>��������֐�n�`W�%���{�5��cp��=}�����>z�G�>��%�O�$��s׹|��~��kfQ�O�m��9�y�J��izH6�oE�T\������
�bo�ͨ�������e�67u��C�#3�̻y�"�����9��6쳻�e���Aj�@�����1�{^��\x��mg_;PK�ց�������J���j��=:�IT���pۅ��(JQ�W��xv�xY�+Y~����x���;Ԩz���%�X�,vI����	�Ȭ���|p�9g�ؐ�3�ѷҲ���	�B�}��+^��)��Rd�����n3H�z�C��9���8� Ӹ�����,"�C/��A	[��??GˀȨ�#|��E��R⡀� q=e�;��@ .�꾋D<��y�.��ѷ��7Pt�-J����9�{lԟ��6���$�#>o̓׏�����U"Ö�9F�!0'BI��l�>Q_;����?<�+�m�((�Z��<�ֵRp9��@�s�&q?�/��΀��ԘE�((RgBGzk��+�  lWa�T�����ϒrb0�M�|��Y�����h��>FN���{���P��h
�:%���� &���ɶ%IɷS�ω�����|�sh{��7o�l���û���\��߼����K��Wv~u�o��a�Y��#���q��`2�+���� �����;�*#��5x Dx 0AB���� `�����.�l%DH�T��A�����L�#�}� |2�ճ&�] kO0�H!�����Mj� <{���+.��p\u=�\�8Ӑ%B�s���ת���#87noo���ZMB�߇�����G
k��*�=�Y�>�<�^��d7��^��dAT�
EM��l<@ k%+ ;���]�\��׸����j� eP�0�R��l���20pۅ�ڊ���3W�Zh�z2�L��0;����{�ߔ�iwG�-h��`'A����R���z9g����43�u��]%��ĝ�������{$��ם:@ 3ws�f׮��4>>)��E~^3k/�}�zswK����U�]þ�si���"W�ȐcERqB��S�ր��X��)�Ĉ�lA�e��TG�M�$Tt�A��ψ(��lmo�6��B^w�#�C��Z���\{�8�r�}�w0��5_%�����ꅄ���Gl��a��v'_I|��U�-wl�G͉ӍD�r��1�*�瘍JFG�k��ёMΑ�������+8�$��1��a�У'�P�	q�ЯCVuS��dC��9�3�Λ���l�f���y�)��w�����>�V3e�A)֐Ȼ]uWܠq�#�Ri[��	�|�z�E--�$M�،5F%8�����8R@�F��9qGm�����Kɟ��p��Iiڼ�	W����z�;Ъ�H�T)��~���~�r%Id�R��S��Fם��׾~_û�;����sPT���1*�������v�}pM�-���ޓ?��+u��hD(WM��σH�̢}^܎�o�6=Ԑ�}g�g����Ժ�򛮓�L\�J�t��
�Šy6R���ƥD8\��YO���=��i&P벚�ޫ��iLhg7�t�*�gi���iSf����X��F8}���S��ӓ>��2j�����i�s }Q\�� ����-*��Ɠf��my�dl��r�9��J���^]�N��zM�â3YD��S�����^��b����N:�©8	�V ����Z��c��=Ef��Pկ/�S_
ԓ��T����K`�>uD�7��<&�Z t������P�L�LL��h����AP��TIj75H'��5�5bd9z��HURҌ���K���e*k�V�%R��9�iMN��A"2��\Ey�*3���=
u���\Y	��ɴ1��@adT���N�+�_Mo�j'�`��@��0��0Vʍ=�d��|�^[��z���ݽK�u��@m�!dM�j��2K�=ِ��{\?x�O�Ni�z�z�
X��.ҹhm�S�����ZdR�y���8�+��AK�T�>����ͻd�QG�xft_��Ԓ�t�ƪ�F������х\��=�8�?�ȧO'r��CJ����f�( Y軶Zh�YG6�ǅfƣf����	�G�p��\����l�lN��v����d|nkg�6�6
 �J�m��"p���A��`S M	Z��xuA P����Ņf�a�H��x�Tؘ.^`d\�{�e�a0���p <Ȧ޼yC���H�:mp��Ji���\��������?�@nks�b���R8d�{���t&��{:���(�em��@}K��Y�7A�3n���|� b����;$����ܥ���hʍ���D��叜��t�Ol�̒���e�X�3���_ӓS⒨jr��,-l�7������f���ށ!2����2����3YaLo,l�ٲQ�W��� ����42U{�4���Q��q�L�D��V��4�kQ�X<�4�u���aV�rҐծX�fX�h����*Zm�Z�X��i���cS@�����iA��>�v��ǿ;�4��D4*I4�2���s�[Y�'Z�c#�%�c�q���*��3O�3��y�"ԠR=" j�Ⱦ@䶳�/��}0��	#��|/��<����첕�i�//��R6h;cP�����f������t��&􀞔/x�Z�gDG�P�� 'uEY{���������7F�a�k��0ҿP�^X�t�F�f��A��RP����������]�A�����B�T�2��I
k�P��@�H�e���?��i��'~~��z�Pޗ|�8�^S&嘵ND�Iu��A��A�Z�Sm����a�s�>�f'[[�M�����$g{nS�����^l��z��i$�l�MD���؜r�����OY,�=�JG1{�ʓ�k,�?χ�	�X޾sH���\޽{+?������F�&�N�f:t=Î�?˽������r��>�G����9x�����r>e6�?�{�$c 4�<�q{�ƅ1��o��~��=y��!�1�]�J�����\]\�Pd�& �އ����Ǐ�x���)�����OK�.6����و�2ӟ��M�4��={�]���E?�R��i�>���J=�T�E4Z� �� T��l�=E����1�6��W�������|�NJ��#�?}ѩj�Q�}s�-���H�m�M���H�s��S��0�T(�HU�
�� �J�ä�6c:��w8��f�:s�����Z�@BT�+�G�88���ck�4�T��ߺ�(l
�馊C ��/�R,t�OFdhh���������,���P�VyNjR<�+��Ȃ������]\j��[��h4n$����`�O�{�t&Gt`?}�Ox6^C�y"�x#἖��ͷ{�ƱO�f�t5H�<@�����&3)���b	�A@�IZ�9��6L��2���!C�σ��;�k�����t)��3ZxN��l�>1C	ьYC=��`�jG)�`�,��N���mn*5@G�#΋��ҳ����(�{-��*}&�.��d���y�]*������V���Q#��3�R	u����R��\�����Z@Ń�eu=`X�'&�"b�"#s�������f�kn4����'hH���6%�D���+BF��P�U\��kE����N�6���Q���F��;����J/F�0�R����~�t�M����"ϑ��˼�*Y�������V_�<��qH�-Op|�]�=� ���d����;�c�-Ua�-Qb�3�H�:�pζ:&�7BΑ��^��rO��MT%H����I��}.j*�*9y��\��iGV���y�S)⑗ꄔ������w�g[���gqG�(j(Y�G���`q���t�f���Qu7G`����� �@���5+��T��"}�U�B���%���mC�A�,8fX����NT>���X�qՖy�̚��_��m�wNy�0��l�.�K:8���"���X����Yν��{{K�"�����#Z�F���A�	���yCRud�7.�N��Tӑ:�6(Ѯ�C�.VCQT�R�(�L� �H����W��U�Qv�~@�"�we=�q�-�W��ip�k�v�b������#x������Lyj�,��9��4���n���wC���r�'ĭ_�p�15��h�О�zf��.�uS�(��5V�����|�z�ra=iJ�~ ݹ�����x�|�,D��i�p}}��і�W�����Cy��K����|����;�9��+}����)k}e
bq-j~O������sw����\I�������-:�P`�?�^e���d��Ų3p�f�p�*�~�&��?����}`��V����:����Ȁ��������?�;��U�ļQ	�<�N��ҐX�Uiu�$k���� f1�Ĭ���7웲�e��X�q�e ���������XƩ�&Yn���>��N�cF��O���A~��<���Fv6�x�x�^9F�)$4��8��y��ky��{��D7�Pקc#����m��N�-d��N6o�٤���ӧ#^���#x��sfn�g���yT/]�;�sO�箲�2g&�7p
����a�.�<٠c{yy�V/}�5��Q����n��hFnG;��>=�绷��ux��޼~ÞR�YOA�����N���t�,A^S]��6����aW�Uq�W*6Z3�w�+�cz���0.ю�  _��ze7�"�J�$�m� ��T3�Y��0*Z��W%i/Ju��N)�tӨ��k�ng
o.��M7��OI�7bCٸ���\=�=�����ܻ��X	5��u��x�V�Q�zL�3�gf��3���l��͇	ֶE�hVM�LwP<$pn 8��'�T�Y^��Z��u�m�u}�i�B��'���������{c�����RTf�W/�o]@�X���U2ap��e5cDf�\��^'�y�PT��@��rU�{��sh�my����-�>�МmO������B&�#�U��� �Keq���r:>��&{�.�T��i���gk7GcW�9j�A��ft�sD���n�u
+�qT���
.DG2�^v�
��X�8J�~W��� ^C��P�ױ�����د����9��:�$-,]��c�a��R"��44tvRg�(��-*�c3�0�f���}���ɛ�-^�{�J;٨��csvzI���r�@��L{S��s��x�do�d�hIZ�*�
��ҋ���U�����UK��Ɋ!��ԟ��ҫ�:�c���4h=�zbA6��M�?]p���?��z��5%�X����{�h�ţ���hP\@@��U�Q��X�=P��Mq�(�Ƽ�5P�/耵�+�;����Bvo�	rƭe�������,+��:��nx�
a`u �'*�2���Q�]��Y��p��HD�J�*Z�r��
%s�;�'_d��Ņ�'�
0J@���x�LמF�s�()��x���'��M��F�+����A�����O�C;�h��8����Rk!�Z����mJhF�Z�{�7liG)ں^�Q*���f�*�H��)R��$V���6<�3��8��@��h{K�Y�o��ƕ��6����Ƞҗ_~)_>�Bnݺ)?��R..����.�����u��R_j5=pZo��>z�ǆ}��i �������3ж�u��}y���p��,��s�_�h\����C�}x��/�c5��`���+9>9��٣Ц���V�� c��pƑ�w�<~�H>{�T�>y�y�㞝�|?��p������w� �f�y���_���|�����\��4Uϣ�#�r�W�|��u��ֳ��Q�d��v4j���֨GY���Xv�wV��c�,@��Wo�(���ʁ;�تCd�K,���qeRĞ�ؘl˃{��ϟ�g�=����,7aJg��{�����2�?��}g�" �o��^^g@0���d0�(�A�|>�����{pW�>}"��O�3�w����:F'''<>��p ��PF�- }�7dp�b08;�����<��'y��c���w�Oک��n�s���7����0�=}��������
��5� ��G�*\���%���P����ٗ���Y����G�3j	L���Һ)qg�݊1��1i�T���ԍ�ң�HT'Xa�2��A4�	 ��3�1�72���ɲbvJ�9��i��M�x[**@K�<��X��Y��/`��"��* �ƁR�`� ��	��\Ԭ"��N�-M�Ȳ
)��x��J�}T���'��E�KP9��}���3߬6T'�T����i]��V!�E�璟W0������_�`��Zh���N��,hmZ��L8�˕�s]�-
 oFk��,�������%k�T,��� ��B�\.�`+^��U�n��}_�l7Pl��O�>+��}��~e5��̧h���nG�R d�`W��S��ڷ�`��E����O��_۫x�Z��a��کl�t�Q�m^c("���h�I��K�+��i�b��|T��@��"g�d,�1q=����lªS-���;d��S�J�`R�,�h�����p�`�{0%W	��{��e;�ғИ΂��z�����HqTN��~M��f��4���p4���E��r@U��i��X���&4#�i�SUw�������'fr��,;�dp���՝�Z��|�T��;�C�ѯ#�����k���w�i���`0��您�j�	�B�zY�:!#�̩6\�k��������I٫J�m�(��"Y�O�ͧ��vGe�>�E]� P*k��O�9��� o��~ٳ�F3������i�eg��dL\�c����fK襢���i=U �}��J12&�R�}��d+�G���M�{��Ō�(k��K6�]�:T��:�lV @⿋;b|������>�~6c�g�T:/z)�*U���q
�����w�&�`N�|�@C�����t��������K��\7~7��R�H)qi��]X;!�ޤD�!��(��@�)s��z_�
ʭW�Ƙ��qas@g��j��~p]���g�jyBI����3U{�Lփ���B��ۑ՞����>���[�R.רO��L,S 't�f:Un���nnl�������𚨆E�5���ϯ(�{�MyD�5i���3��wxx(ϟ� /|I�5�:�x>���y�d�y O���_�: Z��� �N=΃k��+������1h��	��ׯ䇗/	(.f�+��e��?o�>��!�h���{k�j��lѫ��6�U��x0.����|?{�y�O�o=�"�q��1���R淇\%�
���#���oF�{�n���׿�Uԟ�
����g�	����!��c>��s�u���^�̀�-�}tt���*�ìP�����˃�����_��+ �)��>7��a/�}xK�y��I�Ԫ�]�F3�7X秧���s�|�p&/^�$�۟�u���FY���M��'���C�/�5���������yv�d��C���Xr����j 웘��Q"}��]��G�[�~n�y�����^4"�{Ӏ�֞���*��%.�Ԙ���(��OL%��aP���!ZǸ��y��d%�S}"m[�
��>��V�#�K�*�9Gc@Y�4ɉX�(���h=�v�[ �WG�+g�_�
�
G��f�粘_�߫?��&ehз��-U}ԡΜ�@��h���"x~����YeR��d�-җ�6}%��k�����^���t�j]�K�J��G�>K��t��^E� �H��}�������M���'�_T!t������Oe=��K��?mS�M�E9����ދ�a�҈�dƕ������yf�����Bړ�� �����d���� [*)V6�6�"��4�HUF���n���S�)mSԴc����֔d@0ShtJ��
t���h�u�{�ܨ/�݇�aG�NUK,�
q�=�i^����d��~��T4���-��e�VЙp�YCh"q\�Bf�����&?t�|���`�Nű<�h��5-��
R�x�����/=�V���і���	# 85���Vd���u굹��9�$+�/��c�_v��uR���.wj����	��1na8V��0vz�-qg�U%_���-o�Q�}Ț���[{�� 1��4T��` �F҅)����8X]��I�V
�"�Ϛ/�K���eV�	%��8�pN,���d�3 ��8ώ�q��w����s�l�s���{�o�B�/л`����6��z�
��E�;�ܑ����8;� `(�mL�ިA��({�5�8�"�(ASI2\)���"e(���c���K��oR����<�99|������~t����vI��'�c�+'2�Y����}��Ȉv�a��xc��v� k�O
E8F���R=�}e�ӺDˊAc0�7J���B` T@cp><� �Y�]���3U���u�[��Y�s�k��������x4�yd�5��0[:)]�$�`�ͻ6��iT5�b�i15\�tk�W�3�Ԓ=px��ٖ[�������.N���&���/���iV';o��u���@�Ì�����P�.�zJ$�:Ɵ�!y�߾};����<�G����ƺ�y]��k\i�t��&����S�_��q�e���e�����[9���~������5XRk�zS5�3 *�:��J$��Vy�B�]�;�G��g�}ά⣇�2(�%U4��~zN��d KHQQP�kO���΍�w���6Ǟ<y(Ͼ����������\�-H�����9=��P<�h��&�w�v2���o7�ﾗ>0;`՚��4?�;���ٳ���~����G$Wo�J�{����@xf�/	���o�6S�$|](�jw���TrC�����D�-�ؖg�?�@�<�v	J6&9�xC^�˻w�^�1�rX3f�Pt�Я&(�X�5Iv�'m^�An�����"h��A����+h���c2�~�RQ����>��ZfEt�z��`��^�b}��J�VK�(�9�O(��9P2|9��{k��b{�T?�v�o�41��+d�Y���7��Su�� 4X��_�ڦ1c%�`kF[7#�!�54'��̘5�]�gॲ�}���K��&�K��nI�6��8&һ���2y��{D�N�D���b
���.���{ً����/�P0&���,����=��/2z݃��U�*��;K��]S1�m0YͦQ~鈛
%��ɕCZ|�(�0.�Ds��}��
�V����+��Qkt3���npM�᭍��* Q�-2�')�
�WA�U�Q:N�e㊚�
L��xT�}���rYd"�DY��R���������,���|P�<���Xj9���8!�b B���l�ͱF�$p
Y�0ጕf&Ti�m��پ�.���<��yM�'V��@*��w$�c���*�(굷L#�S3N�E��#6���D�k��N��Vʅ�U��f��9�,��I�&���M'���1��j�\Ң�ޔD���c�s�t(w�+(tGRꅭ}��6�ʭ����>Qe�+�ұ��+rM���B`{`��c58}q xw}y�"|�-�	�ɡ�
� �b�кfj��Z��L��T�^նlr;���<D��v��(�
L]&�dac_u���E�}޵�2w�u6�Q�yވ/�)�fg4>L~L�.g�Zd-�^@���"�6��o�|[f��V�{�2A-p�%k��4���;�LClQq�m^�&�Y��Lҵɬ.oW'��}!���P1�9ԕ&��F*x%�uN��~��6X��	2?'kҁ��ae�0�g��0y8�k�\�[��[�j�?��Ή���f��Yt	5��^dؔ-+D
�T�/�d{�c8�p����i��2�𫱊�,=��� 4`ĦJ6����MS�����ԧj[sP�x�M�9�m���=H#f�Ԓ[�:� �B{� �J	�z�J�� I #_=�Z>z$�nP����f���t�(P���Ͼ������9��2':2� ��;(zf�'_��7/yЖf�=������
`�3��g��fJ��57 ;�#�y�ɢc�P����C\�e{{�G�dg+;�4�Kfj����� ��H�
�x"}(���\j�b_��)�J�j��;���W_?�/��L�>��Y,��M�iv�?f`���ʿ3�sfl��U}`tL8�2�}����`�~>�|.�Vn��ވ��b� )�D���� �-����i"�A�w�Y���e/�п��*k��uw������W_1��~7���b���}�'�.�����.�&�A��c���Rt�Ț*�	5rcwGv�o䱈rzr.�["{��g������<~p(Of��4��lO~�����6�i:�j�Y>��9�0�ex��~��<��<�s�A����ڇX�́L�������|.�8���@oϿ��X� 2+	�*}۶�h[z�D
�Dzp�ِX��j�j�����r?K�D ���N_.l�E�L��! b��P1`��X�4S��KW�*�^��{�g�aW��C��(	�)
1��!Uz,3d�.��E-����sX�CQ�
��H� �X��+���l����� ��Q��ƕ�,WyU��b8���cpӶ�o��{H��\�#:X�9�,�,�Y��og�FyNc��[��!����gqڵ���-? Y�M����֟�cn�.��.�3��T�ه^z��Xo��>Ҥ�����3!�ꗤX�/��4���=��}Uꔬut�ǚ���(25�#(��.�'��z4ꓩ`��.\�5F�퇕���8(�Q��1��ۜ�m�a���&�=P�"9�~3i�����i�D�)���>�2qb`|e4إ��t�꧳���֋�Hǹ�֜n�3�)T�*��Q2B�Uq�����C�|�E�~Gc�M�����[)��m�t���ڱD���ѵ��/�F�iz�R��͐����B��綊�i�ȵ�W&eE�k�$���4���Ru�ʵX�"���4�x(Z��J�,���y�[`	-W������R�
�$��Z�r��,�gݛ�SjV�`ײh��7�ȸ�;�,"��𢶋�
?�+99�b����	#�0�І���B$�������-G����ƨ�R�v��F0Cc�I#F:�qv�V��`���6ø�N#w�4����!|��!�@Cx��^a8�g���z6?ro;�P���u}]ZA������]gu(�O���.�~��*t���|X{����)�^��}Xd�}�������,�`��:lI3Y&P�"g�cQBIV,��Y�`�~
����!C���)o��d�������21[3ך,��*��?�7�7 =�\����&|�����X�>XF��{Uʹ>7T�R�ad�2��{�3;(���ǽ ����N�<}���M���Ņ}:b�U������0�;��*��_�fd{�  92&����K��_^P���"�%P�A�Ǐ�7���|���O!��|҆Ľ��ӧ����C���OD�Q��`�8��+F�lb�Ԓ��N��J�r�3���Ylg�Һ��(ͨ�����Y��o�ٳ�����[~�r>�sj¯�-Qm�l�v6�m��T:������~+_}��uky��� P�l@�v��^���J+Eu���g0Z����&��[72��0�����7��.��J��`��<}�(��ۼ��R�V�)M�} �������[�/ "Ag-e������,������{9=>����ٿ�#7ol�V6� ��ڿ�A��y~gК�p�I���H9�qX6p�������B��nȃ;��g����;��:���<ov�d;�avV�&��=ʫ;j�9�>���ץ�IQ�ThEl]:�̳d��fw-8��٩
����aO:qX/�
��ig^ۈ`5^X�4�B���cR��T��lt��N���{��͠G��A��3p�
|}rZ�։��=�������\���6�����q��?8��m���M�@�h����31��02��fH�v�l���A�����=!&S
���;e�h�
�D�<P?G[0��βC}��΃1�,h�NJvQ�A>���Gh�{���ձ�YA/e�@k4@�R=�y�����pK�tY}Vl|TޞY�N��XY�@O�1�v����w�T�hͼT)u��SkB�id��T�Õ({�7�Z���.|�g]��d	�^�m�,�@-��j(�D���P��$��7�]DN�2��	��6�+΅``}p
vĶ$�<`W��y-�����T#�-�:i�.ț�L%+�c3��,�F�b��|@gi�+*u�+L�W��Q~�JF����a]��w�|!}6���B׼9��y�����G��	7j����C�%f�
���Ct�~�![��lI'a��e���B��FT4��A4:<p8�@��R��y��)O�!�	�jM��Q��:p����Quy]�%����Uc�)���;dҳY�q��A�E~F��iT���7�L/��ی��� �?c����� s�h��	�%F�V}�J����%�-��R��� �ǉ����,~��1��]^GY ,f#:@Y@�%}�
�	Ȏ�,�l���d�;��K�ʶd�?M�P��LfJg���5ht(�8�e
���B���GT��
<������$�X������;�:9�D��+f����UKe����:���@��E�I�J@PqB�Jw����.x�uE<~?�s��!�$*�_{��&M�<�,c:V[��v��"A�ja �^��!¨k4�$W���&��R�zk�$�[�+Tݩgs�{[�ݣS;�Ц�}7��&�����>�=�u�-���� ($��t���Qv�w�3��[%Sp��=��N�훇r;�����dA@ �Mv�x.dhCTDG�y=�����d[���ݝ-m<�:����w7��;/��e��ѣ����SJ����t�%��e�R.ON���{y��޿�>[X�����)�g[����;w9� V Z��i���eA��Ç��ݛW�مE�	���'���N���$�����V��zV����[~�ŋ�ى�H������1n����Y~Z���_��C��{v/���#��?�t`�ػc��|B���l)���3e�^��gh�`\��d̓'��ɿ��o䷿�F�?�����ee�[ڛX��*�gt�"���ʄ�0Ǿ����??�����싇 �Π2���ͯ�ܺX�G�FK�Jfq�)2�q/&�]�Q?�?2U���z"7�3��hd��?<�N�Rv��ѝ[r� ����F`hA��j޳0}vճ6w��y�����ܘ�4c����}q��I�֦�����[�ӟ�,���������<��������� ��2�0�n>��ގܿ����<�^���	�2���}�L|F���|�y=�wO�̀�~��6�e͐?;�����������I"�wq9�zűQ�z}b�d�F���>�8���J#�ԗ�#j}Wb�l�2hy���<��Q�\��R�U���mp갈"�S)�Zt&u�{�@:�y��S���l�<�s����J�VdqzF1���΋Q�����g�g���إ)7*����-E��a|9�&��� ���v*�Nk��/FIbm��F�+S.�8�
k8
�D�xos-B��/�(��lŽhɀ��db�A�B���f�g�VRĜJ Dt���]K(�˛�������i�B��论������L1�T�ĝ��AlfU�.Z7�8 w��+�T�� D��f�@+�T��h����FF�gQ��j��I��� �%<�e6UNP�TTj��W0�`�CW iǾx*� ���DH�q�QT��.����p�4�7O�F�?d�1��L����X���h��������/�	�O�Y�9Z��/}\ג�,���X]Y$��ٷi�i�6~2L'��<��\|q��)�/�d����#+uA?�?ȧ�O�Dn�h�
|��0k��Ǽy����>eM;�p����а@���|h_6ϴ�!�k��q�;9
 �Ψ�	��Q��}Q�X�jG^�_�_[J6����9����k�yK�{>��6�>jQ#TX:�ť�r�g<R�� ��z��� 3������璋q�amS�ƭv^7����sFz���{skJ�(M��Ĩ���9��;�e#yz6��Ѝ��U�̫��S�K���"�p�K��=�A��MJ�o�`�J����Ͽ���'[>�D85b��65ji�'���<��sN���f�<�d��i�0I���u�5���R�h��ֲJ�>O��'��^[BZtk���Lv.�C��8�E]y� ���jc]�pE�mQ�^�(%284!�*V�M�88H�@��t�&�l3҈����trz��[��5�F��b�pc���2q�̞;]L�n2�i���\CJucʯIk���T6�M5�8�_�[cM��Z��R�Gɛ7��L������xܾ��E+m{co��M��legwJ�C6��4־U���궿�Js,%���H�~������W������߽z��A��-*�u�HV�1�d���0�P���\�..9��N,x��i�����Ap�k�掍ʻ%KT]r;��}*#>|����h�n��h�q6Q�5��n� -�i��uR�1d�ng���7��~�+����r�ޝ���S�r���Qu����J ȚN�L%��y���
��7�ܿG���� x���)���`�����dJ���-�c��&��xL���4ḇ�"�����&�|�)�����^������ǿ������\+�}_"�;�����62O��B�ֵ�,�f�{��� 5�RǴ/3Ć��wz2��_�y1�2πYmÕN{�`hwx���fm�^e�O���u�L>�ź��A�tFV�\d�������LSmT�^>:��Pe@���qr�^��vU����B�Z�F�[[9=���W���K%\��T�:l1�?\uLגIceT�3j�g�8�A��X0j��K�ic�B�LZ��BJ�#8�\����k�yW��;����^h�_2ۆXv�_UѰ贈~�ձ�h�ө�l��MtFhl���ӟfԁœ$��Z<��2+��	�(w��C�R2��Y��(
�G-��}��:��۸����%1�E�ߛ�]�T�	�&��dĩ���3A<S�������NI���P�6F����S�̬cӉ�`���{�b�\!+��~���CT:g�^e�I�Ϸ���X곂��#�d��g޼N:��&��֝uFꍪ'�5��A�D��{h��D#���0Ң��(�{y���
��t�7n���#r��驔2�6G�\Y9mY ��4�v�x�`��:Ǥ +��q�x?v�!��H��\����������k�
���ʹ���]�ۢ��b�?���(��?#���t:('!�o���7��ߣ� k�d�`���FQ�:�ԛ������$b;��"���/�È���آN/Z���R�\�3����rE��ټ������.��Ů؜Z۫"�,nLY�C��rQW����מa��*fgm: ��Z�Ð��3b�����j"D��|���yCl��2��i�y�O��n�ײqz���d0k}J�>`���Jd��5�L���5��Ն�`B�@ ����{g��}�^I|��_2�B�M��n}Z�+p !CΎ��0�g(�uK�����iTQ�y
�C���L\H�a��x9��1) 0kL���T�"�G���ߔ7���1U��<M��K��&R��:El������c���Լ�@Ë��Q�N��Qp -��j>�>V�WU���5Z;ecUGK��f�aB
(���T�U�">����^~|�R޾y��=�I%|����n�f��&��޼�����x{k�Y�����zA�S���H��^5(��Ea6�q/����d�]�/��:�ݥ��_|&_}���7Q�h����*�/_�@J�<�d.�Z��V��U�Ng�n2����}��9vwU�0���[���1�ha''��%�S~?h���1h��v�r�i��kC�dvw'���#�����O\��j.����gL��<����٬��|/Gr�����'��Za���lm��ֶ6N�蓵�¨��5�%ʿ�����3־N#k ��P�T��Gݗ����<�� z`q�!#��DE0ae,!����j���A?��w�D�3�0�g����z���ָ�6�M1����.�e����h���4T��@�5�Ȅ�=�Y�b��N�髕�j����F���j����E2���˾�L�����{c5����L�jW������`����t��vH��*d��SomĲlb�%s2�nL��)x��F���B�}6�G��mִ*Rd�m�*űU�c�`?Y�o�J��Y��@�[,��>Q�-jB}��l�,VU6)��0_�Ӡ��`�)7g�ޕާ5;/G{��w�G�H9�m��,��{M��%$�g�ւ��C�=hP�<oSdf?3���g�� � ����P�W�d:6�h�؈�-"��y�6���)��H�����d�L����D?:�2n�sZ����}R�#9���J������H0�@�6*��/���>��� k)-���ځc7����J�֣�E��?[m�]t�F������D6��?|��
�����r��=������/G�G H�X�Rr��}���<���$�?����a��O|��v}&e�9���_$� �7#��cY�~������4��U(|U��J#5d�l��=����U;W�!���ΊyWL�'K�:����x^�KW�!��){�QJ-_py���*�l(�7*YW�}C$=�"�H67Z�/8Dٿa�rx�C1ώ��lN��uu���K|��H�	�fӘ2��R��h*�����@�>0*�o��y��W�o���,�'qL��R�jx&�K��e9X{Z_d5vA�v����(7c�S�o9��T0�Y�`�����˽�:=t�P5�0Xc�>?����P�uWX[���h�5�G<`��_\w�P���y{�u��FD���Ԙ�n:׌Ak����_�w���&�o��V!��P.UҸmd=(x����lӐR��y�&��)�hE�
(��슎=������GA<c+��˛W/�ӧw2�8Q�\��KU��� ��8�z0�)��Ca��N�������BU`�,Y]�g�����/�˷�k������ρb"�6M~6��}y����2�ٺ}X;�f �g��#���"�SQ J��X�r����f��N�-�PNev�nɗ�>������_=�`�f���I����e/�������� �o�s�3�LH0 �(��ҊE� ǐ�&�(*�5g��]f���轼�����~̠�2�ϊ�7oܒ�[7��M4�����nI;=�W�Y2�pz�o�䟟�1���?|���'��I���Rr@.�J�iW�o��3��o���w�*?3�%����rxx��W뀢\\������ë�L{�a�Ч��߱v�[)�S�	UF "�;�Щ��í�����16n�ٱ~�`���=�g��������~�A�d$,YHy?$U�40�EĲ�V��`���f%%�F�H���3�'S�L�����q>���# z��MhH�GcdV֢F�-;T������P0�A������L,��B�=Z77w�� ɢ���`��m��a���?�PX���ߤ_�� � ���F��"�Fc6L ��T�X�:�������Z�S��0s�I4E"{ ������vڞ��U�es���^�~X��櫕7����${������)��x��t�,4�A�^��ۦ�s7$���bAW�9;tc`A��q�_���x���XXCF��g�jE��W�S�"x&�O����jiU(���O�����'�l�zG�����{U�2�>�q~�� )��~�j�����	�6���U�߾:f���`���+�(��R��A����AB�!�w �j;�MO���Sf��^�DE3���>�rx~ [;�Lꂞ�}-�&4��D�gt� ���8-D� I�Dί�mJy���|�U���Pr�6���ǯ��}��\855r��3��G�5��Yīj=yCg]Ӓ}�B���1]��'��K+��(���|1�r!)���$��kؓ�J�,�A�ΰ���C���LF����J)��7������� ���Dc�FyQ���l��oKz����V
w���z?�����X����Q����� A�?K�C~�	3��6ӇC� � ��Cko
v���jwI^I�,�96�/��k�*?��'��jR9�^�^t4��v���"oH��ʽ�z��с�_^o@�'��Ɠ��X��� N�q� ���A|���^�FtU;
�m�%.sb(����>����������4��r~.�� "�QPbzߐ,�(��2EF-�9�1�q�󝞝�Q]Z��dQS8����Vw���	���(?�����9ڜ�s譹��s(�a��ơ�H:b�޳��"��~8h�n�P���*�x�u�Hͺ�:�w���w�}+��7�\]�Q�F�Ҹ����ev�Ƿ��y%=���3a�tr��Q�eW�`D�"�ޯ
�5��-� �|��3��?�Z~��o��g������G����������?���������Gy�g] �:2&�4�������=��]����}rE@y������༐?��O�t�{�A�O.i�N����2�ܒ����� }��q{K���
�s��l���J�/��5�d r�Z�	Ơ��9s��������{���_�<=^c:����	�Uwz� ���{��-�f��&IU-��� �؁ �&x ��Yl��
� [Ԙm�����.�����3@�� ve�d���c��m�͚���,�%�OC���	�Xy4�^\���:�g�/�зՎ�����k-� kGn�m�>swg*wH/�2'�4���g��Eg4���l��쉷i�i�#u�g��o+
t���:����
@�c�܄�
}�.��:>9��sN�L��בuͤ�T	T�����:��>����a�n������ݯ�F�@�R���UB��)[�g�\�|=Q����Wn_lߏ��j�
~i���֖�b꩔�x�ӳ>�z�!���@����BA��;�E�_�p����x?(;�\��w�>���S�=��rO���"���=mdJ��t1��6��U�ۯ5��M�h,���O6�늽C�x�6od�6M���K{��9hK*����:-���O+2�ln��f��x�@Z���<IRd�QVU�A��hא��
��G�L����U�t�L��������@A��qs����ZN&��D=7�
����*�sNJ84h���EF��<jǷ���H<
n�H�XH3�W�uͱ3��$>�l���'���sӊ]r:T�t]w {{�AU�j�D��~p,kչ�҄���"(�f�z�	,�W^S�)�`�5*�h�Vtj{C�d1�A��6�-�k�����,���wVݩ��nY�CК+�G��pI��M�P��hf)97�IRJfP!u|���Y� ��(���aCɫ���A�bI�B�i�S8k�VQ�y`��H�:}���R��}]�off������o��qM'���񨘏u�]i}�i@y�c���^��0�wȀ��sp�wf�ϻ���5Xޜ��o��ں0��@������%I�
��|B)5{xz�u-�B�S�nb�`�V:Ȳ�SX�$�lEg�,����s��f�t�-
b�G��z�~I�Dw����XS�)����x�g	���\TjG��t���gk���M~^�_גjqG��ی��&�J�ц���<?�p���SF�ji���5�=鐈���C���?�x)���GE�V#�����E>�9����٦��_f:�HbD�d"���mFy 0�����zV���³��d���1<d	�?�~N�؞�˗/ٯN�_�]�ٜ ���B� %����{oo[�����~#�������}��N:���\]t�������o�&��=�ͫפ���'�0Jo��l>+myv��x�B��yD�Bd��ϕN�15��׿|�L��z�VJ�^%�ɓӣ����6e�������;�(}��tkd%�y�w����b�/�[��&��D3��F�!��O�(zc,���޽{O���{�!��9<?���9�:�����N3x<�c�rWZ�
\4��{`&ZR	&�Z��Џ��c���&S��zG�/j�nޔ�y\�I���,�{`LlL[ʼ�Ή�:�7���sآ���fO:y��l's���#��`��n����Bwdk��;[r��}y���L ؉�Ŋ�Akx�4 ��0jI��ޡ&��վ� }7�^�T8l$���������S�������Y>�+����	�ǳ����0�f�uv��w�Ko>��ι�w�X7;����+Ɗ�j��gY֔<��켚캇�Օ�&�]�f�����"Q���#��4j�0g�ۖ��|�e�Υx�q��z�T���LiP�e(�b��6�;�&��`�����ߠ�]��7��(N������J�}�{b(cP��v����޳]����~�{g�R�H0��|6����ݔM��`'X3p�=�|���AC�	��EP\/G)��,��[K��`e)�`���8p��9����X
�x�p'��Մ��I�`ۛ���:h��<�� E/ΐ}�
$��h���S*�!����R��^6H����^����)`�͖��?��.`�/�\���ȫ����J׮��βW2�d;� ,��� ���P���W~)�̀kVïΩf���ڕ_w��	w�ڍD{�>0�ל�'C�L�S�*��j�������,��JC�e�HD\%��~�n\��N�V�*r����,�1��.���Բʛ�ղ�Ӌ��R6��0�DdP�(��YKF(�RW����Y%�\aA�BRg�U�T��4��_��_��=��_מ�������0���j?�A�����U��FҪ@���ʱ8�s����n__$b]����x�OA~�΋���6���ߪE-���B���g{âƻQ�J:覟�q^fu-���`�K�G��ˮ�t}��}fwу��ɑ @D6)�>�k���S;�Y�37tZ��|J�V8�[����`#�-���On�#������5z\!�/�Di[�<��uqq���NUb��lRj�q�A%���
t��k��S��6��ϑ,MP 	dެ�-�P�h�)
)\�v r��C��P��ۃ�#��f�3�_����/�YU�)��Q���)�wo�j��T!:W<c?� \*�r�x���>h���Md��fbo�������w`�J<���9��}��������� ���������ٱ}����цt�ޖ'���6XqF������Si�~�=E�h����#y�����C��],��� &�zPl�4{ur��](�n��Ǉ� .�BDk�S��Sy�b#��]��q��AF��Ҭ�ݻ��嗟e[|����Y��>�\���Wrx��Y^���������O��\��3cV����'*�5��[��q��7���kXr/A$�Ld��l1��<w��q�o��������"FP ͠��ݼ�zb��@�ʂ�{K�38q����b�:�+���bEZsG�i�Op*�5�A?�<~7v�2��'��k	7is��C�u��(yT נ5f[]����ZCƮ88���u�5�>��tP޼���E3˼�,3ŃP�G�sg=>c�'����n�����[[	���L(��^�2����os��Z�d���.>�������̫%1�uS��IUᴳ�����p_�pݎ���p�s��������ʱ֨��[�+N�L<�|.���d|J�T���r�漐��mn�<��Dcq�$~����pz���րT}i��=�Wk�S�]�O*�Y ��~c��4h&��-�a����0w��1�Hz�����N-v��W�Ƃ<�E����f9�(�Տ�������_�4{}~&�B��Qp�ф"��ڀ���F��e���涱�˱vfG����Q�_A���3y����F�A7���M98̆JƦ~r�b����/�~8I<�m������FdெP帍n�A��pz�#���ԫ�m5�%���]��A$��k��`<��Y2�>���I��P�H��Ah1���|�v87R)�^���F�s���ǲ��څ�����C2Z#�D6�l�7��BrU�o�),��R�[�*>"�JI�(�ދJ�Z�b�Tj�t��<H6��s=���|���3�򳏭Ƴ7�0[��y<�ދg�}TW:c,�D���@��/2�,�@�`v�L�$�_!��c�v<)�>{`-kX_��k���:7�AK�y�P����٘p!*��̻>��V�V����g!�2��΋�3��-���3k���?x�I<t�@��j������ pƴ�&��f�us?���<���x��Q?˲e.��E�@�78�0�����������6���BF�mlӳ,9��T)��Eo��M���>i/&�A��_S^�f�p��y�!�od�y�@	��ʮ9��1 V>�֤������X�Z�1�8��;����F�5k~Ȝ�ϼG��ڳQ:|�x���8��C����A��կ����=&���*� ϫ�Mu|�J���o�o$�y��`�3���[��;hCL=������(��ȇwǬ�A]�7�>|��0 �:'d.�6jG[�a 
R�hҚ}fT0aL��ޒ����W���|�p��{��*r��<ᠫ�);�Qnܐ/�|�����e�-<�_�2�ܡ� 3)��>F�b>y�(��O������˗?1�Ց*�򙣗ם;����G�s�>aN�N�����>��)�2����2��x��&���O� lǨ���9��kC @뿣�;��ew��|eP�R@�jGX3S���B���wDA�a�� ԏG�O������ɶm��9���ؐ�� [��ӏ���W�".e?5�zg�t���6͊��tX�e�Ʌ�$�ڹ�.��h�D��0� %?��� IG���ꀬ���<�!�tv*����5k9����F��V��&�mkO�X��IWUM��Ve�V=IJ2���ZP���]Ջ�VU�F˔_W�CF�|_���z��L��|�i�����{��5eQ$�XT���\������g���o���_[��;���?�8�7�ɕ��:K��g �3^��_�y�*R9C�����L�k��0��|�ξ*e�SqFH)�1A4�g>u�I��~Ncj��7�E���hݺ��XKٽ�2X�"��/o�΃��ĩA���N��d ˢe�l���W*�+�\Qf�0'�\����6t|F��+
_�x�R�/�����dmo�f#�}Yv�&�Y�z%���T���9��Mu��� ��rox�E0��0�o��;�o�M/����V ��8��AF��+x���0�}k]��7:�k�Ɠ�}v�`�ѾNW�8R���cW��4�M�,(wv<��c.����F����.U��E�-�:��^r��3A�
p��`9�L��dY,=o_��w� 7f��4T��>�C���H����io�-�%~�O�0���9�.p�jFNA���k0���(}N�����H�*�)Tc=������?Կ_�szm�Z�3��Ɂ��\,�A2�@��!��,:���)�O�o�T.��-^����)Ew�`'�s� ��x��ѼA1�A�F���̲u����z�
T6���(�&!�����ӳc�\�"X�Q�'3�R(��&d:p-�`}G��w�P�� g��S:]t�)0SIs�qmYH��u��b�s����)ݎc��V��{u�*�!%��|�[[�t	�Z!�#��H�Z�v�pW�*ม�X��N��^6���y7c�7�~�
��<f��ƪ���?�(.�]��������l�h�n��jW��7�]W�������}���xL��1�Oy����QM��-��׿|/?>Eq����AM;`,Aq7N4�F��5�7�����[r�����=�bg�H\APj���N�圠k���Mپ���}{,���ݭ�G"�(�h�߸5�#��Ŧ���ѯ;����s�'G'&ݾ���6�փڐ�ĚP�{�!������H>e�u.s��jTH�;D���%h<Gdif�W�됭�)떑%��Z�:�@q7�c�ַh��L2 ږ�h�"*��*Aj��@~��@a�X�i`�z �	Z��D�Q��-��?��,������ ͢��p����d���k�f�-������֢(`/dG�p��咪���UK�~\��w�µ�ǥ���j�����ȥΑ�g|p��U����Mj ��R�Q�>����GF��,��o�d�uʤR��5Xtd d��k-ڸ�Wp�V�c����i�ޙ�LpchOt;L���z�IHp���	�o��O%�C�~�]����~���%)ͭ�n�@���o�~�D�(x���b���� �5�Gח>����%����
jpc���P�|N�g�D*5Tb���% V	��M���oS]������V�	+~�Ʊ6Y������YfC�9�7C�U�lES�ғ+�^�� W����ٙ|:ji������Ǣj=z������a+�:>�
p��O4��ju$�(��$^K4,�)����#��.��V�[�|S�m�����/II{�z�6��s��g�V���)/;��z�^��>,�5e��Ҥ�Hna�����n_xV�Hl��Lr�E�޴X���׺~�H�@1j��t"V���oG�����΢�	��hV˜�:��gG͸���{�������Е�������w3���Gm�S8x��)(�9�w�v6W}n��#?�NF���f����C��o���N3��P����J��l�E��79k\��?v���#��U��9p`Ll�C�d�sI��u�G{<uTi[���&�hH+��I�Yj�Ud~��f�@����,Rl����k�0>i��R�(ܲ���M�ǛL6dv1�H�G�|�����Q_��\á�H2Y�����J���c�.3&� G-֧O�
�u���:��`�X  5��4uް��Hq��ʘ4�ųg�wP���<f���gg�:�5�fC���]�A�Mg�f�^���N-����}t�6i���{ਝR�QJq��8Á�D�t8�/'c���Z���ͻ��*����s
/	VѼ��.%���3!�1�`d��5Jb�+ؼA[�5c��೾!� &}���:���^dZ��ۓg�z"_}�+�{�����A[	i?����i�U=�s�[�7�JR������.� >�u��J7z!^SdM'����9m�ك�ٺW��Q� ֠{X�"u�\�Ub] ����12غ�e`�&֋j����&�UD��X�(� �,�olI+�a`+�m�:6 5�;�P>����F�.��xfbD@+|V�z1)gF�*�Ɔ�ޛ7����{��B�#N���Z���*�b 
-˼��0HYl��[k�ZNF���c�
�4C�e��L���q~�`���^1x������F^���p��,�ӥ�ה�FC��@�I}�������k�epK+*�����~&�E_��b�N*"��� [�$�u�[- W��ưB`���={�O�2��^9��[�&��t�+�"�o��{1��@��K�����9oBWKL��鍢f����&�=���v\s���\
Ļ�ߛ9vP��!�]c@*X�'�R*"d �>n	���cr@˰�hR��3����()^��91؊�W(���0YJ�#:��e����E��a��6�&
ؒ��ܿ/��==��!tQ,m�̧��Z���<����7j��	���H{�`c[q�@��]УӠ�xj[��l�=sv,���x�M�Јt��L�i���P��&7[���$���]S?����S��u>= wL h ��r��>����jE'�c�5F��J��8�^��-�m$����:�,��ل]�
~BwQh�*ZR��S)Ύe���q�Qs6}��\]���f@[t�$y3I���[��=v�4V}�x�
�,6Q2*_R�Ůb�L���$ϐe���u�D�Y-	�;��N}�c��0PVC� ��j@����2$���c�u0k�Cj,
�_Y��O)YԵ�DZA�l:QJІ�ui�{��=�Xё�0�S~N5����A���9����*곪��b�m:迕�e������a���Y�wֳW:U�"(��N��3ZЌ��'~�X�!�`�6U�0�X;�ؤ�W��F;w��b�t2�1��&҂&cu<ZspA������qvL.�b��\ �e�0�3�1ƭQu�V���N�_�E�)8ډ��x��";|�N���ֶ�0e'����W�<r����<�su��[]���O��4�}lJ�7�􂪱�ç�
�����;��������l�;��l�n�De��0:���+"�cU��;�a�x�@qbm��U]�r��O��1��W����ȸ�>�*��O'�rt
y�|�<��ɦ:͘)�9a���Alj�R�)�46�ƺ�lƍGRm�R�qڟJ�e2�š�Sg΅�\p���lj�y^A�t.g�P�[2[1"s},o߽��?�Q���ȋ�e�T�y7��e�c|�H�j�Vj1wOZi��:mx\�Ɩ���_���&z��6�:3dR@��S=n4h�
ٙ������O��|��ײ��-[S�sT�Z*��$?��:�y�6v�����k��֤ab�j�5V쭦�琈f����\v"	�^��v��`L~��U��ʓ����Y�	c8� �g'r�8�U��>fI5�`:���f>�v�)�z��g��찮La2��6�U�)_�N��Uܔ㋕|�\���!�Ӎd.S�GxM2�����^���^c*{�l+�ў}���Po�ގ���Y�E�,ӭ�rc�nYw28�);y}x�Q�9�Lr��"��-����h֨3t�h#q�R�L �d�O�1���eG�ӌ�v�q�"�
u��<O���X����[����޼�$��ɇOy�����8iI���
�`?���֣:�O��G�� 	Yױջ,;����F�l�@�`� ,����C�c��ڂ.���N���1����<��\Sg2d�T׼xus��s�U�ϾQ\;_��g4���2�b��^R��8z�� �ac��.����, �-RV��NW�]�Ml�����3IqLz�&��
8)l�4�՛�H	7dj{���K6)������w)M��Y���P�GU�0��0ꊗJ�\�Շ,�
�ҽ��4�z�b-�0�Ea�=�u&���W�󒑸:�֑����!�E�����@G+��
:pR��"6*���0T��5�@�0�bA7DK�{e�X���EA��R��M�����'�EA	IZ4�PUU���S�O�/	Q���^�;�Z�|�Z��>8w΃y ����QY��Q��u_�Ή��$�wYu��Y33�ڣ��]/b��4�Ty���� b͆8��r�,�U`*V}�D5������t�E><J��B54gðK�q*���\���W��h�0X��)EWnp��G*�C���1MuD�A
�[�b��<|��;J1>����{�אb��R6>�2`f��_�}+R� �و��1j�}�Ѫ�|*1�`�r��N��P��:>U���N����N�v��cfhd���d���ى������w���+f�A ��Ӿ�+x&W�6kv�`�Խ.//X�tttDYe|���!�g�����p�t���[�BA�@�{�x]�>z�X�3�Z��'��A�bo��Yv��׋J��!�^����	�"�(f�@^��!�pm�8�P�p�P�;=�G�[�]:>�uh#����Q@��=H�B��9}T�4ꪵ[@���5ٸ͵�B4��t{y�o��e�q=c*�Ig����������Ў�H�E#��oH��5��3w����w��%Q�Hx���;Lf�1��� �T���f����������~��޽{O���B�Ы�9b��ꡪnM�{�����Ճy�\I��L�o�FUI1y/�ླྀ��A �x��)m0p0x��1D'j�������_�ϟ?���b�=![P~1��L�7�}�{��jJ�`��5$�KM1�����;����X�$Tp}}�^�x��A��y^G�&�D/�?��8�]a�� ��㡞K�0U(1�TY;'�"� Y�	�b0����]Y���m���)��Fja��^�O���g�����^�Q�� ���d3s �Ƹ��K?�����!�P�O�кDc*���^�)�Ǻ��Z��f+5���q�h�~�R4�2k�yc5 ��p8�5r��o��wx���Ƞ�b �2�Z=D��@F+9�X�!��wmmE<���G�R���[<�0����g���3k9`�c�|�y�|0�`z�z%�D�� ��IC� � BU����Γ�S��N�ѧͭ+�UGI*@L/��;V�z]�F�8Z��__?��@1)�Q��\��ͪ�g�EnE�8Q܁�zYgJ}��=(�7\��1IaJU�4�����G���f�.s���	.�C�%��EݻMl������0����j��
�=X�h77�{�����%6.�:x.@R̾FW�N�2a0ư�׿Q��)v4IޢVj�����ܸƧ��V��Z�V	+��깄��* G�:�-���٩m]��{��>M���l�T� �S�gܖ�	3�U&P!�Z�E� ���K�iv�i���<��k����R�޴���o*ס�{]������2��V@�1��T��:}>,.;:���q[,fW��k6�ny�:���p�#�!�_�S���J���֊�ߵm��yRӿn�uЗ�NV;\�m��i{����k�ƙ
�U�E�$�F���L8���S��d?Ɖ��}���I���O��Y���:?lRۨ��,1�!��&�kH�ZB���Y�`�7�۫W����%	�J�I�.X����¡�.��Wc	���N�����+��$<����I��P�PPy@C�67hqa�&�s�}�&C>C9;c���T�g���uGR�P��4�R�V�-��q�$���XMg�^	�mzbE��VY'g6	o1��u*rl]�N��̆���INT�i
�W��bkgqx���VJ`�2Z�oa�Q2��b0+�s�K�����R�۽�#����h{{�A�(�5�IAޓ�l	Яܰ�Z�`q�V�N���C��\�i��ت�pdx3�_��ts}��#z��	��ܠ�̼�P̓�bk{�~��?�?�`����]��f�����ڍ�A��\� $��+kkg�� ���4T��������;����)M��^=����$T��/�ҧO#)? ����.2 _Za������ɑx�&#!D�r�ҙꊶ"A��e�sŠ�@�
����y �@�g#�tzr��%��r��5�U�l����g�z�4�
� �A^���"rv���1����wp���� �Y�cO�?^j�2����p��!x���%��B��=�OCIf�i�RZ�ݱG&�}qvI�<g0���5����|�>|@s�t�2j�����zfP�l�Q���S�2�³է�%����ޙ�`��� ِ�}�|�w�F$E�'���֣%\�8p�2ȢHF7�óK���,� ����I��R�J�^��)��:V�_� J��=�O�0�l����`ei0�mJ|>���(���:p�X��@T�����S^[��䷙��L⹯�^��OT��b"tI��)j��пPx�|M�K�t�b�S~�9"Do��&��/����B�#wvؼT~�xLd��E��8�۽`.2O�Ҷu��u�U[||}p�8��m�+M�>'����Z��%���:P�)�,�R����GA,:��r�RwC��ɴ� (����Q��H �Z5��@�آP��wм��I�\�\b���W�_\������{%�{��+>�W�M�!B��`)Ư�YC�_AjF�yԻ��o褈e��}�>2vA�l��������ti1H#�HlC)f���ҘS�Y��.�o��k�hk��G�S��Su�J�[	d}���8���JpH�ɉR_��l�^$��,T"s^�M���\�M�[�;Ԃ3��3P�kkA1�z�����,�i��3�DS&bm
���ZR���Ja��x�hLMӵ+@����k�����}a�zWm��!au����(�T�CĬ�\5�o����}���E� PZ�Z�6[����UJQ�=Yh��iB�"���� `�(x
��|E(7bG�Xc���l����#d�*��UE78E��4�4�:1�3%%ؐ�	ؓ�v��4V����R�DA�P>5�G����dx��+�y�xʒ)�`�re̕d��(��ʺ�Q�D����eZZZ�'@5�xz��ɻ���6mm}a����#�T���U� x�$!)"�p`�
�X�\���Z�Tv�D��͵ZN�k���{�����"=|t����ݿOs�<�W�:��y�������_��w���-uܰ��N�Ί0<	f��לIn�Q�x*NN䃬jkk��יx�����ۼIc�,�\��YQ���ٹyڼ�R7����x}� ���X<Y�zG��[W^˳&
C��AM��.bԉk�bJ�y���J�&5� ���XJ����D����9�}�����H<Z�~� pO�L�#�c�4���	�B��=~jF��7����!�0�Z����,-,��<��e�0������0��:Q�ԭ�|�b�S��M���`$k�� ��k�%ʩx������c^������I�`o��i�^`��5�aT�hz6�vF#����¬�N޾u�n�ِ�@�����!�o�lB�"�UB㯐�6�3�0�`y޼��zi����Y�P�l��\��(R�� Zų"�)�K���#2dD�
c���T�"j��s`�o4}�s��*+ʴ��v�Q^�뇏L�Y_��Z?b,�Ē�W}BdfM���� $�gC�>���O���.�Ja��+R
�vctҩCq-���[��PgoS֋�c�3�QÂ13	G�*��$]N��0$�� \��[���<Y����d�|�t��p���
B\u�i݊����PP%a��NV�Z�jټ��*����sO,8�k�θ:�S��O7��,۬��U����0(�R:��z�+j��➫0�K� Y�Zw���+i�h��ʰ�[�$�����i���r~7o�ԦtX�|��{>�p��4i���`�C��k��QhBtpD�'>��`V�F: ��@JJ�)I�tg��:u��#	��`���w������Y�XK2�Әc�	�߾ %�N��޵k�w�k=)�*F�챾��X����t/kʹ��S�0,��� -˼R����BF�����W�2�֓Z͸��^�1t�6�p���w|�P��B��J
�{2�܀|?Vfu����K�bLɫ�(� (�����0@���ͻ*9S	�������Fk�=����봱�!,f(�~q~&
���x��z֓V�#y=clhYص(�M�B��L�1��1�yP�{$ ^����x� �� �P�Đ+��f��������r*�\;���9µ/��x�1ә�`₩�V����>�I*��=%�|*�U�	Ӊ�NFa-�P�`s�2���*SD��zMP�tR� ��XO�B�) ���6���]�FG(� �[��Z�ho_	�_՚; '�����W}3)�E��o���B����LYVZ����|yc�67��ɓ����}���I7nܐ�N�W�Y�W�Wdv���O��0�8:<+�xF� �M��
R��<f�r�wA{�҇"�XQ�����3)p,�3�����s~8��<<���97��':nq��d`|�A� X�f�uյ�Dе!�=m_��i�X��F����r0!C����	�<h�!g0?���O���/���6��S��揲�up x�r�y�_�s;��` ��D[/Z~@C?��?�Έ�7��V�fiuy�V&�<�7��=0���l��0xL�U�]?�:r Q爂�˫t/��;0���|�@KM�/۟ū7b0���L�ˋt���`_d�BeW�`l{z�8[�Y�K+t��=z��>ݺuC���p_B�GR<��|.���٠��Hv���!�U��l�D;\+3<��WE�},����V��svir�]�?|�u��m��W�?��������8�<�~�*��v���O��S��_v�����X�Ik�GQ�9�R��:c��	+J��+��8|,�w(��N��5]������眃�F:*>��(a�Q�LdmUY��f��y��R��*0�-@r��g��:{�\׳ڳ���ʣ?<<P�:�����v����J�`ls}�R7V�Ea	��Bӓʕ�>�:.m���|:;����r�kH Y������C�bHl9"J���k�H$t6c:�-�M��s��U��s}�܌�t���[(��M� ?"u����	+�u.�����B&CZdY��b^�cF킫x3��aŊ�-i�%�G,@��E��6EH�>~yÐ�τUj���@#f&r`ꗍ9_+oP�N�%���o'A�/ �}#�E��hT��
(���i���ן��E�-�3$�&�C
�6V�Պ�,������è,oIR�@���$1�S�z���ȐI����f)!��0W�ڴ��~�뎒���I�Q���z�����	�)rK@���'��[�����Z���V�Ч�V�$�}Y2�㇨$n��Hd���d6&�?kt��fYQ;�x����{WF� e�0 42�gH'�lj�K���q�0��KEf��n	�_8�d��V�k�u�cr Ԯb�w8�a�$Ӧ��� TxI�	 o��c~�ٳrp��������(kǪ�5�	����!�U�&�d�'�'� ����'d]e98^�dm�����k�,xvr!
4r�@'~zv!�A!�����G�,Z�Z�.���KC/��*�bg	�S��P ؗ5�"�<��w�.��/���P�#������1���9��O[���kz��Kz�a��PȘ���ãs��1}�ڥ_{O�Y �YR��AX߾yG?|�����x�P`� �Q��2���ݓ�����K�{�m��SaFm���:�c�}�a ��xp�E�ų���"-.-p�����le�!%@ ��y��x���<w7�ރ{t��m�Ɯ�+ɹ<��_vh���c��*�z_o`��6heq������]:�wZ�A�ph9J�!c�_P�
����	5����r��:?7ī%��ܒO��mq�Hu]�C��o�/`5!x�
�5��&c!�3�&� C�RBኁ�;_��ѥ�g�cõz)d��i�2���,�k���Ѓ��ie�S��X���MC���D�Y!+$���v[��[<&+n�9�Q+�>���-/Q�+Oi�� ��JBYҗ�]I����Vr�n�ZtSh��u���mM�q4�Q;1�&�ycJ���6�1ۀ(��#�W�����l�I5��s�rIo���`�RA�B�p�B#$H��r/iȯ'r/��ε�</�dd����񔜨Ƣ�Ҝ�:1�c���o�gko҃C�Et�)�����J�׊��S��1Z凬qrH�ʮ׺���W�s/Y##�f��Z�Δ[l`Ӓ�lC��J�uU51o��cYuUi`S���2��dr(������{�b�	n5��t�nʠ$��ֆ����+�y��
	�8I.M_�v�]䱸�]/��j�ʶ�t�������Em?sX���o���&�+F�,�.�q4�cP����%*�����,.c��n��m����L�)�2�bl�Q��e|�}%_"�>v�X]{��;��!��T ���V��.��&�������p��Fi?���)����i"_y��{���<G�d��c
�Z*d7AXC��5���~4^K��Z�H�����z�z��%Uܳ��nߦM�?P�?��dx���؂b EH([U|��h0�b�~7�yD��B��=ɽ ��,_seYko�P��d�Z���6:S�Y�D�"�D�B����3 bQ��,�Fb �=亀�\�jMFl�(�wߏJ��!|��ˠ�� ��}u��H \�b4��'�
I���4
��',�P<}�z�׼k�K:����
�K���>����A�u���֌zH��M���T�V&��~yG��s)xN��A�!DN��(&,/FñP|W�!]k��&ҐA�ʝ+
�b�2�,���1�Q��HH+�_��uemE�ó���g�x=(�$W�DG߂���/�˯?Kn���a.�b�IES��ޥ�_�����Yl L���	Ŗ�0��S��P/��7�k@��� �L @&r�旤�����Ȟ�5���h��cR�\0�s����j�/4~�(C���� kDc~�g� �{x�6�ޢ���&��7��M�/J��g����yF8ܓ������&����m��柳����s������%O��g^����ݻw����vC
�{!	YS�Cm5�t�x��r��S��F�o�^���2����P�o&�X]������ ���P�Ë��"l ��C=fv[���<J��(��9��3C�f(�Sa�k�D��t��f�:�}���L��u?Dv���Op}�L� ����'����w]���M�x-^{1�-׭JV_��uAoE�\F��̖gE �����"+�T��t���z�yL�_��
��古�_�-�Ϫ�;�F%�z�cwJ���r}��c`ˣ�,������>'f�2�㡅��[���x�<W�ۚQ�SM��r=K���d �|r�Z���U.P09VQ��3���R $�(��
B(�L�)��'^@Lc�f!1� k!-��P�A�\+JJh��|����19C`���-����N�b�'�3��-W�]�1�~W�ɬ�Y��+�ff�`R3ML9�1m0{��v+CZ�iZ�Qw�%�i�RQ*��l���ڕ��T�ƅ~Hc\���M�v��_z����8c�?ߧuKFa�s�$߮l�;x��Zt�oI6z�t�Zu���7��2�����}�+���Xx�-RL�N`LΔ:Y�Ca�)]����&!G
QmgI�j%��0)�'�S!ԣ��o�I������E+S���:�W}-\�CVaȀ��,7)$P��*���=5���H^|0�[9�l�x�͑q���N�0$�i��I�V�5՗0CX_'R�B<1 ���Os<���(���湨�C���[�E1��Aqqq&�S��o���X�D���{u��MڸuK h�%7����s�r��8�׎�@ѝ	ZWkF��P��G#��(�G����X@Tk,�Q���X���X�`S��J��75�@å���
@_h�t�}�"D*螖#VP��Z�2V���Me�5�c�so)�)o
����7�J��n$�Pjy]�
�,�?3��[�ſ?��!�p��g���6Ä˧hL�5yq�N^��Q3F��M�6�F��S��0���7�
���=~�>}Bw�n2���:�,�!�i�޾�@/_�L/���-����:V@ ��F����z��� �3��o�~���=��>����R(��{��>��ѓS��ՕV��4�6j-Ó�c^���kV��o�)$��]�`�.,.���"��<����hH�18V&D��łY���Դ��@kyu�A�����v�@#�4hz\��� B��k���=���c�{{�V�fy�����6}�ޢ�鈆լ��D��"æ&;gy�n�/�\=�wn��'O���ZY]U��kߓ�=��@7Yh|��۞N!�M[����JX��s��x��h��J����:�8����T�� X �"l�2�0ɒ��ȏD=K�@O4lZ��0:����ʦ)��g-BQ��h��)۠l�=5�G-��J޶ɝ6{*�K�!ev��B���t w��Ώ��ĮW^�Y��-�E���'�s4'��*V�u<r�vij��)�� �0�ۧ�dp��o{��s���3EI]�p͘i���W(�E�L0c\���;>�A���!�n�R��`��������Y�nh_z!�G=����tڔtք����z���v�W��r�MgB��a{�p���<Wmn�Fdh<��N���<
��C����Z��2Q�}�`����à��zu���rn���Dz@)�R0eOw��Z�q�	k�K6�>��`W�<�����V��D��]�Ok���>���l�g:��_6��^�I��eDz��㺰���۽�Q:�qᒇ���*D`����,&�틉����i�����	�Wy��k7m���k��]�����a6�5�_���De����N�b'�{���ӂ�'������sa�Io�{�6c���u W�-��% �s�J`�!z�0%5I*���A��Y�>�˴M$��ļ��5��Cn��UV���S�E3�;D��$��R���wK��^�g	���Q0Ƞ�\%J>0�Q��S+�[����gl���~��u��])N
�����#�$�w�i�.�Mȵ�w�.ݻwO�lct��"$�#����kE�+�B�P6�]��nN����ũ����x�dG��!�0 ��F�Ov� ܨ�p�(9i})d|�
��X�nz�r��fG���6 ;0ƴhD"�~��1�7�5�7dz]�B�hgE��KI�譬H��^�~�(� ꙝ��������Z\���E��ب�t*�4�=��[�)kn��N�s���(�ijE.[}��)�h!�d�w6��/��O�?��%�nǁ����w��痯��}x��œ�����Ȓ�� !���sɻ���@r�1Cqe�"@�Tk{�e�F�ޗ�:�Ik���V��~Q���(�wzzB��r'9DM���M%�%g^��Z]]��e��B������I����\g%`i~���<r�Ԙ���?'��=�����������ڸu��M�ok<�}�,ޭe~o0Sk��,|x�}n�H9�gXwY_��g�����t�mlޥ��5��UoM4�Dy􇤼fP�s��,�C�\Eυqf4O	A�����D���,	y���w�j&"� ��� ?{SY�/�D8��T��v.x͜�sa�'�`�������Zu:���ju�c��i�Q���r@Io/�#�LI�>?�����Ͽ~$������JgjG ��y��L�vM���#�R�}�dvү�TJm�z�:~��Y&W�\C,k7\�$w��*�Yy����w�/8v�����������xק��X!����h�-e���`]0������[�V�a8���h��Y�_�(�e$ZA�_��n�^��!����V�*��Ҳ�σE1�q�,T�����%՚ɓ�j��'OJ|Q�G�ݐ��9ޔ���V�=1�S�n�%m���&�]KLnz�g#���~�<J�9|�|L�b�C�P66QI1�g�Ww7��]�Ғ�����<���s[�n^<���Ụou��y�}�M\zc���EKO!I ��.�� "��*� ��{�Μ\�-dE'�=�B�Q����PܴmId�p����	��b�a�� T���1�]
�ot8^��å\�}U&��O������{rt��[�H���Bk+�_1��[ĳ]nb_�F��{�y�*7�~�%I�BY�Y�F�p�������z��?�kȜ��DQ��DŘ~/&/�*@���&(!P*�vV ��Z[]��>99��D�+ZBA��1�nnn��G�����ρ�yX�Al�\���ma}CQQ(���N���2���E����,_?1���7�C5��F-T�����Zkd)ZO�(Z������Nd!hnՄ�>��P�kZ��J@g�2A���^�0&`�X�jZ�I��^8�SW�����h$\����s�LUL���B�.���͜�G���V�oJ�W��֞xp��J 	JT"_�U�׶n�,�Q�L!%�j�>�����	!�s<�7��X=�?��;z��sZ__�~vv%����mVo���^���vw����rxNzF�����`�}���Jj�M���r{��|a`pe���djޓJ1�����q�W��Y]�!��7�h�b��3\blY8>9b�-�� DA���=�8c�����7�:��q�H�q�ӺKS����'�f`!����QWq"����8���C�jP���3��L�����eZYEX�'�7J���wf�Kj<?���3�h&j�Q��۷�����{��kfnqE \d�^�98�MWM����ole��-ꑳ/xdQ:��0� 2�GO���*��m�1�,P=�нS)rݫ�t��pB桹�X��>��O��)�5�eLz=3��S�S�s�����'x]���|�x����(&/]���~��<������;�\a�.�Σ�-y�����f6&�ś]��I�2QE�_���J�k��%}�u�N�uGg�w�\�����Ǥ��t
����H�:Sy��������q�RW�E�ϕ@�z�b|�{nKN�q��`��פ�mw<�k�NNza�{v��k���<���>���n�N�>�ZI;����j��<C�`�d��ڗ�Z�TDr�$Y ��pPNm�abz�[b�x�l(�'�E���+q{�`��Dcؕ�#���<_c8��E�#Viz`�"Mx��*<o^�#^��|�^p�.Ql��1�Q�ɖ�Ґ6P�v2�hb�,���C��c8�02`��Ҋy1�G��u�x<�b�����Z$���֠d!M,���6�YJ����i蟬��AZdD,
�J1:�
h�^E׀��|;�#���Ū��RP0���& "{�i1c��u�S�f5V`])��3O�:j�Ap�m���ݕ�\���N�~�C̆3��*��t3�x�B�yT�R���,
-#����b�-D� @�2�����������I�xr�ʇ'dvL}�t��r��t���j�rb�~_�ǘ�R*��ub�C�I�%o�e��b�����k��W�І��hĲ�,�v�UJ>e�(�A^P:����	IQ���]5 s�a�ZVS�Ղ�}����9���ק۬�F��4/���ʲ*�sttt(�
�"�J��@F��~�����gz��+�G�C�dC��(�!X�@UI�ub� ��W����G���3�����-b5�^��ANɗ��Bn�ۛ�B��ZN�a��z��p.�{�$
*C9�B��(���cZ�2-��A�2xia�Pś�묀�(�������>���<������ǐ���_0(d0���G��9<���1���HΚ���ZE�©�V�~a�H�noH�=���-�桸1r��#.^8=��R���,�n�y�ڶ @���V����7�}��X��s��Oh{���8���K���j�B��5����|�jp%<�i�U�n����RR+Hqn4��"֫�����&=r�=Z�����+�{������˟�& ���T)�͌k�M�9j8�4j��t|)��uF��ynjH��sP�g������@��D�Hi�v��y;�}��U�yk��k���<5߷9�+�5!�l���	��⼑�B��6����t��!}��E����rJ�߅�99�@f�\���9���������<yD�K+Va�Sȭz��myHsKs�{�r���@�&1%ss}XC���Dk��n2*�17#�0�!�Y�������Ȁe˖���,�hum���*�����	j<ѵ<5f�����7����N��o�v��Wyn_)�A_�r��h�޽}C����ayqpr��j�֖nJ�Q�੥��V�>d��d�}����M����1��3��pd�Nin~ 9}j�����b��|���H��z�ɤ��(1��f��{�����>_ 07Lo��`�R��$}&l���+/�MD����W4Q�6�nA!W��8�?��xd�
��o�6�f�g{��Rh+�=Qv��cJ�lU�3�Nٽ�,�on-���֠�~E�Cȃ��H��Iu�)YX�x��o-�>c��w%���`��Fߵ�W���\猺�R��!Z�zݚ��"_zٌ~��MTW�Q��D���l=sE��i�Nߘѷko�*��k�T�zX{�Q	�QO�4���*��Rv�ZcF����P�k1�Z�j����,�<\�7b�������
&J�S�������'���P,�	L�~�
���".�v��L��:�4lE7~IMN�R�ʰ����a$�A��&�cZ��FU�=�n,���",���cR��Qp�m��'o���翩�>�+O���S<ܥ�-E�Y=��:�oZ�y澚��z�QH�<��|�u摼	�B�<D0	|���3�>�
��t��U��C--�%�K4�aג���V�C�6��r\0v�e�x��!l�Vw����ϒ/#���Ж�Mc�B!�z�<�)�]�Y��0|E'���!k��!�zJ�вd@ ����p(fB|����nӚ#ۏ�*hcZ�B�G�atސ��⍺s玄by���~{��Xy��CΗ�=0޿�^�xA/���6n�����<�K���G������������	�8�q��q#q�Ԡ/
��bܺt����hJ4d$	�ތ� ��!d���������������?�;�����}�}[i��E����i�5�(*3�s?�Gp��^7�Q��<�ux �Ϟ=�y�B����iow_<$ �5�G�M����pC��KI6�3Q�5�P������VV���e���@H���ݗP�_}E���y�d����Hs�:ڕU��ޓ����@�������Uz��>��O����s�o�7<?k���'���_���W���k�.GS�@I�"i^��SDP4���De����f��SO�l�V�`6�p�{�ٯ�o8������e�7��'r � T~Rޯ|�E���L�e��yg�@�W�D}!G 3ߝ�;<�x����=:�;a٠�R;@����y^s������������?��@�̆+�|y� G�@�0���3h��E���=щճ���J\csa=㉢��?��QK��X�W�<��T@/<Y�7p4�c��'���16����UZ3PC2g�^��:���Wx�/�~�����/���W���{�a���a�~��޽+���\���=/do�l���ʹΞ���D�J?�a*��o<��59��ɣ�Ǳ'
z0��>?��G��Z�����o?�|��
T�Wϒ��� ���ſBi�����
­�n��.hC
�����C�]E>�7�Y���rt�7B�ú�+9{˿��aV�zt@�zV	₫V��]ӫ�1�L ��>%�ϗy�(��v_�g!~�H�C��yMW�ڽ~�h@1�4V1U<ه��?����\����	N�N���R8��z���B���Qxj����!���5���ޗP�P�v�D��/�F7���PY(xh��B8��P��+��J�K���Jqgϕ��4�1i���!Zbc,�U�	���n~�@���q�� �����ZSe�Z�w"������-Z7ȕ��3G�/IZ�&� �.%pJ���i��K�������/�BS�N��B~���[�YM����_�e�hG��[���x��yni
d��'���(�=p5�����Q {B�3U��˶-|r6'�Zx��b��7�uM�X8Ut�l�A:��-�dg���F��� յ�}��^h$"�b�e�l�(LbZ<(1h�_р�C��l`�-.�� %�q�#�er��	��*z������ \�T7��X��P�����e�J2�,$�R�`"����h�� ��B8  ���ڍ5� ��%{��x�@����18�π�ɓ'��K"�@P���6�z���������J)�Z=�I
Sk�3B��@�!��Hd����A�~M�h�4^�ۛ�������?�p�`,����ϴ��B�$��q]_ߐ���L9J4�H�x,������fk$��c�vKx����{��ٳg������ν����K_Ծz��~��:�?��Dܠ(�Q��y��aZ����)��6?��ylVto�P�h�EMw����w���{�<7�D
A�0`�iba�B=,[��`������6
< ���������~��w�'��З��+�~��'�������+������n��h95�G+�	�*�7�\��O�m�ڲ� �����6.���.��Kc��+Z~����K�Ԧ�O�����%��5����B$352~��}b�z���JK˷$��:hϟ<~��
��}�@����]NDO@H���5^��O����'t�ƪ�a�<o��i{�����9� m_�&k~�ԥ���dP�߱H���f֌ 0)-#�e�0�����a����p �����3��tqcͼ̩�Z�D��J�P?0��P�d8 ��]IU�Y&k��Т��{���y{��>}�������D��H���G�����k����>|�=aӃ ��l�΢J2<:A�4\Z=��GVN�ݺ�ѳFΨ8�~��]����e���߲!�\�NJy:V:�)ǌ�6��`�T�+�%K9��1�BT��4ÚWu��eDOzI=���Q�h����;׮���3~��4��������~�b
݋ʁKw���/���׫
��AW��ӡ��L<i�=3`j;�%Y�q=�л|�=��x!�W�F#�+�-j��n�H=�t��b� �AAVsX6exhT��/�b]ʆE��z7�t�q��78�<�wna�f�$�V, +mBmb�Ѷ�F�麳oR�VJ�P��n����� ��k��n�C[�<,�*c9S�n���䥶�ī�P)�~w��"h���!��������k��<��R\ �M	�aj�OwA���1%/A���֋�����NX���=|�HH��R�Ĥ�֑�4��$ ����i91��Qeq�/Ni��H��K.H����ΓGc�ߺ�uA� Tt	aiR q���`)�%��r��u�˘�v��E��3j���5˳¼MJ}5<��ʬ�r��|$����2�J��d:�^�P�3�
�ȇe��{dMY�A��*4���~xX2`�1X@��:+@=1�\^����>+Q�$���
��E�t�8Pam766Ty���� �@Y�HNSCY	�m�����S^n�·�VkU���
��4�7��<��H���;9>��Q������ksk�P%��@�g����я?��>}�@�g'��)�a_Bռ�<^�5�E9�C�� Zb�u��uOj(Cl�z*�\��u��޹Cw���o�Pzs}��Yn�0�!�O���zxQ�9+�������;tqy.
����i:�dR�ȏ��{����V���Gmq��ȭ��ۧ�<������3�� �Lc��A��,?0�H�G���^��[�Aͭ��YB� <�k��F�y~O%������{��$Qҕ1()G4/9yT��K���p������{���������]^Al3X+۬8���5�����7�D�9�0_Q$Z[��*0 ����9?��F�`@���cz���#�s4 |��!zW�'�+j�f��Y6��b��w�B5�4��2Mr;f�]r8\��[����^Al�����DXW�x?���0��K"z�wu��&��gi8��y:�_ļ����=�K�������3���xm.)��gg#��r�c�Ko�~��|�Y R�!�U}� M9�̈އ��m%�	�q Z������S	�D@��1�3�����|R�JP�{>�ܠ��O.�=�J ��*��NS��`՟�\��.s����/b�9�ߓ{A�ݿw��?{NO�<���6���#e�wq����d�b���R�i�-1�~�Qk7d�XKn��L(a�8zvR9Og+%�u7ڒ)׮���m����MQϻ$�]���,��l���{�!���/���܏���;KO���U!���q1X�D}�w
��Q�+|����l�}^<w0�_,��[��C�R�G�6q���u����ǡ���V�vR���N��5�w��q_>��e%e#ՙ�l�sos[�ؿ�o�>D�A�ɍfIi��{]��13l��Z��hG�a�1	�#�E���;j-,�� p Ė��hi���yq���꾴��Lj�T�q��6���[w$q
X��|h��P��X�h�K�7��H��^ڏmZ.T�M�Ap�K�J����@P���3e]�;�yU��u_R!���7���Ȋĵ��"u�:{�������%���N������[f��ŵ�%���$���u	wlӦs�U�\^�g�DZE�\������J,U�� �4��B<}��P���JƏT?�Ș�`	`k�2c�Q�B��M�'�1/�{�wQrÐ?㌟r��<^�%�Ρo�,:x���N@��M-f_��ܤqѨ�b��:~�3�gE�+��K(@z9���v10dN�7�<)�;ɱ�@5�Ǡ���X���S�07��eV���'�����9�1��L\@�Aۛ&�,!Lº7�B��Y���P��4�4���6�$b����FRK�ѐ8�����0xZ�:xt@ ��ht%����F(���g�� �W��_��7�嗟�m�rOI6�����MV�.���H
����
�v0�mn)$��yK�g��Ʃ�T�� ��e����=�����qSI�@ų6��~��W`k�<�T�|�y
زP��B��7��V�k�۫W�tI��7�"���8,�M��&�<�3n2Hø }mf:�=!�P����+"��
�t�a�*R_���� ����J�g���w����*�ٌ,D]������+�<(�����Z陔��-%��F]��A�&(����O������?<���o3��ϳˆ���~�����sgg��}�	������R�� ����H��@Pį��{�����c09��6iyi�����>Ӈ����H�2f��aN�����{�?��"��+t�A!��PVƼ�z֊�!sR�As)x�Ծ|9�������3��u��=>��d�k`v�A���n�ܦ]��5��n;(��l���j�6B>�����𸽗�ĳ�K�8ǚѺj� ���� ���~�Z�iȥ� 7-�}�Rz�Z��<:���yJ�a�K%"���<~�x�r�܀$�vb�f�=�Ԉ0 ˰���E?:<��#
�d���2 o����ѣ��
��\��b}hʅ.P��ə��Y1��mg�{υ)Պ�#�r�����[ �敵mqp�aV��*���BL��"��=f
�$���V���BD��t�\�3����R0׍B�RWꯛk�w����g�Oe��ۉ�O�b���}�S���H(�)����GLzZ�Qa�@�Z�}�Yߕ���қ�(1�f"����G<�˟�:�}(�1��d�ۭ�!�:?�#F�����J?�0�½�H4\�W2�t�I:�şN�]�X84�ٕ�$p`͝�T�IҌ5a��&�)��T  `�5m��m>�b�(���b4!Đ�V�F��'
��%�]Đ��`h(1�tWj�:���ܨ��b��O��y4	��.ZT����
��1v@- ʂ��]l��Ut���uW�JH둨�h�̃���;k�W�&���VꃁI�L:���P"�Ћe�W�Gٞ�mK��Xl�h +;Q�����R��6;��T�y�p�bI�j�_K��,\���s�hW`�x +Xج�Qs�y��F�Mdy�.@<L*ʚ��֗��R��ei�)��v(�[���Y\fe{%I�ky�&Z�X��e��v�9Rae�V$��S�� ��[UQ���&�^�7���r8���X�d1�F��\�^%�h�,CF�0\ ��J蘗YiX��F7�V$���dQh�Q�
(���BYxqZl]��$V+ˇ�@+5�>}��B{{{R�
�
jJHw�o@5yM��lo��q��-�9!���v�����[;���� |�aN��H���kW�_��=m0�}�_ʐ�,���P��<���{V�n��[� $k�<h��R)����iK����9i����AaF��f�@]IX٫��q:�����, �>mmӻ�� �aXS\a�	�	Jt1������ B��mEڍ{ë��@tU�%/
k��x��sW�u�@ �H��R�g����%0w���ھ�@Gh���/������Zz���a���6nm���{Q����{���y�4S��4�N�EQE(}-��������Z^]E�t��{��Nք<jl���ӓsǼ&�L˺X��x!GPvG�F1����7��	�B�Nk����77à����
�����_!��B�P�����������CV�?�����G4T����t�J��g�th��R���7b%�:�C(���z���熐� ��X�gy���h��b�G6�B��h5��g`A�X!����#���/������9�7#j�|+��s�K.��m}��@�h��-ޛR(��)Lkw~@�#/ [D���I^)1����@L�l&�W�'>�,���=�I�p㆗("��ٍz�p=�	³�~�E�	a��}}��x��#
�����`d_j�W2=g&��zB�6�꥙���]�����H+�甤���K�Y���v�Z�>���d!J��'��Z���F���1f�!902-#�G� ���=)�N<�z�㋢M����.��o.x?�_2�&���S���hu�{�@>��))~�k��?\!�3I�3�E��^C\r4R9��ʧ��- �@��C�P���!���JA����g哊B��\�Yp8�-U#E.U���|�jL�Pғ<n=������1��	J�
)� C�B�00�'x�L���ޤ9ɮ=�琇��wyeU��/0�I�&JZ�}��=k��3��n[�0y �J��&BY�*'�� ��Ĳ���ү͢a.�`�W��wi��m�u�䐍�v+YuY��^ʿߊ��XsH��N(�w���G�l>s��ro�5��C�­�<���)��6V�4��|K�i�Ew#J�"MkCj��QW�Uބ����<����İ���dAP�L�����_��p��?�wؓ8�2�^x]�Ȉw�A���&`�y�E�8�J�r�F<=�4��%vJ�n�����iO�ѠT��T��\�@[��R8���&�G�u�a_ydx��h�vS���)9��`~��,�	��(�Pk�I��k=݄B!]�Dy���C"|v~��
+%[��~!lY��Cj�pD���&c�sG�)X��-��Y�9TU׭���˖ ]DV����"^q� ������3�����D�ֳ���ua݇��|#���~��޽}+T�Z��/��2	zyak�1���ӧ-	�ڐ�m��Lg�3���/��B��{J"޵9/�g8 1Ȳ/AFYVHONϤ]?�������>}xOǬ��4+vP�^�zM��	mږܲ�w����,^V�gn�P!�
ߠ!G��Ѕ��V�oJ��B���v��~�s���GY��s�A,�^��eo���Å��8�E���aac���4�z�F"�jq��H��Y\��0;���+���QB�*K>mS�W,j�M��Q�`�H~�����	����d�$c����q��rE�� Ъ(��9��r�p�d �sxC��³�s\�j�W����//��u@��C	����x�� kB^�hiX���V�d=yH��<�ᬆ��R��O[_�����R@j6� 4����%���@���-���1X��� 7n,�8,�����2�� ����y�_��D��?�����%��/��� )w�	����ؽ�ޟs4�����<���s4�w��h��-���D)/ ��eO^c 4���S0PJ�sA/�7)�k���?'@O4��06P�x�{j���0V� m�A 3�; �e#�������#� �G�Z�6gr��Ѻ3��x�V�W����d6�Wtuq%��R�OX�ղ(�\�&�%�0U?�=E\�5j;�\�qcbR�]�v!�'OL�(��gu�,��t
�\�.޳3��N�=	)}>7}te��o@���ۮ�;���}z�iJ�l,���U����h�c�B�*� ;�Q�!��7�J����;XV���C�%].�u�B��	�Gՙ~�Rp��� "�������t��S׻��+�j�.f��3/��X�e��z%L�l�4��(X�J�ߙ�Ô�h�Ee*Ҡ�(购|3DMx'��+�$U������5��V@-Uٺ�J��*�����{����?a�{b�c� 0�_�3 c��0#��RKb+,fʹ2*G�kۿ�L
�~C�;������\�����d�g�w��!W����j��!US-Ti �&0X������j�C��sE���hs�p�o��NO\�_]��X�'v���D
y�P	��$L�
�P%p�y��ڕ���`p��z
�P9@N�,J@K=Y!�+��cN��o�}m�;�G�8�ly[��ࢿ6CM ]��
|�&�_rLE���d��D,�:v"TR�}�VԆ���J��
FSY�2%KZi�����ߏ�����`��>����`�	�~9�j���J �ｙ>��a�b��R�D��H}+�	�D�j�������/�� Z7*{�%�/Le}BI��� ���H�i�XC1��)�1:�}&+H�i������q(�g(iPvԲݣ��%��<>�-?���x���%9T��+�� 4y�C����P��h{�3���,^��`S�+�`��Ç�C���r;ЮF�o�bYu;<[3�����zà��˗�3?�D�lB��32� @�����A����g��xƞ�O��d[)���pr(�A�*�<uW>��v�7o�(%�Y��ê�!�E*�	��t�Թ�7,�o��d`
>B����YY[b�F���Ʒ�sLg'Jiک���C`�v�j�%(�ȓ{��}���I��,��I����b�!�r Ww�ޣ^����Ԑ` ?�0f�� �P������^9E_�6e*C� >�e���2X�7����U	�G����BY/E��xX�Q�Bx���=x��?}Dw�n20���C������:v�o�L,�l�!��ى0r��p%�3����kan���=�4޻����.-�H��`!��~�~{�����+��_�w�>1 ld������dwO�(S
�^fI�ݓ;K��X�B����\��r�2�s��z��恀���>��tqBtq~*��3ɟ��<h���u�K5��S���{��&V���`�P_���A�	������z�縞h����,��m02��Ix`$��ԺU�8H��~n �xܐ�5�0^�\�z���BV"�mbaϾ%_�\�q��{&���@\��SQr6��܄[�k�sEِ�B��4�33$���s�T ��@�� [ű�����{�˶�w*������cy���l�4M�b�{�����v�sʾ�(�]����������I�.!��5o�#S���KI����DpQ�A�mC�fe���,�*�Iţ���&4��5�՚������D�EV���9�%�U��6��n@mku̻.ʤ'�������� �j���3>��T��F�EV��S�aWR�����{����,h�QOu '�(�.&c$���3��,P�|P%�d�F�֨�[V��^Kj\�	�^`�%e�=yš�UJF9�r$A��^��R����#$���� �������GǓ(�/r���' �
f�hc�:�J���(����{������U>L��*y9Kp�k*�`�b�y��M54ή�Ԍi�:ZZ�����!�^�Cr�2��>��N�W��3ot+�,����b��2���r��������)��H@�LL¾I��ͭ@�C|ASW��-ĕ"%���G��irɊPZ>K���+u �ܺ�F�����FU��2�ɱ+{LSW�(V����K���`o��7Z��2(}}P�Q�����X)��p%�N�6� h��#�/���%�Bc�K+�дBzpN_X��������O��dmw"�9�Z��}5"�.��\��(/h��V���}��Q(�_�~%��
n�߷6�jS�� ���ʊ������ep ��?�
�����	��d���� ���JC���U�F���������������!��8<&�痴��/���P�y�l%ލ~oUa7%L�9.��S�K���a"�`�����>��'�11�FA)�����׿��)��<����v{"��o���TB�P�ރ��2�~N�����Ǌ�:��]��3B1d��˺�~��+�K����=z��)}��0�!�G�va	[a_A�B&����Ν39O���j@�$�����f�1��/�w��o1�>��K�	��PW�x���hc���Ɗx��A;VV���i��'��+�ȭ�y`s<�}J��;w����Ҝ��Ѹ�5��.�?
I��הU�*b���0<��\�}fp5'��E�x�Qdx��'���YG�5x��wtp�}�D����׿�L��~�]���s�7#^��4��*��Q	 ����{f0g���� ��|� ( �s�<?��m^�~5���H~�C49��R+����ھ����x=���/H�� Έ�j��JH�����B���0ɡ�,��o�ߤ�;�����
�{[r�"��&�ΦwȦ�H�~�0���ʊ��6�%t�!��c%�q�T�j�G�NT�p�*9�JZmf����o?�Uv�=����ua@5����T|������A��*�����5ݨ %��g�}O���֙r�C�3v��-�G��nX�i���\o�x�Ώ�=C��5�d�/��	�0���fZjF��*ӿ�74�s�_=�&瀷G�2�Z�:��+��S4hs�� ���+�������I�֘P[L�H�Ia�K�*�΋#����1��
 �������T,�.��#(�_�\r\����|�e��M-�C��"�0���
.{\3�hO����h�.
�N�A�^Fxhq�,�j�f�y=��@�%�������YG�l_pk[7B��B���#����|�̫5j?�� �tW��k��k#���b�_-��#4#GKs���x�<�M�FIh��.�cC*`��P�\�V�&�{�P���ZP�$���R1]T!$�
7ɏ��=U�"9Rq ʶ���PLd7�ήm
@i����*d�ؼ��V�� eoq��A�\*E��Dp����u�XIx����nkD�ٲpKߧ�vA�$`\i؝(������7At��X�lTzhaK�l_2D'�KIjX�����~5������T�v�~���( u�����>��Յ(0H0�Z]Yb�lV�,!*E�@(����9X�3=�� /"��	��M��@с5Y�=�dQt�W��q���u>e�[QF�+0�{���p-�/ݽ{�?z,�&(!W�#Q\?��������a�!��T�1ݫ����4L5��Y|_(<�f!o	}F�ٻ�����-V���Xh4҈ �(w�HK1c0��(��� �7P$�Ub|a��}Wi�d�d��x͟��cem~F�$Ǚa%y=)�9�sY<Vgc	Մ�fv(�5x�2�Ax rӾ��2��+�B	��N��C���\�B�)�����A�W�{g���>yB���H ��B_X���
�e �� ��=��FXj�j�*X$A�����#=��=�Gk���=����kyJ�ךZ���<x.A �E�KJ	���c~(���)�y�^���`~��1�����}���������G��[ⱉ�2ab��e��kx��
��Z�[�������^��Yx~���S�t�y����+a��h����<��M��^#5� ����O"��޻���=��g_䪟9 ����;�>nѯ������R�E������x�ʚ��Pp�0oxB&���^P*y!�V@~�A�LJW��2!�2-, /TA�dt��($.W��x��ĈY��`�`�a��c�X=,: �����Z��`��V6�^hd�{��}�T<�h�^pz��5FE��k:�ݐ��[�7���� O /.�/�	�5F�8�$�M��]/�,��4\%0�Z��`��d��g{�m�L��E�Ęs��SNX��A~FW���0y��l�(�nsJ?[~8��1�U�gYxwr�H��^7:�����Gko�^���IE��Q�rV�����u ���um�u j�mcnV.S�y$�w=k#��Nґ��>g��V�����sA�҈�@�q9T�ߣ���c�VK
���!{���哅Gc�(y*�pX��j"\�ȭ��>U���X<�V�фu�a�EYGmT�W2���N��j�����<;9��������'秴z�"1��|� �
�6��m-�> CH��i�6�f-ͱ��R�!\x�P'������}f҈�\��X�%�FcJ�OI���h�V��*�x[Q��D]"�6���8+��o��z�5�ԋ �����SI.������,�Xp���@���:�.�'�m3���.����*�����)L�,DE9����M�4K@��pm��j))]bI���I.�VY�za�٠��WZ𖬁���rm�N%T���`��	K�&�$�|����=p��A�T!���P`mM��7I�k�]�%	�Q�����@Q�G���J��N�H��̸!F��4D4b1u�ZMm-1�e�,-���F�"Ct[r����"�"U�ȉ�ʀ`m�*��(WR�����z��.%��L,� =�U˫�_�F�ذRQMY�a�n��!+3��g�������KZd�oia^ԑ_9�K�"d�Xk�)�ҹ٘�
m_j�)U?�m@+�1���WRP�D9�uED�Mm{��Gm��[�ö�dq�t]�]�듷��c�V�`�����
o}�P8(ħ�Gbe�2����a�E�Idu�P�Z<�jZ�H�G�]Vp���?2`;�SV��<;e���EN+�����xb����믿��ÇBV��I��pN�
����;ZP~@�,�����3r� ���=xpO�
bc��<?�ڥ�<���k���;V��<X�9���:�S�p[��9����Jp�W&�Z�ƼBa�<"�!��;<���χt~2�Rث�@?9�C����2����;7"��;��	 f�H�'v���2�����-K`./��A\@��y��N���E���aHK�7��Jk|F��Xf%��%�����`����2*q�:�}u&
R뛄���//�38����@O�������((��e�|f�������Kݘ]�����S���G���~��/�	Aʙm�)C�(��1i�l�y���c��/F��������O��۱B��"�	�"�=y?��Ч�����������3�M���[! 6b���
��3�Z��W��F۞�n'=�^���C�#7�/���,]�c�:
��jg%����k�|�C�O���6����=�;�S�r�@��~qq�^��'c2?#�X<jʴ�cd��+	��ܼ�iq���KTueaO�_�s:���;8���g�ߘ�i
#�y�<�����l&����gR�Rz����S�7�wLO���1��tV����X�Ы&�) /�_�PZɋQ�ߏ[?�=�W�n ,)�
I������B9�!�*�d.�E��dYԍPTj�L:H����B�>��a�~���M?�3�xJ@��e�fA��G�y_�~�o)9��48]��z�0
$�@�'My�`}�/x2;ک�t�y#�U�ͬS�H��ٮ�%1�5��$=ud R��LOml=��*zʁ���)�gzq�?�"Q�d#���&���9�&7�C�DYo[�h�ԇ���1���VCcԂ%�%qSa,�:��/���:���
W���u��!���X9�sq��0��;�%�n�T���A�h:o�+n��d]5`5�J��ˋ�X���I��Z<_"G,q�/���!�^��Ѵ��E����+���.��k �ݩ�Qt�:�j1�l�u�7b%�@��]E�x+��0�קv|a D�VY���riԢe�}%M���,V�T���-?ʀDaM���`aȪ�I#gt���@V��0:�	O�$򢥡P�����>tb�m��d��4�bsF.?�*���I[����.6��z���A�̨�J��U��f�Z�RRfe�U����I�Y�A�g���$K1% ����.�����́4�T���V~7Zܩ��|�DQ���J{�罨���dI�u��3 Xk�9T�Q�>K�`�B�QI>�D
nj�Pf3H���� �!�WRc���a���q�T�����W3�������u奘ˊM�Lp0njAZSDn�P�hx���@�ݛ7�%dzwgG�?�!d@GqmL����6ա��
��ayk��SB��/���/��[��Z�7����ݼ�.r
�P3 ���>J���H�Dڏܷ�9G�*�L9���5��c���>|�'�ak�����"Y�o�xOj�!/9i(����7�;<1(����+�66�2ȁ���\�� ����(�xSr�T�hhU�ʱ�aB���:���S  ��IDAT̉�><>��_v�4k`d��js��P>xL�"�q�M$G����i�u_"���������bZ��gE9RBY9�j�P���r&#�X�����ES 2�oo}��Ľ�s5~6f�pK�9 ~c�O�@��9�q�G�Ϸ�W��B����	�-z�����!�O���ؒ���~ۤ�r*�ڴ{����x́IyA 7�+C!��W���6�7o��/�?io�9r��"��Luu�o�����I����x�n���u��<�x��@J���K[-U&�# |8>�?�N�����Z;wp��������~\Z��Y�3�aYý͸6M�K�YJ�:U�^�{�O��?߇���K�>�Fz����>������ 
@��� ��)�"E��3:t�G�fOBO<���d��鶗˽�k�\m��u# ��S��~�,�%�N���������*k���[��7��ҟ߇���ɢ�*W�9d�C��H��ȫ_�_kmڎ�ݳ�~�R��)��h6T�u6)Ps�iȋ$d�@w�@�r_ r��d��$79B���3������6�a6g��_�QCa3%�� !n��!p"�q̵�JO�ڣ;n���!�q^X��_<3��cd]<"����j{��y$�/������(�3ƋgX,|P�s�W����GÁ�)�8�:�Ѿ(lh�h�C�46�֍��2﵆[*�R�鸉�o�%�XD�0��Y8H�E���j����Y�!M��
��;QZ�~�����v,d8���D'F����Rh�Xs�E����?]4u�v�oYL�˞@..E�����A�cDx��K�k��f�����y��#��G�S+�,��Л�5�f z���������MD�ax�^���_�|�$wEA�ׅa� `�7SB�1!(2Ȳ����t,;M�R��(��o�kq`&�G-���l�"Fx5%��	���`D�<k�!��Q���X}�!G�X���{5A�W�)�j�W�T�Eo��8�-K�m6���fAeM�4������}X&��B���7~J�ؘ�ƁtU�}�����M�4��W�g�ʵ��p!  ��* ���B��)=�����<7��E����d5��n8RAV ���p������$���:�����'��Z/ɳ����>6��@�D�$����
�1x��l1�f�Ɦ6_R'a5Su�5W�̵tΜd�p�}cS���fundN �}���fE��>߉qĩ�y�t)�:�%e�7�ނ�Hk*�wsxX�/�ʅ�g�4nd�|�2�ӽx ��H�8�&I��Sl����ԁ͏`q�d2�� )�h�� ��������q��Gm,������%�pNKb�nH���a�E#X�����0�U�#��f�̴X��9����l�N���J�b�l<J��E�������;G����D$B>1h�*A����9���An����$Փ��QN��1���L��;Ⱥ���-��}ׁҍD����]}~���{�{f�"�؝Υ��i����i��}�u�7�Q]�?�C�?J��$���j����pv"�9}�w�l�_		�Ή������_>�_��B��ؐ���ԁ K[��%Aѻy����w&�)�\��^�3X'��w�}�ipMz�}��cY@������C�˃��a��g �SM��H�F��`�g�Ʋ�{�ݾ���W���??t��#����?�[�)>�S�e\�L�Y"<\���ï�j}�w���E��x-0��ƈ%�~�ѥ��,̜B:Q�7��tZ4���'�Y�!�,��z����a������]���Y���=mo�hs����j��\� ��� �i�u��~����ׯ��펮��r��QIɬڠ�HV����y6B�l���'6[�M��d�۟Yޅ͚ı9W�#^ &�O��ϰ�B-h,�D���w��o�Z�b�0�N	�]�C��W|/�����W��S��[i1�O+�L�^��ɘ��J��3�T��T'����#��Ԕ��X�7V.����L���p���T	�ſ��
j�ɽ	H��A�`aji�����Þ<N;NF��D��a$�ﲂ�}�o.�qfv�ñ���z?��/���fZ�.<�1t�+`ⴘ����T�??p4�=�.����x��w�~�$Ju��B�F��\�Kt��L��F?��FGv��(^�XM��ه�kUKך����~�&-������=��~�W�*v�L�/�Ҿ+�CW�@�/�-Dd�s�\+�pj�՞����vY�1n���wxQ�X J�ӳ�٘�ٌhX�Xj�h.�x�f���U$݅���F��M��޴�����S"�|�Xr�ݫ�Zl>�}ZPȦ��M��/(�
�� ZF.��~����`ƟV�T��c S������X�<���c�j�F�ؖ�T�E�z�}]2��>�5ፊ�@q8�� v@Aafe�B|�=��b�p�M�ZDk����Q)*��unI��Aܱ��'f�c�0w������D�W���`i��jS��ҍ���Z]ܩa�
��������(�����[4����ɕ�r�ԟ�k�WB�`m�`.U�#�l��-�aQѹTZ��Q�b�
�ES/&�8� o��:5\��?��0q�/����:r��E�
�h������?>B���!����h���oZɌ�I�e ��gC�C�W��0��8hq��!;	���e=�,fB�Z&���Ͽ��s�A�F(HLB)�:o4�5B3xc�~k��j�/6��be�b�����-1[������ sǇ1I�q10t�(�F[g�@y�� ׶Ѽ�����R�6I��(���P��@�n8��2�?��Hm����g"��v�y/�5���9��鉃��b �����s�K�_����h��e�P?I�������[YR#Vt�ǯ��:�痝b�KϷ�4M�������`Q�� �˥��;�p�׌DF��m?G0/���r��e�Ao�C��{������^Rr\q��Ԕ`J2^f�ʌƎ�z������i��37���~G��=�������g��׿w��W�GY>�"D	d{��������B׻�~yw��у ^H��������ϞӜ�|�"��3;u�n��w��92k�n��8�"VXK�� ���紶�l���Ѷ8i����D��|>v���.wؙ�v��5j�����b������+!���%��tIs��h�ns�ן���,�e�:���,#�S�3��
t�69\�	�|�?f�%| Am����q���
h<8��b�`h7��W�(`5�O�9ŀ�ܦZ��r�,���;�|��-�l�>*��J�\K���e(�l+a��R0G3ta��S�d6�Mj%��f�5��i�'��Sƣ��K��_�u�����>��^�ĵ$����<b�[�P��i���t(+2�
'�T�\�BF����!@�5K5�GC�g�õ	��I���׃��a#���^���кy���9�_���rz�k��ه�����pE�},w��h{d�$�^3�9Ӯ��=�2���KZ�W�hij�(JzH.j�Ա���zE��#��M7"ľt����.|?����E��[T�Bg�۷R*J5�m��`v�S/~U�mp!Mn��v�(�C�g�����2��i���BL�%�7���h܇g�J:L�t`qV�`kV�� ���h��b-AX�14Xr��J#Z[JxWdY�4�� `�ջ[b3#�^Dn��QmS^��G�_�x��⩃��^�R�bϘ�/fM��FyL����rN����]���QxlP(���\屮���n �Ƚ�y�UYrt��$I����0���",Ni��I����}7����]�Ԩf�ũC[6^�ĩ9ӹ��Zl�m8���f�r沓��ٚ	+�'i�`m�lM�p��5�s�5�����k�uX	Izc�lAn�P]��lk��$��Jgn�~��P�9��^ ��%���t��KѺ��|�(��pf�UW<,�����Z�N�L��;�R�E�M�<ZƆ��R.���̕D2%���h��?�O�����z	�@��в�������{��	R�G�b�F#Gy��D啂f���3Zj�*��^��"�d햲,�w�5�oU�B���s��2��̑�B�R�d^tN`�D��1��/��IH[n��Wdq�!�1m���T$r��N��A�߾�g7����{qH0Q̾���^ +Y̪{<M�?j�M�<�%�L�Gqx�zd �����Hth����jc4�[1,ذg�;�X�y�[(n*�`���;}fq���Ϭʾ�>JB��s8��h�X��<&ֿ4h
�}k��OR�z>���( �jx-�V�����8s�$�V�sa���T�����mצ�;8����k��O��?ӟ�����-3��Chf0���~���&:��>S���Ӟ������it����{ӟ�H�o6���+i��鹷)�������Dl�M�kI3d�.��|"Mc��
H70��Yud�s��͍�$r#Gy�3�������J}������Ͽ�����?Gq|LS�����i��|�Z���>�L��ng�^��ׯ�����;�{&�8K��I�U����<%e�H�0�9�(�޴��d%v���P��0���f2����l� ��j��@�f��9 ��Ek��_��F��Lq�P(�_ �8Orz&8��ui~�D�^/ca�t�mR��"��q�+����QʺjI�����>-�*���Iv��oώ�D�S���6J?�^4�˾ی�y#����h$��kh��>��$�/�j���Q��� !��Kۈ��.g�p\[QL�jWu��٣�!�2��\����$\P�b+���99"�=I8��s�y�P����٣ָ�y�ǳ����nН��>���p������Khq&��	+w-�W"�+"�5'��Hz�����#!r��Q#�e5{"�i����.?���OR��������p���i��B$"�Y�k2x�6�7�9E$K�e�ۣ)Si�j����n��౲�ɣX���L]H�b/a������N�#�q H�Hn��s��H�� ��=�@�K@e�C9wp!ilO�i��)�����J15��`r��hhIjp��z&��,m.�O�fP�4��,��7&3�0�X�](p:$�A��dGEcuX���B7�z�����������������j��*���7z�=�{a�tP��Z��
�H�9uP �>LM�����MQp���d��R�r�{e��f�I���'U����S7D�U���@�� 
�k5�d�����Vj����Ϥ���
�{U��ښW��1�"7œ���G2���P�\�)�#�N�2 :YT�A�px�Hif�7�93
���WС��;�O������k��R�l�� ��=�歹�G����j�Ǡ����Xg��U� ����59r�ԯ;��Ԁ�ApJiU��N�A���|,W���d,E}�P��Rܨ�D*h1:'�{#@����qv���tv�#���nS�HWUֹ���IKI�T��f�Rŀ��i�@��Y�l?	��6B�>g>���8G��D���]w�H����O��G�
�T4N�UgA�(;oΗ&�OH�6�y��3�t6eq�.���(2�Z�7 "���h�~m���Q@ܤ�N�R�u>[4?׫�[���ΧA���4c�_B�"}�9�&�7x_smS�t���$�Uk(H�,�nN4)ʬxl�X:O'e/e�K�����@�����~������~���Ы77⼙�6!_F�a?�?�s��G�� 돿���?ɹ~��?���}�#�cx?m�o�N 4��Z��2k�-�K5JL�5��[z��{��/��/~9E�/?�W�'9�~�w�����F����~�H��/��plt��,6��rK�� {v�tJ��[mH��Vk���޼y��o�Ї����$-:�Is��L��l3��/ dY��Dg�>8��;���ȧ�����l��o\���J��H���0VcPf%5��$��:C�7^�+�FS1.�*O%㥗}(��"Yޗ�%|	�Zb����MY��<=Z��8�->v3��[+a��q�
'�}۾��H�0I3��������R{Euq�@��Jq&fՍ�'0b��]�"��
x�"E��l���B����nb�I����E� Ā D��1�=TM����fP�{����/Z0y��y�
�t�3{u�����R��7�pwGGk�'1a�:K��x(��=����������j>�Ë=w��k@,���,5�u�H
�� �5�� d��r����/7�4�9�>�n��d�bk��,mR��H�μt��O3���
:��Ѧ� �a��9�3+�Z�Rf���-�nx������M0 ި`�"Q�-d�~x��Pý�u0��@ S��)fٓ���d!���b
#��c*���󨛋Ә��E��ż�&���N0�R+�tq$Xҁ��Ʀ��P��Р��������F��Ʌ f��\����BANzD�8F�� [�3�jQ�:j$K��ɟR3�#����wb_6ݰ2��,F� �͛[!���w{=Юw��F�Z��k���l�����K49�J��zI%jVܯE�*hD�ܘ��j��c	�Z�ee�![�𶺠o��DI���ãʎ���!��6��!"ZcA�x`��g�Z38=�^ӭ �Kx��F����=\��}����"WL�����D��r;��-��b)A��5��ا>ߓ5��Z�4�V��=�>P�8S�V�,��jT%�7]$j�^i7H-�ϓ�Ċ:���:�~p?�dq�O?̃��}ux�2pq�.�g���@��x[��}�,em�u-�z���$/_,bXl]i]g��{@��ϟ���G��9ʺ�te��ȋ	�������˹�ck#��$����r�m|<R�w�T�&��BU�UЋ�rNATGZ�y��<�U���O�>jt4� %/%H��A륙�X���쪓�]w�@R)��5��H��4RVd���R/�=�w"��)���[z��D��m�j;p��>���p�rmӯ��mW��?��?���i:.�k��k����O��%�i^/�+��e���܊��SLPss�)�L� Y9��y���E�Un�o;��N;���h� �kp}��<H�λ�A��8-�K�_�l�e��./��k���f�dvM&,b3i�c5�ʨW\J<�����p.n,�����&��[�5��k�_3Y?��F�P3�h��dz���)��i����+]o�~��A�Gf�M��"/P�$�e�L�\���nYA���?2d{���3����3v����_�.�邰����78^�
�J�lS��<67���B����#=�4-��3���'��fmXk�p0����J1��rʻ2<i�:Y�	<�n�"$�>2��6YH�m
i�J$^�QH �@؞�sWbG��6�A�]�����P�U��)s�W=��x�t&��Ȼ>C)[���/�20<�j�L�fL�.iq'�1��3Dv>�"��4G�5=J��� "=��'U�H�)5"@���ym5�Q�O��3�*��E�XT0���/p�����*���" �ٸ��p������pQ�Y9���D�#��$��B{@r j���b #��62?	[��`lN�h/Jà�FÀTAU���J)n�CQo;��[�7���s��0����M��s���H��#N�H0��yD�`�Ԋ�|�k+b�P�Ԑ�ؓd^��ޛa[4R7V���d��쀪D��T�ԋD��ջ0��JG��bg��U��I�����k���ry%ulL|fB�&��k��� ��=)kb(8t-9Af�� �����4=���nyf`�+�d+�(���{���.�)3�H��2�5�c�;_T�{�twG�t�+��' ��֓V��ƞ�职����=32�g�D�s��K�M3^ԁ��y�	E#��Ob�_��j4��ҵ<K�*`	5�x��l���&e9���:��I#�7�q$�.I�z=�6t�EJ>@h.O�A�T)�rP�6�-*�~�^#fD.����ߋ�ІF��P��T��j�.7ZGp�y�6N�9u9*u�耋da��;@u_$���S`��P3D5P-�Utv�#�4r<�b�Uu��9>]�1�N��� �jd���u;�ѻJ�r��PN�Q}�Q9�$B��j�K�7Z暻��[ڎ$�r��d�`���JP"@�,)��Q���?|O��o�F��AS���6c6ع���ͩ))��NR��RS�&Z�Ek�X�����)k�~d<>��������������Ҩ��w�������iډ�Fō:��gà�$N�42)��=&���i��9�h��f�Ҟp�N���4%Yp����{���i�ѶŖ��r6<ۖ�3̖�@X���(9t�v\��ٚ���t�(�]ƸЎ�f�ȋ{����+���������s��-�,�ګ��~�5��ZO�ث�L{�8�;U;�V�J�Ɵ}|{տ��#����Q��@�b�7�Q�ƅ\�C˹�� �	�'�e���F�OA���By�o�^N�C,�Y䛈΋v�,�X
L�j K<g��$1#��*�h4���I*�Vu�p�E���ffZYn��78�w��I	��q�T�y2ᥑ6�J��,�
5 ��
���C m��եM6W�K����"�iιQ��ʗ��f"�Zʳ�HV�6V,��H�J��Z#.�q�z���ᴲ��M �`(����2�ūx��(�� �9��mY�X�fT��m��I�,V���l)w�F� K#M8.��"_7BC�qa`��:x3X�`Ăv\@�f�j�`0)ч�_���I\�1i^�F��p���W�9�+�Â��g��w����+��*Y0ގ���!�yb�В�k:���i
� A��lt1������sc���r�U��3���r��*\�O�A�?�_�|(�	���L4��&�I��.��SN�>�ȯ5	L�՚_&�٭(pm����+s�n ����ѵ�F�U�{ehp���=��?�i�2� K=���2����-=�pZ��{�AOӵT���D¦9� ��Hu"��K�Nѻά]G�f&��4��Q��ƴ����KBb��t�N�k�T��	�4�<)�{�����H���ِ�}�g!��?:>��̉�C3�Tv�<�S&��My��_�j!��T�Ct]����@dMf�>N�f)��'u��b�Ҭ�],�y�0�����)�j'j����2~�6I�0l�p6��T"�p�U����Q �D��� ����S��R_�3P�D3G�d�Г0�im���J�BAFƬ����X����me��z��wh}�]Vw�}�6�{��7>M���3"I[�쒋��st鷿�-��O�~���#�߲��l�*{��֢�ɬ�6��F���I-���ZC�i�l+}��I�7�e���;�����W��O�J���t`��#�B�a=�xl�ʖ�ҫ	Iپ��XS9�h�2ʤ)5j�YI}�1�����!�'�N�F�)Fb�,l�d�&��ζ~��#&:������grV�RE6�؋E�r��#a�d�ǆL�Oj�l�Ȳ��}�9f_�n)�8���`p[+��tP�{X}#^�f���f{,����H*�{�9����5�u�G�i�vB�\.Cp��#S�G��,�}J��d�<^�W�s���Fu��F+�lS�;@r6+eĎRoS���D���D�D���Y�=��N��g��JF���"
�1�'OG�2�M(�B+�HX�=�O���N��u6��� �d!;�g�2�)bF}�s<�t����D륤+����nV��([�EU�
3�̈�h�V6��ї�,�6/ܴm�%��*�Xn�f�xj jK�䝯y$�$-�<zs�"�i�:����Ss�3R���f����}����.Wf��e K"VÆ�r��q`1�r�eQ	Mo��8������H/��M���0Y~�p�ų%=j֜�	 K<���g{��u�XA��jQ�3E?"�T�2fC�(�F3��H�ٌ��m����^bh\v;�-lB�@�E��^X+TN�@�f���ԏ0��9�wc��'�W��#�dt,Nb�wC�[�RH.b��p媠�Z�P ��T3���k��`��8��y4@1b?cA��&c�~�� rK%�{�� �2]0�Y"�3�d=�h� �@ `"8�,������Q�,�һ�� �^�5��E�'�!6)Ϭ�e�ً���d�{��0��
p��j���-,@�3�~�B��aIg�@�6�O��Ig����1�k�8 �ؐ:�<� $Bđs2� �Mk���u�5"=��5;$�\)N�$Fh}!5\b�������S�ST��Պ�Fn��.�@�"z"�����1��Z��sP��X����OY�TgJn�^�����i���lp���$:tk�}h�����1�
.������nNRw�La��xGu��c��6h<[]�<�4�>��2i��(���������ՙIm �]i��ka��¼XrJ����tu{c��B����R�-1�fc�$r*v�R#�����l�>~������&��3Q3�>���a�-!���]W��k���8S�B4�`������gЯk��}���t�
C���iy����ߐdL� ���0[�f�-^�2H��ʹ��@ӓ�?����k���#1R���j��x)'pȀ���{";�ln
���}f��,}帖l��~/.i���L�����\������|,��jp%@�^5�+�`��9����g��������B�~A�?>"�w��#�xw%pb��:캬͐��{ڴ~�Ej8.������1��u6!Q��w�W2�#K��V��f��ӣ��� _�,�ZxX�ޗ���1�64e�b�Z6��2iL��׉D�q�u52I9�^��עobr���.��Y�ॷCO�"���lرTcSrg6�'S0��ۈ" };
%[=)���	H�a��lYx�����3ij&ϝ����>l@�Q!M#1c�<��)*��f:������g�Z�۫ \�W�Ak�O�\}��髯
Y���&��F����j��e�+/(�*�K��,4�k��y9�t�i�x�`����E%���ה3�@�/��W��e���4�1[��c�S?�G�4BaS�G3�������=�D��hF��z'�X�D1̩���f���t�TE�T����-�O��*����^�Q6NK�V[D�̶��D݈`C���?�Զ����ٻ�[Nfl��*{F'u�ؼ��
5[��7��f�u�bc~����WCY���{�5C��% � K2�y��6��l���΀iW�.���+f��hf��H�O+���S"?R$\b��&�������ٞu�juʑ����	)�� �`D:N����PCY.IK��;ZPrOБ�m�f���F��2�fn�G՚Q̈� 2��!��R��Q�� -C4N�#U�$�ȠP�+j��p��B��q�ܒn�<w[
됬�("
:d����9�|����?7�d���C�3���>7S��YJ�|��;���p֕��"��,���>ǚ��L_b�A�pa$���S���֨R]��Z�ό����*p��׉Yt��]H�@8ⷫ�4�g5����˟.P�������׏^��[����n��R�}���)ά�6r��D��|�}ݝ������ N�����=�2���A!����s�������>G�t��ʞ�z�q#���������'9gYS�{��^1�F�eo_��v4L��m��n����n�����e	}-�m�i=q����HvW�F�����n�js+{�#���{���g�������5q��R��ƽ�s���א��0|e�*��2�S`�d[�����d��s~L8���p�k�����QkUf�_ (K�8��a˧�P[O@cp^�߰������L�;( +!���'v�ۑ¹e�ε�@�5���q�ؽ�6)"���OC���l*���P0w�jJBܪa�0��sVK�.G�� 발&��Z�⎸��@��Yd?N��avU��L�}�&����5�:�q�G��f<�<�aa�/U��E�@3�vH�0<[2�9yF�<~d�6&g�,x�?���a,�i�~�?�d�N4$E�ض�Ľ;K����h�k�z5�axM�V���45H�K($�bQ��/��C���@Ϥ�K/�	�W���E��W%�+����3R��X�W���� cPfl�x����(<��蹿yme�0!36�ʢ䩄aiFX��.�$����%��D�Jx� p�Ir�(�Z�)���H,R�Eb�����z���9�l�����)��%�>C�x9o:�5s�[� �v^�!HB���w�=�%lS��R��zp.��b��-Gij���Z �g��tGOg�2�qc�����r��w�����K�r S`z��_L.�ΌM�:�S���Y$(/~x����"�XyP�n������>&;�.��
�sA@a.C� ��E�Fe�O�W�c�.��~�w�~޲q��|^|�p�Xg�e_k��$�t�l>#�tz0A����������(�x0��dcN��(��g�����bbk�[~�n�{/��x���j-KQ�$�9M�B����/W��������Jk>���3������z�s��Ŝ��V��zY	J4�0j���r5�/m��\W���"+7�����1<�C���,�������΁&�����;Lf'���ST��.����.���i�y_E�@!�4���������E����֚*Mu��!�U�^i�����o��;�t��\�����n�9J'9�G�-��Y7܏������k
+�r0P���^zLt6[��F"���{*��܋�m�אR�C��j�mSB>ۛY޺�=��l]3	��K�#U�Y�NU�#��_��D/0spY�����^t�%�䕧��Op���H�s-����i�*K�xn��j����0�+�4Q�=G*8"��:��W��^h��`[Q�!F��RS҄��N_q��ǝ�ǲE8Z���2a���Xĕ������HX�b��ٌc�)�b��6e�����O�5I��V.+i}�F�b��8��@�_�_���	E��`���jot��j˥��������ym.���\F�\�/1�νXZЀ�[�l�n4g���^��D�=K��7p�i9"��S<�Q�bf��b|�FKT����N�=��Ȍ-�tt2�_e~R�/^rI��������9d�ژr=���̾���j�JBek�����zl,�F^�.ml�S�}�p�	 %y>d�䖖FdLY�ʎ'鰳�aJLE�P�&���ԧ�g)����q��F� ޵�]Y����G�D�l��ɒ��}�ȣX�
5Kj��>8i�%��\ �gOaӾD��~��	Ʌ�[n<~Q�����}6��#�Y�[f�N��֔�;M?�k	�i���y�_Y���m�ձ���}KO��Z}�ϟ4��`��[qG�̔0h%��#Ҝ�/��\��4��}�Q��~�9�{�2�}O��qkdqy�k?X�q�uq�����4��SJ�#	']xB��i:8V��Gs�`�'�	��^��|��R}��׌}a���ƫ��W?M���)E��E?����c/ғ�HM�E�O;	K G ��@۫�v[�m�g���`��?����ʺ��dZ��JM���rwG~��~������]�y�S�O�=����,̤Zfa0D� G?�>��I��؁Չj9e�)��}\�Ax�E�}�����~�������[�����G�gg�|B&���.�9���,3{�웦v��1�}���v��,�}ΔZ���a+�L	�r��µ�R]��LSote�C��RD&���u����3��o�/����p���mip� �麒7�}C���R�c|Iqԣ-]V�s�M�#�M�B/��L��`�6��o�8n)c4p���x�y?%�������5gcK�G7�d�X|2� ����V�I&��-&d�TQ꼙�i������pV���܅�
0֊N	9���v8�·\��~KE"1;�Ӹ��OV��i~��/g1b��l���M��Aɡ��d�⳦��x�� ��A	����\��"�I�z�T��mo�e��H;��JO�T�YD�TI��ڛ~?�Ft�G�D&��V��!��`n���I�d!*3�F�1ҵ��+K$�_gw{#�J��C�r������E���E>p�_��.88"���P���D���*--�un
]I�pi~"���J�+׌�������3lL&�LR�B������|��|��oi�Լ) Y6��J�}K���2^�.T@�^�t�ev=���`\17q��/�Y�}��.8���Չ����1y�)�Yh[4yV��Dt/ʨ(u���W(fpjZO��q큥D���D򇅯��]*ך�'\�O<[�����H�_&)L�TeR�HK��G���4�.���-�[D0��I����R[����*�b_��g���s6��,�vh�k�0o����6ʓT��#ti�����fD�,�dl��i�4��! �5y3Q��|-�?�-xώj����,�V��b5pN���j���*�AŖ��lu��0<~�a7V��5}��~�||e�o��<p5��u[���+Z�C�|W}&��9b��="Z���͖5Q4sF"_��١{�6	�P����g$?���6dmh18�HY��#��>d"��`N\�p8�݇_�������u��A"�ls07�z)�����%,���b�$���EK5��b6���R�z3R��h��m�o$���G_�'穃A6y^������3[�ՠ��Z�u�����r�%5\9u�k׸���R�	ӖN͈Z���ľ�E��%J�j���j�@�꿼X��5l+r9�B3�e��-���� О�@���W7H� �%;){�Rʵ�i�_��g�웬�s�R?f}5�m�C�>�����
ף��5"p��<�Z�P)�+]��,�`�V,�u�)�-�JmB/�R�:��Sj2/֔w�HV)���晥*[-����R�YTl��@K��p�	?K��DiVxu�
��Q�u$"e�v`j^*R�qs{K�߼�%�f�m��) Y�l�g{W��6]�p�L�]`q/���\i^&��dF��Mj�ظ ��L�q���Ak�T-��*_c;Ҷ��7J����4��_ǣ�0���9��j����o��Q�e�"c�Hg���g������qcR."e�.\�R}3���iZױ9�2���� 	i;$%��H�WG�� Nx' |YH	=/��C�o#O6��n'Y�D�x�ڬt�)��.�c�֒aޘ�
xYyͳ��7p,%Ad��(���$@�s����� �4~����Y./?Vu!	���� ����l�����|�gL�j�TI�[�9G�"H�~&�g���:�'f'�-���.��� ����w��[��W�ܒ� �c��b���(;(0�P0�~[K�����3�K�Y�'p=�PZ�_l�O���=5r�2�T�EW�F�\�hF ��{G"5�˹�Z@'��@v݈,�C��� C�̇|�����Ն�/ Y8��v1 kyޗ��i�U��8�r/ޛ�KIp��o�`�Ͻ�o@�;�(���B�!�]�˹Y�Y̪���<X3X���+�Ϥ�z�nv��:>^��� ���C�g���F�R�bĎn����qs% �)ݙ���������{���>9]8u[�ö��yRL�KݬQ{N��cc��J�������p<��R��A��7;���O�{����>~����7u@نm�}�?��ǩ}�@��Q�R�~c�S<���Ie{��jE������ck��[\E_m4鷲iZl���ģ��N�2�y���n��lW�%��K�z=qO}��t�K���_�{�X��~���u���!����9~,2�}I��	'�G�Ӹ�=#d�Zk^h��W#PMzAj��b	!V)��b��RgCE��0p*�mέP�<��]�qc�y�T%UG PHA��;�3���������w��/=gEq|��7���v"x���N��"}�8ב�c^�^�u?�b#��,����ة�,N��T�"� h�q��N�p��+bVV'3���_I�ُ�-������]�F��
������'���"BdO�f��mh~�T?j&��U��4�ݨW^ݬɥ�h���kƁ@M�o�LR~MKB���l�Qɷ_m��ePc5b�Sr�������o]Հ����^�d�-�����u"43��9�c�� >�euN_�n���Vg 43�
%6��K����s�́����Kz�w�O�x[V �#�������3�f�hQ,*�,��~[?�����0~f�*iHqMPW��]�cPf渱�>��20$ XYY�k�۲z�E3�k ��\��$&z��0�Xq�E: &�`�Т��T�u�gJKe�~[�z���S/1�(R\ᜐ�# �9]���UO� y�7�_Ȣ�I`��@1y�e @��D��:�b߈��Ȕ��"�|5���Q�C��E_�~<�g_
�J� ���X͌���&�28�f/�p�Kk��Z����ۢ3��뫼̮NN��>y%��F?�웑�m-�ϩ�U�.%ֳ�.	+�U���ݾz%��fk|���Y������5��R�$l��q���y6��p���8e��������Ý��d��ӑ�rqKvƾ�7�[�O�H
�Q�W�=SN��,5f��ݽ��\��� �gϬ����L���;j�5=�f���~���=}�l�͵~��DSy���3G���u����]&�M�m��>��/�t������������>7;���0��֩�j�D��7�!Mu�p�@�������[�b5y�`ľY��[�/��ao��V/D-���lz��2�x�Cǯ��}d�������M\B��k@��w�	����vYLq��WG+�[b.K���p�%���0���nB�Q�7M/TlYld�:���3պ�	l�M[�h�"�`���RT%*�ӼDgs ����p%_�~�`"6�A�e����4�RA�h��t0g�C�~���Q\i�(��ז��J�}9{(j)pQ:hUL�J�����?������7��4��w�EX95��bv��}rcW����r⽲��`+�E1�E��lk��u�y3�~�A/BX�mQV�d�p�����v'�O/{%o��t=�1* �0f�33|�GX3#?��p+����� �ആQ��<P���NѪ	@���r��Z���4A���D��>e�oa��t�z�U��3?sS��ML�V�s��=h�m����{�I�y��!��grD�X��z���'��xj��0n��Ϸ@��3�t�PH+�ԣ��k�`�a ˭K�:�G�P(@3���5]<��"��x=c�_��9Ӝb��>��TrƄRn��+��̴<o�7�8"�!���h��a�8�K]�=�Z!ڊv�!ӞeM󿗢5�.�6V=�?���;GB X�o�,��랆�ќT��l�c.��~m/,"�Ͽ����BJ��~�k_Q/��놑�p��6�fo���ߔ�di�P��h�)l��k��Zh�Y�v��oz��][�rΎ]�=ą��ʀ��*f=��%N2a�4�A>3Ď���'�_�뿄����_�Ç=}��ȹ�K��h�Ӆ�w���+���M���<qSa�v{`2 a2�H�a~q&�A���hC뷊�>�޼����4�?���v��wwCu��v��~�t#�,f����.ۍE�L��w�hہk���x�h�o#��y���͖+�ֱ���T4�C̰��F4A���N����A���{�%�}n�'�υ���~���9fm�@w'���6�|���;틗r�M 7g�	���2�r{½U�V�߭�o�k��*\[�֊ke[V
����.�� �Vq�*��30*�ƺ�_�zi�e�Fk�(y�~��&!B�!ۏc[y�%'Y�F7�*�a[?n�������� =��1���x�6	Ո5�ZQ#ɱ��9��p����4����W�]��.�b�D�6���C��W����׊q�L��#��$s����=4���B�1�Y��k��g��q�?�_��.��5Ee����\S&5b֟K,"Ͼlcx���5}"}�����e��Ә�@�믠!-�A]���kzO>��X��Rq�7^Ki�2,꼗�(F��ϗ�3��m��!����R��ĺ��i�����@�O:.�nT̀)*��r$q�$ a�7�7�>i�� x��2~�{2LKw���A�?�֤�{8d���GjE�T������?>��16�(\�b5�PI�^/��F0͘O���^��hq.�z�d�����������t%��۝��9���;�i
��f��ǎ���3��6S!R�́Uc�#��
[�Ѭ��{�II�4tUq=��c_�!:������C%��T��龮c!,�"	Z}yx�֗C��Z=q�1�=�"����Ʉ��Ky��Io=����O�/m��Ǌ��0*��ތ���9L�%���J�F�ƪQuflL���\�
��0n��;:s�vQ]�8�t8�����#`�y�N��f��rՁȅ~��gz�+��t����^M�;:7�L�ǠuNu�6�L#��{�s�=4ay�(�T�ڼ��d���۸� l�����<צ��������ˉ{���Վ����U���n�]�T���"��\G�j�yg�.#�b�L��E�.�mƠ)iJ/5[Z�U/�Mԃ�C�I	A(CԨA^�˺���P�2ÖY����u�Q���ٷNa�Q5�,C"�8V���F�����`��~}|�f�`}��.�R>�C-��Gz#2|п3r3L  W�^��<�C"7Էi��)Odx-縤(VF-@���o�yi��ت��	�+��b^����n��J�8E6"Y�m1�
�u�Oּs������SI4$�S����/�|������r�y8bé~')����" ��j1�`�8�(��'i�)�wq��T�B��c�%����sށ�fT�W5"�(Q�N}<'���Y�5g�>���2dʠ�t8ҥj���i!D腣��Yo��&��M4�J4kF.[[�oL���KEIC]YM�i�Ya�6?��;,�LZ��F��ی~xu ����#Y�[�Hx�+��C���YVܾ0β|�;_�ׅ1+�!Ƹ��� C]P\�u��y]{s#�g�����o%L�H���.���K�V#��oZ̑�����L����=�-Q�%�Q/��If���j��C�k����ЬY(�@��\S�SI����1%��Φ7�j���RIs�s��!��W��W��iYCZ�-@��⓶��m1z���6���A�os����4��$��gfK;k�6g�h"�p@���FX:?9
����.פ�a��,��=��gq�4�b�ɢ�A�K���K`�׊�����eV4���DgjQ��+�Xy�|BN^D��_�4׸Ƕ��8�e�����s�~�\�1���|��/&C3]�	0�~���&s�ʈ%�n�Y�������n�k5�'S�a�/�`Y_�tw�@�����z�A��~G%��:p���{�����2��)w‘�<�jKĮ_s�2���H���q�/{���FG�_�7I�)f���ҹ_���0�E#X�F�X9S�<��@��;&+G�ͩ��-������5W4��4p�j6,�7�R`��s���[�Bp�Y>��=!�x��k���"0`UC�%y���A4�/+��N�4���y���w(�~_3�� YvD��Ul�;J����}��^m8�w��+=w���?!��#Yf�/��������$�4T�|�b�ػ���0�w��`�|�Nq����'�$�� t�D��2v[OC[��l�Yɏ@��<���|�>�J���1j��X��Mn�ť"�xC\���m�����E�� ����O���?�g�%#�����Q�<��oN�8� p�Z�79�@��>Cd�TMkl¬7��� �Z�l�'3N5ϹM3�Zd�?��;s��dr�QG�[e*S9�d����v��q4�CJ��|�ד��^�,M������A��+��C�������aa��z��Z)z(,ms?����'68��kk-�[������K�N�uSY�������q.=^��-���)�<׃-���!y��i"����3�������|f�����aY}��vȥ��ڕ�����j���$�yB�]S�渺@��5�"9C����Z-��$� 3�|��[(���N���7׶iJ���»���_&�f��<�F�Y���� D=J�Z]����P�8]5�Q�tl��NvM5�[S�=��3��� e����`�䵼02J���ri�Q,�稷M�k�=��ј�Z�uʨ}� ���W�l�X\=�Ș�${��\��笯��fY~u�2zՓBL���3kV���d~�K�KF��u�;?
���Rt`q��(��e��C��w�'[G�,�#4��#��ǚ5��e�e���wN�c�.31֣��던��x<	9���$���~߯� mT�=s�Ij���^���L�>0�OU��v��{�ƿ<���@��Z�]����X����I��s��uWG�$T�B�1rM�e�A���N�}֯9��z��Hֹ���[���H�9l qW�bByv"�&v�$�zj�t葴�IU�d���󓟭^z����E���~�]����}�Ԭ����������N����P�;!���P�6+����C�]��S���;(�읭dC��#R	���C*� ,�p���V�m0|F�Y�&V`V^��t9M%�����&4�r�5HR4y�A\��¤$���L�ߵ�T��_i��,|������*1�����
5f�aA�-fku��?���B�z���6IZ�ty�s9��c�5Wωe'5c���{_��2�f��w���#�� D�LA X��W�G7��-
��[�����h�b�!�A�;���-n��4�@��ECdPO񅻧������<�V��~^����*�i�a�\OV��=`�<���H���Ʀ�XD����㴖v�1-�Zl���G!��`������Abѿ�j�����xH�bl��Da���d�5W�P�޳�����s^(<0������焒�!0cRy^5���X ��J����i���"�[�6'��h	²r�A�����e1\,�]�?AG�(��VN=���%��raKB������������aV�)C�7x
���} �-�·��k�Ҿ�Ɖ�b����j��,�4���q~I���MB��x�1��pK��᦮��F�Eܫ��bOD�1E8��x�� �Y���	7��Bf N��Ʈ��gc̆:�MYi�n�����XB��:�ůz����QU�"}�GrJa��0Vw��,�v�$Q$�̄>��f�,���:a��cL�50���f�ۆ,bC~e}M-����������QS�4�� ���L{��s1�v���%������J� ��ܴ���]��?�G��\=����27g��09�+:�Tw̚���p���U���- �8��`2'1@���M*cL/k�RԐB����1p2c	�}d�4���z�8�����]�v�0���e���ϱg�x<0�n?	�����6l#:��>��,��_��\Ӊ6ӡ/W����Xg�������u��;γT���]�үה���y^�5���
�>ڋP��х.N�k�� �T	2�a������z$}#�֐G�ڼ��dl�dz�@��W���'���j'Ք����Mqc�[��۟�gg8��[T<��~>�N_Ƶ���5R�P8f��^��j��u�7o-�,� �oBo�mm�L����yK�d~x��^�H���]>�����w�2��D̥ޫj��oM��d��d�p�����бԦ_㲡�-�ڌ�N#"h
m��Ƶ�,1�Y�qCPښ�O*�m�P���	�w6����h���z��,�o��lƢz�����v�ܼ�V�\Jϋ'}o2�*��3��Rh!Ȱ![�i��<Z���)��R�V�5[A5�h]jd�!�k֯KR!X������E�PmS�?��� D�(l|/�/�t�7�1�o.P�N��,z�h�)]��g"h����o�F$]ϸ�\�����=�|gAQ�EV��V����N�����w��kϏ_�!�1l(�ed�$E��s�Ꚓ�L7f����X��ă�ZknԚx5Cҡv���� FI��>���x�\�,p�{6z�^�a�<g؍�((����v�B�qv�E�T(��Oc[�ƪ2J�\�\aد�Ӱ�� _��W^Kc@d*�q$���-IS����xB�*��� l��gN�"�Β�G�X�PÚ \اgg���k�M�s�\�� �z��z��������r���-�ULCv�4�R�����(�X&H��1�@]̦�qۏI���6��������z!c�G[܀��^��Kո�l֋��daDn���LFB�T��Wa��k9���K��q��x��M���-��0��h�,���-}���������o���r8I+��z^�CA�)�b��ii�Q"[J�e����&���n1+3�����X��	&���Z����G�v'�^�_�i{u���}H:�%&��Zw�'�S��6c�7Gט���n�uka<�:��<�C����뿷�3����ҪՌ����0�)x�Z{�&#T�$������\;T���)6��ߒ�!d��"E�@�3��\�o]PFa�s��'_v�d�BaAI{49�	�A�%͋���
���/?:_Kc\��&E��ĲF���&'X������Wn�e���C��ӈ��c��X��
�4���ζ����}����0V;�qC�V�1U�S��]�R�x�F��"��(N���{6FnJg��D1PW��F��Q*��*Z�7h4#|��L�� V�7jS�K:&8DiJ��	gD��r�H�Zy����.l� �T��U6���t������)��Zq�偦��&4�V�#��$4�CI������6q��Hd �%���hk�C�6X�ޫ*)u�-��[ $��yld,���xd֥�j�0_{�t�ǧK�����`��K�mXx��(>y�s#�H���j?�#���x���Lq��`�ưKK_���R������Z��m�H��J���s���� \n\��1��A<`��,�z[��k3}g}[k/Z���X�H������h�(�1����w(Z�{���y�\���u��!�n�A��n�<�?Ͻ�?)ת�6VL���ϳ��͐σ����2yo.8����%MI ���K���'���ޝZ����9�:"?fV�f�)�dj,��)43��}d�v��w���Rf��qpTP�@�ht��\�J�T���u0F@�1O,g��=���q���o��{s���w0���������^�̭RfI��=��(��+@��^�&c�v1]���gw
��T��;�R��,?��qh{5v�s%}>��O���޾}E���o�����y�r
wv�"#��-=?o��Cu�?����V�p�$���̋�iW�������+�����W�27�>}�H>|�O�?�;O�v�J뛭�m�<r$�J@ڍ�%^o�d���Ӈ����=Ng�$2AӮ3`�[�G���8����_�}~���(��Ͷ�o~��޼~EW����p�R������J0غ�����J���َ���o%l�G{�@Λ!ޒd��zj.?�ڭO��f6�I"�]���6�寕�jv�pL�m�/���f��n0${l�Z�7����o���?�Y2�2xl����RA�H����wV������I���?IƵ�7�sFy��%���h�������Y��j�q-�n
�:�� �Z�H�z�ʵ4�a�)b^���Ƶ������h\l��4����"Ki�菋/��4t����n2
�>苡��'T�_ϓ%�Ǣ�P�"�J����<��Zg���8.��{Mn�;J��lB�&m6��hih�<.����}�(��j֍'}��A���G	gW�^�"k �B���l��	T¥ M���\jja����
���!�o�w'Z���+j	��T��I��z�M��r<!���X�`e<�>M�Ԙ#��d+��8<U�`�l]<s���y,-�S��Sp����������������k��k%�)��f������@[D0�܃e�V��񅘂���h��x��;�m����O����`w�g�u���ʓ�����|g����t���S h+���q?<�k�Ӛ~�k&O� `m�	��y�ߕΧY���FE"�T�K�GM{�P&u�P�ڦ*?#��6�<�cieQ_
8�RQ#ܞM]�g�b�,-���V����]�n�5�8�������O�0���@za[\w�׺Ο��#��D�v��Gľ�-;'����sk���O����s:�0'�o\^�^�S����4k*����:Qp� �%
��<ď7��HyY�l�,dn���P6ү��L��{{M���Ex�{�}M'��?��xq �߹� ���c>�Nt����"�Ɯ�T��r�)P�:@z���� ��τ2���@�cH���+}� K�_�LKF�W*����,��I�`��Ӆ>��u��c� �pI��k�)f�^B���NR�����':�+����w���~���������؛+�oU�k�T�K�3�9UR	��z��ƣu
C�f����
�C�ւ�b�����{�A*�M�nF�)9F:l��p~,X���I-խ�n}��R2.EM2�VN���^�yHuoy�%l�b�br�䒋��<-K|X�~_G�>���$�"�W��p~ζ��*���،�]�;��R]��4D��*	N�b\Xm6��'�h�|�j��Y*��zS@�s8|(��<ۊ�tӌ��/��\�D�
Ryd��l(Q�-���`�R
�J�cy��+/�L��0#B���b�*w�H��҆��4�e>��pe�� ���ll!�h0
9�E�~���9���5�:�@��f-���bt�>�&�H�(�Ř7�@�Xɉ���������A���e�i~��o}o�>��'4�X�/��r��#>Լ��I*�,!|��igN󗎦��)�!�ʜ�^�b>?�Q����ɥ\B]��8����|��O�eGj��#�9Ra�ŅqNN}iOXj��R`T�Gc �QYX��0L^�|�ρ,�C�>�_��߆�獽/��H��TX��>F��'򄞑��zdSn:KW�v���g�?#e�������U��f��3�Xcj���=H�
,�ʬg�����X� ���,^���%�i(t�I�٦P&5��P4-:�G�2�+�`֠g��Fc�ϐVZ�����OiQ��ҡ��qU�7i�%�X�7j�#cc�
eߙ"��i�~��e.�ҿ�5�e�Jq�F-�3�����YZZ��=��U��6ը�$ �-R����Y#��h���.&�&k���oZ��mP�����U���=��o~�W7o�O�W������w�@V��W�JnũH3�6�U�Y"P�`X�`K�3Ri����ۛ�fJw�x�10�h���`F���\lc�z���������H��}W�Il���+p4l���r'�Z�x��6W2���^�p���$y}��۫��H�fv�J?��3���`��>!��VߢQL��B?H)�7_����N��ng�ba.�p��[ġ����u�����~a 5�eD���J�/�B�e��'i��D �t�B/�{.��j�����k����e�ws����¶�ѡg_�=���������?�s' �3P���y�SM�'G���jӧ��j4�S�V#*F���yl>�id��=�Ց�����2�5`��JOnJ���+Đ-�y��<�)��D.�����(@x���2ΔGd}�2�	���6�y�X"��iwX%RLHŃ�(��?Ki(��,Bz��k��� +�23�����2�-����#Z����r������X��ٵ�X�P���2��h.�4��y�����7A:[�oF:��|�ۑ_��BnT%����W6�<s����~Ԕ����a C�w\��a��#� 1F`p矀!.h��Ye���`ͽtp�b���Jv�q�����ҽ�J�Y*T���n��5�?�\P�Ӝ�ԁ��5��>	" �ҁ��PM�T|�)���9�װ�l?�.��xS�{��j�� 1"��}_�(08��J�B�������S˚��i��d8UP԰�2�N����'��f��뎺����ٵ�3�����㴩}Y�9�P4�'d64\#��vk?dVZ^�s�o��� ?ovҵ�\��8@�_7-���ϦYS�K���9���(�$K�cÖ=[�u�C�&ǵ�?"5Jj
RTa1�hQT��HfT�	�T�CM�@3�Z�N�|d#�vV'1�ޱ�v���$��:ZOL-�W*�ɜ������L_���Hono��̔��S�q��۷�;����Á�؛��I��N��,=��r^)�g��H�`ե�<�\�Ա��Z�3p�����72^iD�S�cC��g���Q+�z_��a߯s�:/�-�����LDF��^�pu%-j��t�@k����1 =�JCev*l%L�dc"d�FnJ|����Qkc�M��2$=�ka�&��E�,�/JС��}�"R��՞.��k3����Wg�y���s$���n�YQ�~,�#�g��C4XA^��Ung�������������g�=	G�l��r��$�
է��#�3q�����p��~T0�Fjf#����XEc�ثD�j��~�U��"�}��� X���L����T�C��G�E��SPAm��'�j��S3�e��D[����f6#L��lv��`��ɍ�Ȇ��&�t�8<j�>��(�� �.�
��h�͞� W0cK�C)����dC�$�J�ڤʅ�����{x8�f�N��2Bާ�+"$3,�#�](R�
R^^#t:���1+'�r�� ��"@XY��Q�JT���#AV5T�=�j��bn�� �#�:���a��ۂ֮�(�D��j[�d�Hn�Ry�2+MB��_J�+&���PI&?d�u.�41i�K������eD�|MQ��GV�7*�;,��1a<�Q�Q$�o0ِkj ��lMy>`�&��� �O�w�W���c�b����]�o����[�_(�&� N���z�y�C���r~�˷�<�k#��Ð^F$����@����W�o���s��L�$N))��ܯc����UQ)��uF"�Ym%�9X ����؞��X��G�s`��N�;�¶j��j�[��/��<�0�t]�b�:�0E���D���3��I�.�p����P��h��!�s@����b$&�%�چH�R�f�?�X�1;ǳI�"��ȋױlyYI�dxQ��I��%?��V��̨&p��j��xι�q����"���oh�9>}�pO?��+}������l:��w�u�����'��e/�� �����:���,��}:��R/&��R�)P��k0����s�5-R"T`�u�)�y�8R��Z�Lv����,i}�����v�f+��#[�M�2&�،[���ͱ�BNm���Pa�/\&����]~鿛ջq�a�7̤_�w>�}����:к�mJ	IZ�O갯
��d���^�ER���K@#�>Fōcb.��x՚���>pc�
��`�V�^ނ�R�r}c�KY7�Y�vFY��hԀ��8��j32��>M�e���c�*�0{!w�^:��B&���|>������bn&�~���[�w�AEpH똕��:�c�d5`(%ճ���lAB�L"�_Y\�P������?�8Q�\>G�f��s�`��WY�Na5� Q�*���`���EP�I#r���oB�
kv�(y�͍eP����z�0<ܠ�\��B!����Q�bq<s5����I��'��E���s��T�n���]@�pԄ�����d����Ϸ��r|�7E�����L3|�-�V� �KX.���F-�oŽ���Fs2l\a.u<B��$3��~oV��cܳ����Ec_\�W[Z���l�-��֔�+�F@��O��CUdkx�aa
���S���ӡYE�Σ=XC�z�1�󃺌<v�.$�njY
��ZF9v�p�y���>���
�N�4�a�k��:�eEU���yq�/����S䛮Yt�l}dY(H8��ga��[6��������|�}Y*���0�"�s��_�
�Jڝ-��P��vnp��.qv�)M4��������k��^`%�S��v|nѧ=PB�y��gJ��%֣�jzcK���*�s��Tmz�?�>���˲�,��a�{���ب�^�\W�\�-1�����J�(�k(�0Jt�f?&�C�]�(ͲF�ߓi�B�9�ˤ̶\� �M��%y����6��)I��H
�EOh�Gb/d4z������{7��ñ��M��:��8����=}�xG,����ݻw��ի��/Vw���,){�
���ς#^�$�ok�X���Y�	OV�6;���}��wd�0aE�sf��/g%������d���YA_5�u#����k�Kt$W��� 3����7�Y, `���V��+h�MwU%����<�Y��>�`�q����{��}��~�xw���}�,z0lD���^�8X�g߳��6�������d����9&?>wo�3��֐DG�Fw��V�dXT�E�=xP�a��=�x�!F�=������<�`"��_���!]���./�o�Mو����|;�wf�'�5{f򴐕�le&�������3��{ �4�]��?�z�S<�d��g7(�1�٘ధ��3�N2b$`���f��L8�l��+*ٔyD��������zH ?��>��<�A���ES��X���{&}3���8�V] [�.�u�q2�ł2�� `�Af:}� ������`�9��7�?9M�1�p$�2r�a�CL1��F��X�J-*��\R�b��=�g�e���c����ClI��T��8�QEھs�>Y�^�_Id����D-8� ��dX>Ԕw���\>p�����q�M�"�g `"k#��6@f�
F��X�������:�~q����4�_����e�Ѯ쾮������	L���}���n����J��k���K6��TdL���a��l�`��s���ϰ�z�=E�ԧ�L��!����I�5h�ڞ>���)�)g��CN��nL��`]�a4�@0[ӵ�y��>}�cK�����u���E���u�����1�H�e^�o4+�g��O�I���� �(��\�t�/g��e���^DL��C{�d�Sj1GxV�#Ac�7�)) �_\�_�jd���cn������;�9�r�m��6���A׎y-�H�g{��A��ǴT)-<h>��E p�y�/+����a����� 8>�$�Y6���,Jc0��=����^��$�X�O�IS�c�`�g��#X�1�q�	;�Y@�g���
G��6e�N�lGK��1�e�2 S�������|~�L���8����-���Oo����&�������������J� �3���.�����cG��}�>AG��,���o�߆L�g�����`L��)o��Ck���^�3H�(��C�=C��}&�Ȉ�L2��T�5����{����>,��,#vgh�A������qXVlYr������>�����ڻ�3֕ɪl>��K/0;	���Wͤ�3�(���>�������xN{I��X�c�ſa  �%�����]�0,g��U����k��-�Ev�ٵN` �%v��L
6'����({�6�6�/L� �v�7�4�����x�$��/��t���f���Q��2> Hd�q�w;��@� �� X���B%k;=K%y>V�5Ʊ�vQ�{$33�Q�}� �h�9��r|�ϴ��W	b43m�L��/��~g-D��m�̀�0�,n`�u ��́�R�)�f�
wQ&(��0*9��53X%�hZ�W)���2��Q�q
������e'�ߖՍ�RĲ�i��\攲�4r�d�P��2��dhص�P��˃�em)�Ң��I\h�X;��f��-�ӫjڰ��h(.ݤ:}�:�8�9qN��?����k���s.\���282���{@5��ε���p�>��`;0�,͆7��ÓJ���<D��;���2�i6�K��o����� �)]��^ T�F�~d�,6}����:��ڗNIǥ)���Y`��v�L#�����Ĵ�������&��#��6�PDڄN�&�6lY����C��`���%딞�x����'���9�]��S�*����y
�'����Hd�p�!�mBh��� ��X��t�F=��ؿ��ٺjd�]�C-Β�U�~I���:;�G�����l
�|Oc����r"e�xYK�~1`�g�4���"���8�X���&����� 'p�*�udv�V���d\[��,�j��y�'���1���X�>?x�#x�ΚVެV�Y�����>S�pÐ���n>gk�-���p���L~��#�K�3�ʒ��$���X��?ҏ?����M�$A��k^ӟ�����;��I4�p��u�GR�=|.�Ѳ����r9�s{Gs��Y�f���~ֲYv����5��0~fc�T�v���/���:���_��<-[�6;�]�ΆZ>X�ˁ-���7�o?��X�����D~X���d��U�p'	�y��=��YX�#��_�T̸�O�B�3�LO	l)������+���ffv�Z&�i(�
�����Ĺq�tHp'�X�Y��v�~�6�.k�MĚE������G�@~w�=����	,0&mH����ZGX\�O��}F�>|���J��O�n�-������d��;��w����%�7�i��3P���zD��;��kُ*��t����-������齾��i�Ǐ��ֵ���Y�jJ�a>���@AO3Y 
{�xA[}���v~��P禯m���Ȋ6{E��TwD�2�eG��!$��1�008u=�9(pg�V�V��/��=4������#����������4E���IfʲX�Q����	��6
��cH3t:�;�
������-�Á��^�l��L�s���j������v��sgϟ���0Fk�tV�1js����6%ƶT9�$�:�E��׮��ߟ�-2�}�<n�2�?3�<s�F�� g��H�� h��a5H���ٝ2�㈧B�q�m�ߝ��w��n��֬�������4m�q@�6�K����� ̑��.�q�ı:XP�͍I�:�:��U�V���* ������^��ӽ���S=Y}�9�V�B�!���3{8�yi-DpF��9K��L�d'!��8?� c��@&�����sH���S�_(�ߧ��{ ���X'�Ԯ������v���VOa?�{E�۸^�F$_�V́�@˝򦎌�:�y R��*:�f��(�C��=� `�pk]3@
n'����V)lm��2�#P���s>���$��|{![`Ү����4�z �ή��u@s�&R ��9{�0ԑ��b���Y�A���uK�tZ��8\@2�����Z�<�t�\?���k�'UX���3�V�9���qb)��<�J�_�[�/�R��eeatm��K���hI>ꐭm��C��7��I �.��B�̓��v!l�܁a��h�j���lHaϝ+��3����8���RC�[�2����9��y��&���wg���`���ͤ�l��O^�.�(��g�r�B���~�q^ε�U���y^{��5/{��z� I�N�g��G>q����g��w� ��D����g�~�y9���Hp�^�g�;�<�Xw>�>32�Vwۚ����Z�_���V�2��0��h��`M��vaC���v�dR&�3�@x��a�'I��9M����^nA2sŉ�a�w���~>Tb�2��;.3�(��~M?c��p�\��+<��Le���ۼ�1�g�7��ƥF������=a�c���QB|>��#$dP��T���v�8|f������|5��d��Pܝ�{<�j$���|���_�/��ג�˹�����=�1�iy=���iH����������g��s����:(���Nx�Ͷ5�춦I��CNbl²##��,F@�f�/w������T��ڙ'�2m�hM�ƗQ,�?�d�m[��%�?27Άt������Zpѱ����X��Yw�F����.;9�JRF�\�@$>c����1u����E�Ƣ�S��bl�1o����k�ͤ����ۦ4ɀ1j?.��BL��{2 �8��fW��Ej��?���ϛ7���=���������d �ۆ<�ւX���p���1��h���2���#�u�%���|��K&���أH�,�<�_$1�����Q�=s��q��6j;�k]��/Q�>�_k�[%�#f���!�X�`A�O�aY�S'���M�H_��i8����ݰJ򗧬*����>�ufG��`�`��4
��Y�ܐS��QfeЀW),�h�8P\RH��5�����Ĕ��7�Z'����%1��Q	��Ϊ�{��e8�Y�Vp��,��Ӻ�t[�� "��c0�(Orp@������
턚�}̀F�~C$eO��Q{�8P�3������k�qNVݳ�8�6��ـ/�D5-�%�o�qsRГc��)Hn�/�����������I���� �r�WbP�� �� �
�W��$2lCM��[5�Ώ}|Ě���p"o���g$�כ�M�Ο7�j�� hג�͛5< MCF�^ k��FӺ?�6�?/�����������:A�р����B���mD���V/s�z2����jX�	WW�=K]��VM�Ŗ�X�
<������e6 �x�������z��@��B��B�а�O<H�|��č�	L��[� �vO�Z��G���}���Ϣ�U
��d]��Z���JFa�ڹ�E����z=],3󞶷��d��<[ق�)�%��ygR��~h{Rv��֪'��W�g�?4b}1��bӄ�}$"�B�	;��c��A���,��� чn������W�ִ�q%���m�y��8�~6�m�M'Q�S
Y�t��/��G����6��h�S\��3#lB�J˨�̬���q�岔P t6���<����VGM��y����-��_�H��^N�Z�!������׿%c#����_?̨����MCg��;X|y0}ѹ�{D�ݏjGpQ'�ߦ��e1�R96�l &4`����C��Y�	��,�l���e.a��!d���#X��Qa�6�/�2u��3[w�=}l��gK|1�y^2x�J�R&`���Ґ�\ٚ�Z6v��r~5���������A��v:��A��!~����i`O��>�L/�i#�l:|3�kt��d�gP7�N��}���r�]fv̍mt'�2>�F1U�U9���s\�7V��U��M��')�� �	Rt+�Z���هwu������*Xtm0��Y��5���@�,�$��|�R� 6�Qȸ�POP"�?�Ǟ��ٛ?[�g�^G����7��=,;$,^H��֎}�ݧ bޯq�Tɩ�k�C�9�v�9x��L=3�d#e�|?��X�)Y���s�p0������Ҝޗ��/�,�=���c�a��LdK��Y&7�R��)�';k�a`��7>Ypo�>�ŵ렰�
\v�v����e�� ���V&o�kw��?>�.��x{����/{ۚ�eo�7rҐk�@1��<pd�(��l�@x0�y̹H���l~��w �gd�q���ޒ"c&��L��,f��^_O�\��	o�z�g�����q�md���#�pʠ���~%�Um�%| �q��{pmA�u��9�0�������A�	� �h@��S��Y}�ͩ�������,��֩����-���$�AP�q���(E2)�e��_���}�WqϴV�Q= ������}3�Ӽ�N�$�D���S@Oӥ �������-��{jY]�u6n{L2�Y�{�g�e���������0�t�mf{�}�΃f;-�2�&�ڷ����1�l�yX��ϑ�D� ����͂x� EAV��ߟp�E�\�6�z1"�쏭ӝуd�2'7�Yf�uY����ڼ>,:@ڮgdIAa�r���m_\�.�}����l��*۾�<�D���3�`S��_��Q 7��bd�>��['fml�=�~V�e޵=�P����h��1�sP�E���E�q��Fw\����!�,����`�~?ptS7|����[������o�ŏi�v��oo>I��G����H?�O������pc*�ʉ��V��d�I�n��<���j�R�L�
��L�Bg冰���jf�vv�I���T8 4-q�8 0�3'=��� J;ke*$�9��֦E8uK�H�{�������	Tn_�-USð�A�D���7����<`��dz;/fP ʳJQ�ղ�����d�ߋh_����|4�2s� "Z�d0]fSG�X�7;�p&M�� �s�{s�1o��f0�9�BF�~_&�p
�̖����c� ���<��qNb!�(Q�?�k� K(�s���_F7(J=��k�9_����^�Y�A��>�������d؝Q��j}����p �{s�g�)�{��N���`�F�2�h6ޫ����Rݘk[��Y���[+��� P���T� S5���ܧ�9�1^��
f 8��Al��x�����S�`�)�Y[��f��k��$+in�����:�Q���L1�^ #	Щ��/!
�{�,���od)xUW�-���� �DKZ�\��m�:�1V�E�h�l�σA��_�5-�1G
��0�Z����]w^�z]�t���xm�@|8@�����~;�uv��}��v�J g����2a~���l��t��ㅀ���Xw܅�x�?Ab�̌I]�!�ln�c�.
tV�ӧ�G� �I���a_��n؜x����������1n/�a@2���m�?�;����3(ѣgDV�&ɖ��u���Ԝ!p����~�Y���9^������4��2ɂ�j�Q/~�6l���Aֹf�Z�Eֈ�Rg��։v>h�3�,��@���Y�|�؍��_����ž�#��d�H3�ȸm_���Lo(Z�帐k,(�(ݱL���胀 �[��V/�hDf&�QH�>��+���=�����;,Ve��J�qш ���9�����ϢM5�����1J ���/�geA=���/����q��H��oه���{�����W��n������m��5n����(�7�0"��fa2g���&��rd�J�%��i
�
�Cm3!#%���7��!<��� ������q�,�Ro��Ih��ӌ?�'GPw�B㐅�M!��v#�3eF,s C����A:�[F#���A�r���t/ˉ1VS���X����	��^����\&����Ӱ����j��:ۡ�����ցn5v�83)hY��c%���#9�ZL4nF9j{�as��o���7�`T�B�Bc��@���X ���:?��>.�>$#�)g�)N�hb�^,�{�XoWI�(�c߫fFp2���E|[� Y��l��8B�a ���>�:7HP����دX|\`��Ӽ�̙���Rϒn)+�hUD��<E��˸�`/:]�ra2���z �ؠ��"3b�)�|<��: �N��Ui�	c�3��Sf�F�b����]5n��#�F�� �-[;淉ђ3`���Ƴ�v�	��2�����I�O�g�Y�n{`C����d�2}�!�||^�iئ���z���0���X����Or]�w��t/�;`�"p�,���e7$EP��j�s��-��?�CH:��쳣f��� �}���<�6�r�D��Sm�ϙ��ImO!��� ��3��5%��K��5>��M�wI��-�_2�Oҙl������Tw��8 �d��3�\�,)jҨ��3��M��[i;�ǤϞ�8?_?��]:��$��Ɛ��F�i���ll�56�*dzE\����[e'bEsc]�t��,ɝ�7U,����9�`at�[�8@������e-�B+�I�"
b
%Q�۰��*o�ߐ��^�@@��׍ �g���/�M�|� �3�?׹H���/��X���ﲃ̵�Sd-%�\=Z���=2 ���#g��׌�{9��W�����P~���j��Q�k{�!9upU5�\�?�:��9�n� �,n;O�wX�����ؒF=��(��|�A��p�/�Pn�,�p=y�@�bJOR� [�iJ����g���y��J���MA��g�1v�T����H_31a��P2$��5���:�MJe���ʦu��ݳN��T@iY^��w�:H����?f��5P��fi���D���.��1 ��s-�|��氈�&���X~���l����b�&�+8���q�.A��t�8˟�B0W��陟I)ݖ��8�q.�2`�]��b"KF� ����I�W���&�~!#)�h��\��vF^�YV�ۭ"�8c�#��c�%�fA��{��ype�	����dޭ��{�ĩĢ����zN-p�D�1�b����cM�bOς�$�n�ϒ����}j������d�t́����)�~����9�D�%5Ӥ+�4����=�y��n`u8a傰,������!Δ�Fv�Á�݄�A��+��܍�rM�ϱ�w�{_��t��������X��xV��a��5�7;s��]k�2KR�%��TOsv��1R�f��(�/L���\+�tC*��Z�׶�X���x+wJ`���_��gn�1���5�h�����Ɠ�JA�`1�2{���e��������<���|>{'��y}�4l�@&A�5`�&ʹ���o��1�+k[�3?N��p�vr��=�ޣ���Y4��<��y�͇�b̩�����r���߇������d9�8��V2�C͍�!m�oE:��E�5��+��i�7���c�33���a�e�)�|{!�N`ڍ��|�Ϛ&���k�G�ˬSΚO4ZX��C���#ö>���
E`�'I��}�f`�1V�Y�9�S��E�A�QF�-�B��]dݳ�y'&M�f{w������)���$!u�NmHa9! �t6\�=��ᫍ����.#��p���<���H��ߪ?OU���o���c��1z�#[h��پ�fK��l �,������+��G��g0��-���\l��dǻW���b�D��_ $���Q]�,(yy�#DV'L{���q_�$06�˓����A� ��u�Z�wϽn[�0��R��]��>H���?0{����	����v!�0 P�ޯ������^%	csO�P)��
j�
�}�B4fZ���>?�.����"�?���v;��`i�P/fx�|��l�Ҽ>�1�b8��=�4���L5oPa�8��{ty�<�������5����S �4-�=6��u���Թ8��P�+�h-Km��6o����ȳ� ���2���#hM�[67�u����{�ӡ�j,䗕as�sڼdG2"�#Ic�A��桏�����P.@��@��CAe_�a�Z�Ns��]��f~�]D��\+�rGS��|��`��N%��c�9N!��$�m��ps4�h$�V���>ajp��J>Nd%�s�dv-����2� ��S'�{	r�2����O;�wJ��l�٣����&i4|ks2��k�Q���|�=��e��:��/@P��k|�U.y��)	����Wx/����T
��n�&n�P�L�+���s���Y�.�Ȥ��6hX���[f� ���'�"���̊��.3��- C��̌��lHQ���y
vNz���+�5�7m��O+c�?�0<��H�_�x[Z[Ԉ(���Ե0�X���}*�A�� d�.DǓ��t��:�.�dTcC�<:4A��d!huOR�t�ۂ�m�I����s<N���3��H.����;�ct L[:F95d3FVA�?4�mԵ}I���L]`���e_�:i�����)e����,��O�)�˙YI1��]�P9.��ͬ��������j��MX&fʳ��y&�I�Z����N$����Ug�t~���7�� �� �h2T�oG7�Yz���a�,������؍z���رo�@������$�`�^rY�YZ�O�q�N������2]^���c��C�|3e$qzxZb�fP%K�@�$N�}�#ٹ\���fޫ��f�l )�P��o�ĉ#��\z��@Į�{I4� |Jd��u��}{?¡�%��f��v%�l���7��i#�w�� �5P(0��>�:�f"�Y2������1�sP� �`�]�H&U�g��؃ �}�i�H��۞8m�����|sҋ�%�1��e;�u���"�^$��}q�Z�>�;Oy�R'��l�C��8�hCҕ� 3�l�`��ݤ�݁�u��jo`�Uq�� �����yl��<����ŐAI�� �T��q*� �[��k��; �Bѻ���C�q���j�efM��*�*�$ںm�O?2�H� �`��T(5�z?l7����r�q�uW<A��;�9�$��D�(+h���� �wq��U�~܃��
�fɠ;�C��:�f+�?�����k�q�u�����KV#��fsn��݂�-�_�*gC��ף+LL�u�/���;�C6���0r�6�@8R=��k��<�hsV�b�݊���RfZ��A����i��=+����T��@7�s9e㷴����T�K���{M ֆ:����54h�`EVN˰�%'�r\�}Ee�gH��J?s�P%�o��ߩ�4" �c�X	{�d������_+�3�k7w�^�5���m�j�QeTv�5Dۯ�9�돡}�Yu]�F#�v"��5�`���_eQb���;�/���k���@�5�FV��ư_NH0�|lh������a�;�*�����'9~'�b�
���L��A	��E(��iĀ ����ut��D�@�oZ�g�Y�tߧ��	��b<q��a�Х����&��X��(����v.{�{'�S�Q��<�㡝]G�Gz]{X;�r�7g���F��<�����l��}填��[��E�L��H���~�(7"O��g��o��˵�_�fNC���oC��Y��<>�������	`�z�jI:����z�w;�"���=Q�%Fĺ8Bg���Z<>��A��tJ�b<|ܿ���V�T���!9S+��LR���N�1���ҩ���X=j)�M��E�ް�<��
w$m!p�}��2eH�����4Of�j�٭P�S��Y�\��/$Z����0�<���fV�wӄ��_��]�o��$ݜf���9Z�ɉ08����G��-y�ݘ�cH+l��Q0��(|�÷��1��=��������-��u[�2��qtx+j�2bP�JL�\�RcѠO�����fy�h3����ʂ\���o??���%������k'j�,Y�)�� p�N)2'��|��
Ճ�%�f[`lY��n�53�F^_��O���:�(�������Y��V<cP'۠��g4��M'��r�mc.��2���0����SAV�K���w?Qo�Z�Q���-�-#�(WDP_dAU��!��,${���o�٫�3����/7�8 x�
����gMx��KTvd�s��| 6[��&�m�2aFlZ�È��FDyC���l��%56�#�P�
6�t6"9I� Z<L� R���ϴ�����,Ka�@���p����p���/�Œ��آ�]�����u�si4y0�h����3�[w?�σk����v����ȍh3n������75P��;� 2�	l�Z�sj�7f�l�X�ۺ��C��M�c�V*ز"��`��@��e��s��7���Pn��� �H���j51d1��$w�������] Qpݬ����,��֊̢Y`�aǗؙh%�(����je�t��e�FP���&cN����J��A��V6���n�%�z'��J0��,b�ʵ#�_���m��l;�� ��QC���"�m�ڂ��}���o�>�U+�g�z[���fj�4�|���Gcɐ᧐9�IHL�d�����!�L��v��#A$_ٳg�gx8�D�Ğ�ւ�~:��,���H i+��X���{vxXc�W�2�M�T�jX����^�U]#�t6���cC��~�{W�~��`��H[�kq[hG�Z��82�0�&	"R�������S|^q����8qX2�b�&AvHF���}%tGB#<u!�vu�m2�YF6�]HIG<���E��/�v�cR��U��ԟJʁm.O:�������;���Oip��c��p�(P����CA��<0�{���e�XoĚ%�/l+_�J�S˵2���H㤭F��F$SF)�nN���Y�#'�����R����f��z��A�s�lHmX[a�³?��i*���
�� ��@�hJ�Sؗ`��d���W�-���*��L�Bd�w1�9�,�kР�[����.E���C�V���Ԃ[��m6����dg�����%ż婭7Z8�?�c�Q��}�5~[F���,ey��Νs��~{M�%}~,鱭I���fq�fK�������A ż��c	Ш�%r8n�لCu����`��y/[=���EY�Uu>��rIjn��-y��P.����A�k��g��K��{ٷ=֝��s�:/"f��mԌ�i��w8�l�i'۝pQ�77O���` ։���y�)��,` �Yu�/�wR����$\��7w��b.��vW���)+���@�����^_٨b���#{t�'�pm((s�ǘ��|~b���ܢɊ~n�y�m?𲫓�u�L.7ּ�.�j���F�2$���-I^�w�n��N� �s�l�fl�GÁ�%,����Õ1v�����ϫ���ϻ_�l��o�8��#-�׆���ٌuYY���+Y�$�/&` ���^i���Z6a=Q��~ν�UBpF�ۋ)w��9
[�7d�17�q�_�"@ݭ:�dÚ��ԃ�vy�R"��u��'��!�Й`��؀H�!�*���ױ{S���$���]Y�ȩ�4�	��f����O��F�@�3-{�hתg����vb���^�S��I%�G-��ܯYc�\���I�//�p\7�͵ZA�s���Q��b�NID��5��y���YX��Ȧ�V&�	)rʨW�yde�=I�����-H�����\�w��3����,��l�n�����{���M1�l맆�lh-p�|n�䥉�R�8j��g2���u�^�����H���1<���k�}`��Z/�_{A��d�u\`����d�˙��6�����Ć��FS,���-���̔Xg6B'�c-pAp1g��'t��3��I��'c�P �44�2����uT
�?	���25�����E�R�N��,��h(ceْ[c��,�N�����m��u|�� M�J����h�����M`c<�������x=�����}o�
�b���QF��:��h
 F�i�����#+`�9ǹ��W�/ms��(���8n�(���nF��2[��r��X���zs��c��E]	uߺW]cy`2>z	��3O-t���$����E��
f�~nI�b�ͺ�����	��&���B��`	i����-xH�!�T�S@��SmQ�Q2��_j��٤`�z�`#��pS������At ����@�w��j1l�,j�����c��FM�k������>���j�2�)�Q�-"d�>����@��1dvfk���$aYu��R�긌1;t��&�t�y��!9�W���/@F�5��()��?7����S4ZZj�q��{!�R���*ӳ������O�A,@M� k� �h�=�M���tU��FG��7��ݱ�&���Z�@|�5��O����e���,l��Mk�b �,a�H��� ������o9�T#V8lNk<d�GMm�
�%����@��:��l��t��������l�,
"�`{+S]��#�k&�gu�侲���_q�ѡ�KTy���_�����xp�]3��Qy���5Z��@�$43B�I�,��� �.�i&�� �$�� ���T�A�ƾf	����l.LZZ��m�ӹ�i�ed|m�X�,�%u�h�l�w6���s���,�e��t�'a���|�+��Uh�O��	�'�PO���z��> ���՜��X���p�K�L��ΥK�,��7H������_(��+���0u$�Ϙ�?�:�Raoa	�Ov���j�2�Q~1�٭X���]�ި�|���v}S�"�o����W6�S��M��$�6Cu�<�K�ȏ������=�IY�J5UAL��0����"��zg���~���r�    IEND�B`�PK   �X��"�IY eY /   images/63ea08ea-b384-44c2-906e-17d581481095.png��e\�-��{p[ ��[ �\	������%��,w����^������ef��7�5]]uΩ�0%i4d"d  �&+#� @�  �lD���������@��!  �J��0<1@� јUw���� �~��A�,炳�W9���O䧂;>���o�~������*�j5#O��y��Zm���|)�i��;��׷�9>�^r����y?������|�
\=����d��ִ�ԇ��Ȍ�l Ix~���6�(``i��@��e�4b�-��\�N��wBS����"D�^���_ku�a�H�c��ΟK�_�wYC�Ѻp���8��& I���5�aǵ{�޴���b��l�/����䍚Ԋ��ޒ�aÖ�¨�w��Ce�R���r�AüE�Wq�������D�L�����mImkI���w����c�}m��à��r��?�;�{~��IRB�'uϔ��4�7��M��+G箷d^&Y;����_&C�'�Vk�4�f��o[q�(E�����5j#��a���ލoI�����jȓJ�	W���k���$F��v�մ���5R魍�˝�\�M�N��VK��+�>��18���Uw�۵�d�f�O�_���<.��k˭G��9�[���w�U�4�ԲM�py��A}�U
?xP��rP�(;p�-J#��銖 �ixLD#=A3~�|C4���j�*!Ǆ#��y���7��v�K�#��G��\���� �4���B�8�A,����R��@�	�<Sj���qW�|���)6��
G�fW�&gL���-/��-M�D4���"�(��@�u�hD#B,�2��F~�-Mo��×}j���n�e��F�
9�y��rPL�"@�*4vO����1�̲)��;9v<��s%�M�|�.�.f�*b��j3���al͋�58�Խh���L.���*�����Q9�S������-�l�t���D��6���.�A,6�����z�_X >j!B��!�Vxܛ�&A��V�ˋ�*V��~U��G��1q��9l�Q�"6.��Xg��_��;�6Ԛ|Jȉ��m�ұ��;�N^?<n�>��&sb���-�����������Iչ?S�=]�V�y�w6�ԍ��(e�d���`��6^%Wo(�]���k�V�E�����E����ңm?��-û#\ٸ �>�}�����q�����/}WxA>ҏQ�~���$9v7��4����D�h{{P�%v�ۿ������o�-k�_�8����<f�h����̶�(}܁ ��$-��#�S/�.w\�way��O�^��Bl���[O=N]��c��?��H�`GͿ�����d�b_m����J3�V�_����1O�%���O��:]>kj����)��	6� 9��h�~�,�~���Խ�q��|m�̙='�T?�-"����dV�-��M�G��,�'�8׊<
-����^�%�	<�V����J��׿�gO������������/r��[U����8�$�cLf{�兒���_$]G@�H:�Gm5\ݜ���
�&*9Ǿݟ��r6�rKu�TNڤ�>�%����jA�\:�������R��Ф�|F��ᝥtx�G0fAo 8�M�����僰_�F��s_�b�Q.�'X-��
������/����E&�,�;��ʀ|����S�ѹٗm��&�I��d�kE{ι%�����*S�|��: �a��O@I�s�s��Sҵv�j��b����O縉�s�\�z���C[�%׊���kL�����������|�%����B��O���d���˰d4�:���⢎R�e�������.�[A"���e��?
��
L��Z�?�{8�����l��%��R<e-�Bu�0���z`~�]b^�E�����vhE��{9�m��y�nϩ%�-���N��y�}C���&�T��ӍBw�*��ȇ�`2�6&H�+Z� y�á����y�"^��e_z����s*k͖��U�5����G'4�NP���L�;�����<֯o������q��W�"Գ�l`O`�G��q�b.����9b�K�zx�]��r��a�V��}Z�z�Զ�ZC_$����f6n�GZa:�9jQ�	�$[�GE}��[�������� f��MRӃ_c?��y`�C� ���/�3�2eg'�Z^���mob�xH��E�WD��3Y��y'�l$1�Z�h�m�4F3G��RQ���OO��u���Y��n/Pl��A�X_H�]�m�����>��?��/@����Z-3P�%�̯uRk�T�H�����P8y`���Ca�[�ZP^~TJ궴�Ǥ}aY��D<o�H���t�nr#1�Q���'�q FRۍ���QX}.>'�g��R��h�)�-^�739��'6_M��
����tjez��`ԡQc 
H)Ň`�k�<�� a��On�D�,������o�^܊8�㈃�#��b��a�k@cї����S������]ZQ�qYڬ�h�u��|�}�~�@[��}iފ,���V�q<�D9L�B�y��D`�#:j�͊�@0���m�ș�.��K�����z1���� z�m��n�b��\�� !_P���aM�)6�!X�pJ�.����{��3n���/ʲE�J�Y��W�_�L�d�h��,O����=��@E��2��h�2{��AקL��V��bf�Z�?��Y�����\�;;J�lw�\�<\ќ�L�+z���0 َ��)��$�S?�n`��lW��m��M���@�g�����f��o;J�6��������5X��뻈���t{�v�p�B��Ll��+7lkD�\O.E?�6��|�a5�dZK������]��@}���EI��/�9qk��N@o�Y$
es��I�+F�����U4K��-	��c�w���~�X�����cM��:��ή
v^>�j"��<�Y:�������l��5,cf-`b��ǭԯk����)ÎM�dZ�F*-{�X@ɹ�Vju�Gg��"˓DU��W�0����k���Y���.������Be�����?:T�O�VI���OOO��������U��.�W�q//
�uu��WTD�t�S�	�����|�eH�s-����/�4��ٽ�V�y����6��c����e�&qt]���xy�%yZN����S��`ՙRC�O�ޟ�ó�C�3���ܾ�Z�Vepۢ�q�"��<RYnUt�ν�v7��u�x.����m�Ε����W;�Ț\���%L�����몫I��z�"�ك�77��(F04p}��Z���}?�ՖX�d��mɉ�*�:�����*�:leאs	�up�5����R��/q��WZ�&��^�\SYUQ!S�h۩SRe=�ۣ�޿���Ȱg��Fۻ�~���l����T��.�5���̧M�v�msZc���7ww�G�Xb�J�r�G��IwK��l �Ӯ�3��('c��F�Q<��(^�ۣ��y��Fk�U�۔�jy�� �X�^��xb���h��"�|������b���9�s����n�fT~yu�U)��5�?(�\}�����RÞo�#m\T����c2�ƟN]ݱC�	��Y7������y������� �
S��RL0
TL!>��6�ɱ�0w�J@l3�in�u>U�4	�A"rwʗ�	�P���ԙ-d��T��/��$|��	��k_>0����_��'�u�'�ؐaZ
Y�ۧ{�3�f��O�M,�k�����8??��Uk����~�gd<z�,E�:�Z������~kV�����%�k�>[��F���¶09JS�@��&W��A����x�2��=z���8�*��8<�Z����7�C��J��%oE0$v!?N�܆���"DtxVw�t��V\�~�z�׿u�����+6|��=Zq��P^\K����>30Q
��F��ۭ��7�I���da-:VG��e-�˒�kv��,��B���}	<�'m�`������)�땏�y^}�:�i�>��?���Z���w�'��#�T7��tT.'�m�O�i������~�Ͽ���ۧ�~ ��2���b �E4��?ؤ���[$�>��#|�d C�w��P K�$��*�s��7�	�._�®��:�0Q�8ax����D�j�*T������!�Ժ��������6�]EE{W���mH��Q 8��F;!�V
�dv�?U��T(�����z���:��3B�d�G5�==I���7j��zK����/�p[��uJj�z��^��d��XdRe�m���J@��a$�7b.�ϑ�!��%/W`Nd��B~]Vշȹp `�����~�`"���)�_O���MF肠�,k�h�a��x`������N�"�+�bΩ
pQ�KR<բ�<��o/��SF���J�X��4-ɍ[�{��A�]?V�0���H����i�4��|����)pY��Q�"703~��\>�/�\NI`d=oa�-OO�F8��t��D�9�<�'S��܆��8y��=�=f�#hy�|M�뮁��k���R�VL7���`lM���}2��!=�n�?��ΜH�繁���2uf�o����$��/eJ�n�!z,v�G0nok� $�ew�c�5#���ikˉ���Ŵ-3I�ihR�h릢Q���%�3`"�B�DD[������a�|T�%r������+W��Wօc@�����8z�N�G��G�**ܡ��.�'��-ϛ�(���d���
�Oo�0�����k��+��8*��e4��nZ	r��a-�T��������{?��z�o�a!��sB`+�|�Z�pů��r�1(*�2n���N�}�W������_�R�q,V���,�R���ItzȠ���]��0Y�*S���hBw�/��|�*sn����y�C����B:�Ym.Ϣ��o�!
MLA鉨�CՆ�L�� X��pۚ �F`�w��06������_�Z:FI�Y謨v�_Y�c��n1��ϡб}b�GĴQ[��~����^���)S����|��/:������q]:� 7*eFD���������<�r
�����v��u[=]hu>X�]i��[���R�q�z�C�����l�����J�<v9��h���@��q��r:���'0mN��ʯq���أL�K��Y)09&G��wd��8�Uw늳0��!bC����)BT+|��u);[�j��1`� ��&tNW�I��62΀��@WEV܈'�d:�b�xּS�$`y�������B�QBj���J�Ť�T�Ч>A}��Ak��>����7,,h£CIg��	���³_��R�06���"�WO�"Ʉ' �$A}��	���\�p��[o	deeƫ�<	W`���##FDM����C���ȏ������wS��s}��Y���z�7��i6g&AYd�	l;�����S)���_��2Ca@��O�Y?���ɸ��ƫ��r��+�)�|��m�~��JG���Ƴ#8�c�{F��h�rܯ��c8�#�k挒�t��$0b\�@�v�����8
.݃�Xwā$��ǋϵ�3�.�L�3�|���]\h���C�(9@�N��n��q��X=d��&�;:��F�V1��u��,��rB�/1�t߾wm����U�(�}��$-坴�jw�pk�Q�J��jl�o��Viяk��$Fxm�M�]�H������r�}Y��oP�G���
��iEjof��'U���[����6¤
ڻ/ (.���W�0X��x����4�	$�IH0��o:Deკ�t��u��%�o+�ԣf��d�(���X+�ˤ��~�<�n�q$?���|��(��^s����Ӳ^�}��o�=��^5v>A�t���F� ���EC� R	���+SZ�"��+�_H�%͢g�@Y�����G�:5�g9�:���k@k��G�:K��.檡��'p���(�pj38辕��J��o�+������������>8�: ���n��=��<�O]�L��}��i0��`~��7���؞�/����چxp�?Zਔ:���� ih+��0I��R@��5K������yɪ]{�3<�f�:KN-s�U������5�r�P���'��ŸhK�i�x�ҹd�>���U�R�g�1�qۦ�i���s����P=�e���c�V�kO�읤FU�w�@�Cڂ�;���!��> ��P��'�"��I�@�<3�JyJ�Q0e!�3��$HD�$L�� ����Y�����(a1���;�Yn�&�A<��^?��]ݦ��,��L=�5�|9ЂOS�#L~АQ%��~-d������C��5F80�`���a끏��핎�W �R�v;��n�^EN�s���Z�����l"L9�9 �,��cWrw]�yk��i���27/��{�H�s�ְ��8_��
1�?+>�Xu����A{s\<��m�|RJShQ2����<ؾ4���
�7A�
���Q���A�YX�P5��Q8���/@Ze___Q&Ǿ��R�C^���RU}�]I�o~ïUC8�p[��"��Rə��N��;8І�郋�,��Sռ{�,��^_D-��$�FU��2�>�����UQ$x�]@�Դ��V��v��bU��#O2�o�����?�j���Q�.$C��l�u��c��7e�|�9�:ϯK���S���AY��
a ȧ�k�Q,c���^�_6��D�����D�f���UPqX`!��1��!jF��yd�T�>�������l1�xy~�~�ە��.�."!��A�ޮ�5�pG�ؒc�7&<��1v���#�4˳�����~_��!��������U@��yT���c��K��,�s� �|�0�{���ֺ���~B?[ȬiS��cҾ��{���� ���75#Ŕ�Ւ�h��HOq8ڴ�Y���5�5?A��xS+�5�1��<���9�O�gW����r]'E#x���c͡a֨����Y��E$�;L��e����eꙛ|��L�p�/���F�Ij��ڝY����d���(>ٖ�����(���3�?C��?cr�2p��H�m.v_���7�y.[w�����˺���gw4�u��������W�a�Tq~�`���y�%�0��	l��5d�����Ǆv�/�f+,�>vf�i�BW�!�Φ��V����@pK����a����P���(�h�c��,��A�L�)�mε��<nKU��>��訍�(�3�=Dp��Z�F����z>K��0�Ц��L ��Q���-WCug�B�y ��rt��j�bmqh�#��U�h�*�oo7�������mΣ�G��qJ�u:�N��v�L2��	6{���il���:�t�?�c&LS�
#(���9�׮:R+�j� "푯��&s��2�O{#�}g
e�|�36^�ls��ը6&Xk��"[��Ğ�]@��C_(��M!#l���L:N:��I�զv+��9sSMwޮJ>�k@�"4nE����]���4�f�Z�&og~����;��!J�W�خ�|��[��@ ����+F�����nJ��`�<�a�rm�3 ��J�ޮ��>J
��)$y�a�ǩ�s����ؤѭ_�Y׼ţ��b����S�VMlU��ʲֳ#Y��|�$�d�n��bj>�VS��K� #�?����%N��+�����)V+$�R�5������]�������,�W{������G�"��u~�����5��*񐲡���=b��j;N�:�#$	��֋�G��!!�9�Z�Y n�`ic$�r�܉��p�D���(������G|�6�KJI��edI�^A�4�|�i2������jI6��;���c4z�3>Q��+s�/��Q>�a]����T��FT��+$���F����&m�1�U���ٯ^g����Tc0s.�۹[���X���}[̹�@=�/�^L�.�sW� q� ���6�2�P b�|�������`����{�j��2L����T1���c��ߞ"��n��}��,��Q�b����UC�A���z�H� ֊����me#��	����P�Χ��E���
��A��t6e\L��h��:h�Ԅ�P���N 	�$��#z(�m,X��ͤ��J����x>�
%���K1z�H����~`1����=�Kȼ?����?-r"��x���En���8'EG�Z�������{�K,�6����aƨ���3ڥ���6~�����T��rT1
s���l��6)��I�q,���*Ċ�WZ�$����~�T@�ڷTs���~�X�k+���`S4�kϚo #I;r�iV�~ޕa�����
FàG�c_\j��F�!�_�Wt�U�1��c�?����KZ��ᴦ�u�p�9�r�f}/��d�3�$����J%����e�+��?tE��V膇����x�a �@*ꈌ�R^C��ݖ���h�։u�����;��c
]5ARD@!��<����u��<Py�m�u�ά@,a�X9�7�������w�E�?��xf�\��1?��vX�P�V=�K�܍�kN���Ӄ0���L��.�1j"���lvJc˖�"�%X�>�~;3�f>��.�+��Q��5���u�h�ӷ���PL��g\F�L�e�Q#'}�界ru��X�jn�Tac=hw�o��g�Ii�
ì�L���ўK0�$@o�������X�#�K
����e���C�B�=�H�M�ύ~A���ym�b0o��*�i�(�K�1ӊ��������U�/~ͼ8�/�?ԓv��Rם�u���w!O��*ΝM��p��⭮�靔���?�Iq��N��\Mŧ������6�O��q�a������`�|��:��tVi@�+�HI �s�)�˘F�{2
$�lE��Q1�\\}�e[ۢsv�N�ug,��(�T��
�i�ޯ��Z8"���G�9�������m� ���-�g����llV>��U��E��x4����Aq37��D~P�پc��^��v�֦�\��u�`"�>�Ľ67�o	�j>��t�[0⃡�d����8'_F2���*o��B'��npX���eٝ���|b���l�7O����ҰY��3���e\����aԗ��<' �}�$>�9�Ͱ�����Ԍ��FDD.I���jo���B`�ˁ!|������^F/#`O��.f�LCwr��t�#�Ӄ���O���Yq�vK�crI��}���l�:���NEv6�,M�ǻ���*��fb}�0L����V�	^���yu�&���g�!����������$	��Ws��|�Q��|���p��[E�@X����?6�c��3����Z�������nO�/4w�$.�d��ג�p�9�⩛5�"�4apo�ఔ`�	4�cJm���?==�(��%R��ҾO���k� w$n{^�H��c�R}�Ȅy�9�5��j�UBs'/Čb�\-}��|���ً�*Ϛڱ�y
8�06��,;�EW���d�[�~�����.����b��^��b��{�;�X9���d;ޝ�V#�(���UxF�C�N�ǂH��ʵ�o����\���2+��ջj����|�닞¬Ь#�D6<��i����b�ϋ��e~fWsQ��K��\3KK�j��m�04�H�	���].U�v�m_��JK����b9#dPi��9CԴ�^_E��Q�ժ^���tdG�w�hp]��bs�lѦBU��)��>�C:��U�;Ξ�YWw���گC�phёO�ˋ�~�(+O"���誫�|�!�+�p��y�GyT��/����^u�l���l8��Q�˓������{�C��\$�M����`,3l���	��Ήv�엻m��P��KE��*�h�*���`�����(j��)(�kK��kMc�-�<�_�c����F�e�-�;�E��N��Hٷ�#K./����7�����!g� T豟��]�4���m.���%������֐}/���=��*Y~q�<�Xu���gE�Bu���(C���Y+!o��������sSz���+��a��ٲx;,�@3G�r��^{\u7��n�4��""X����V�pd3Ič�!r0p�+S�綘�<'w�7/RP�St#9(^XX�8�7��b��k��naZ���^�ZKa�
�hhEA����'����J��`pB;�B�\FY@�����翄c��s�۔ظ�p1����Y�&�o]\��h�6K_�S&ĸ����Þ�� �xqE��z���l>mҵ��q����P�������+++�J��7��ө�j�}-,n4~k��N�m�d[cC���3>U����Ku�]����L ���h�\���jݾ��i�E�+�6�7�dH�=���#tJϽ4�yL,X�N��|�K0a�1)F��ql���M#Q�YhsԨbkC�F����t�W�l~�UM뺡�f������F���ea�m�Ŕ(�F�g�]�7F[q`(5%b�]0Ůu�C���At}��Ԅ�BмM `$���O,��R�n��)<��F�^��1BWC���'���v�Ĳ/�W[��~k�ʬ9�Ԯp��3e)-%�Uh">�]�!���|e�J/w�`��%��*��p���g>�j;�!%M)̄uh#3ޡT��1VF}�ko�@��-���w��w�$�d�|�xS۾Z�QJ�B2�0P_�`�U����g�Np�����7b��7��y]#���/�4wޭ%�(�_O6�rs�Fr�o�ttN|�%�f�קb-#_��r�����%.��r��Mg�~�G8��)�ܒR��V1��{cҤ$�\G��ߛt��رg����f��%R��*J�[�fY�i�`�A3ԤN�f�
k���N7�ߣ�@�]&�-�^ɮ����^�ֲO(/��	���"�%��y�:�6����C�v+��k�wȴ�3��iM�������b��S�*���*<�j��b��V[\\��-������#[k�o�$%�@�����;�Y���ş��N�Yd��/��l��@�@��ގ0N�>3̻@m�ņ!����]�֐9C����B�P�7��C)�+��&��p�l=�\��:B��p��/�|���[_l]{6��L�B�C����W���?0�eWz�\t��8�/]�eC�t$Y�cz�����D���7sUo��|��:�2��@2��������wל@�1'ܯ$lK�����4�$`ocߌ�!6�di����"�E,C��s����^�@�;�m=�~b9��3�w�i�)m�#3�Nu@�����u@N��V�KcO{��+�<��#|�p��ܱm�%�~�Q��.9ܑE{=ɽvq��4��ց�#�P�X����vaF�u8�����J;�Mk{YDȕ�{��P�JC���L SX0�P��`�����G\4.���A��U)7(�9c~Vy5�h�4�+�'��M9ZWz��Ԍ���A_�����*�6�a�$Jj�� ߘv��.�����`]�Ѐ<k�J�������V@v8��X�c9���`M'���A=��ں`BKH�e/`�d�]0k�����S�hZr���`�����R%ȁg���B��Tl�$n�������K�@�rߍ�n�Y�����ɶ0�LA�I~pe^�Bw�I�ZG'�'�0H0��:�N5�u�Jh	�Ĩ��5�c3���M��lL��=�[�MY`�����q���gDu��p�A1��:S��2�|"z�4ݦ���ɘ/��,�Ҩ4�%t���S�$�LO�Q>B3�NL��2_;U����=7֞������&/���i9U�a�x������"8�Foc�caEޠ�i�
X�a�v�x�]����O�5g~1�i�+�zk����FD��r�qD����p3���i^��N����� �����&�S��[n�S5�H�5ĒJ;+�"� ��g�����B��荋x�?��J�bC׋P�+�o�#c]!n"\
Kɚ�T�
�6�i�3��p�\}�פ�a���O��Ltg�D���-ͨ��w�,���2�W���P~j��$�N�vsu�PpN▹�PO-l(G�Ƿ��r��mQf�a�=]C��_$4&1�� �Dܨ�(qqѸ~�)��:0���E$��ZK�����|LL�}&@ս<?����+���?��A�|
Ke�):�O�c7_ ƹ�x;��4�� �BĞ�t��?���]M]�����/ bs��O8�����5�P���J��GnifY!���j!&"zr�&�5�<=�Ԃ�
�ISx������pa&�G������
uGG��	Zv�����ȳ�*�^��RB�Z�.�j�D��f�n	F!1�֝�3e���@VK�Dێ�Bl �@��^h�ց	��fw�bJ�4.��晌p����ٷr4jm�{��('�'�7���@��G°��Z��q+ip����%����Lm^� 1��ZDQO$"/���(΂��j�.d%@�aW���8��Y��v.��Kc�����>.�g�ܐ=�ְ�����&��5\k�
��}^�szB�9�P�UK��t4�s�����c8xg���RX̰�3X~���o�\[��ԶT�v����y�t�y��;�5�1b(G(�mB��K�7x�c/�X����ʎUP�++%l�|�NҨH8َ/Aǫ��~��e��H�,�A�׽�i�#J1�C$2�,$+�Q�@������T':V����$R�tZ����yђ,���Ԟԟ���|�c������'���F�{�wk���7�#�5 ���Gb3����i�DbwG��v_��~FI��TlߜA#�`ґ	��A�IҎ�3���O(��]'!p���g� "U�`1\�P��eu�	m�F�~�ʨ�;Z��vDG��B�޳"�ˀ ����E��4�_��U1�o~��65���{u�E��]�8�HD~��<�����oGycm�2�?9�!B�k����%6�,,h���8�?L�ZB9��ؽ�z�I����|0�j~��ށ:�TjR2ѽwR ��(��bր6�X��TD^;�Q S�V�i�V���~��l	�C�@�>~��Ȁ�қ�uDo:M��V��+�SKL��a��l�hQ9狅<��x�)8��d3�XXrhY�G���%��[֢�G�F���"�t�ON��)�S�5sX��db컗�������|��ɔ�����59�ސ�b�HJ�4�*Ej<���r��:���:��Vr�)F~i��q\u�F+��s�_�/�rN��U���K2'��2��������.�N�"���;��U�
%��T��v,�}�i&)n[�o7%��2A����r���#�P#���}h��4�%���'��P)��)p��@�Ts#�^8�st^��Z�����)�CE_u�J��E?�+cDTJc�QO4
�-����w��,T�2�;��R<���;W��/o����"�e��Ʉ?=t� '�SH:�O1��pjK��L��P�ۣ	eCI2�2��w�$�6â�T�H�cB��O�j���X�>���S����f0���sh���7���	��;���(5���?���/���3�ny��_σ,��4��
���׻eN)��3�6����n��ARw�����H�I�w� V?�4qJGI���SZ�T���������m�O�J����W{���<�+�<�C�?t�Z�AIA�3� 6�����PRb��C��j�W3� կ"a[}�lLKl75�'?��Y��u7w���;�}m��fy_��i�P��3AwH��/��Fw����18��C/zyX�u� � ��c�@���¼�E��ge_)�5���>�@ �a�%?��<��!�8	ikcc�Ņ�_Z�V*���:c��@�އ�4�A�D��%-!U`G	Zw���Y�I����8Y���3���p���!�,�T��獛�>�z�R��0��D���FN�����l>GJ�_��?�n
�kY
�5��|O-)~���!�7}C��HD��0��q1>��I�+�!�Yl����,���LMƭ��8�Bq�Lxb�L����]ꐕφ���|q��'��S{�c�P�׿�����EEu���8v�z�Ν�9�����Lς�_����ȝ7W(nC�z�����.�� �8l`
����yw�4�2k�P�NQQq,��
�����#-G����� �[�3���\�Ԋ�/2����c��gp�>�V����]@�
A�#A	�����^g�Y�-���F�Ʒ���GrlyC�!6���U_��`���Mafm:3��*o�܁����v��q8�����yVV35�}}��Wڢ]���S�����P�x0
r����~�ҍٔ���+� `K=�x�[p���Bz]�x�@�d�V �! �M�	��X���n͈i���A���E6�-�a"pH���cGB���1���L (�@
DS�.��t�Bt��5u������h�ll@z��;�h�����d�Z�_Ƅ��0�t��?ȁIWQ0�l�a�J���.�*�%���Hl0q���
�����!�Uua��S\��сDJ�����	?�&
a��t��n�No�y�<"$) �&��~	�.�ͧ:�	�f,�]�旇�Ů;�豶���z˸O�*���EG���?m����Pb���ƣz��<�� w=�BҒڀj��c#u{H�
��K��(Ky�)�6{(ߖl6dO1K(���d6f�|�>��r�e� ���B�}��4&��ڃ�4X[o1�w��g�.�A-�0Lh���<�*��4,"�y���'Ii1���-��蚶1�����F���]���I�W�]|E�0�{�dM��ᶡ6�������������~�$d0�����D8W"%b��[�R���3��|�ؽ�IM�6� Ɂ����aۼH�Ze�ؾ#.N�����f�@���r��s�
�hd(����Io�j<���zH֛�z@�ɩ����_�uE*�'�V�ap����h��;�~c�(���!�M)Oi�)gt�]Lxg��	���#��g�0��B��v@*f���0�,  �K���J{9J��p;��ì	�_�y#�@*���~�i]s4���Eh�����z���{��'��ݗ�����J �s�+�����$\sR���*���p������Y�0���d�,>��i����~�ڼ�'��=��0R��1�,��I`'�#f�`��CUj�S^���D�;M$4}���y�<��0�48����L���M�qb�����BJAQ[���a�4T�h@���e����Y嗄�J{��+�i9�%�ǢϺ_R>c�A�$ @�P0A�#�����s���vr6l�HPFP�i�2̸`�@�I:F�-J]-8�^�h�?a1�n�)�fX)
��5�y��UD�t��@< t��e�悙�/��n��i���@����������i��ԡl �?��BZ�mB���v�~xMDے�3|Є��;S���`���	�z>Ø��KK�ٲr�'Y�k�[`!t�ųK�P<��zK��:m㞛�0@���EMN?$����}�A(�V�����F��C�I"���BC{��$R��KQ�$�?��?�N|����xC=���ql���F�]f�tK������ֿE�9ת�Ϝ��T�i[Ռ�����|��٨gU��+��@ZV���Ģ֧�LN�fY��'�sSvmZ�q���Zҍ��!mx�w�!0���3�DGr�(d��(q[��,�ַ�Cd �2%�p�A���\5H���ZY1�l���Xڌ*t�*��;<��SH�j<�+o}���Mk�ە�1�N���xe�G%t�kk"�ՀSr��y�B�kίt�_$��oZ�T���2eG3X)~������84FL�k��o�-��wI5�d2��jB�g� j)����/"�kS�8	�UА�kbZ�K6D�ǏZu�H�\�hc�ɶ�8�p�}��G|)d�t*Ȝ�=q�'�yy�0��t��
�p��*�)A,�E!)�[�w@Bay^����$��we8V����B�\-� r��,!��>cH8M��o�)�*�4���8UJ���"����>���������`*��p��{�n�h]Fg��0T�3d�f[r�*"��.�r_���iF<�̼3����ƆN�p�������N9ݸ��ք�nI�2h����&~7�~�e)Q'�����{�Z�a.J}WʉB9���N�-��v��of��.�\���U6L�=�Y@�7�	杀�s�Uw6-ƽ%�4���@t���� �t���v`����A����h;X� '�,�B�E_���+iC�� Q֖-[�q"���f�w�}7�ꭈ���]zŒ�+
�3�Z0��c�m���)�!�2)jUs�>zu�˴j�f������B��*�'�d��� ���B�n"ɚE�=��ә�/]��c�/��b^#m��<4@Xw����X�,���*E���v¥tՁρ��'��`��e���[�lP�����h�޸� ��6@���qV�KX	j�����p"I����]��oo�9K�n���҇�p�g�r��C sbvG������h� k l�"�J��o����"���z�N1(��g?�g��فo�n钥�Ϙ1���-�Od�@��}�m�N��a�9�DGqgQ{��g8�/q�ೞ�Lt�=��eˠ����y9�H���̝;�Se"���{.� @C���+3���Id�Jh¢/sSv}����8��4��+���� �C�âYn�?��]���X"�$*"�� ��c��At�_;���* �&v*GG��L�P�&Gl�Xad���^����_� ��!C����f���������d`��X�^�#�Iރr {B���7�#m	�Z~�u���(�Ţ�@ =fi"���K����ԔT:� l��_�}���~�#,G@@���`1��*2��5��P _��H U�.p��1DO��'>A31�3v���B\_"���9܏�2��rHY��p9@��\記YAzB[@�]��tNY]��㡝���@��"3$ee�r�p%�D#�L�P�=��,G �����Ѹo���� ��� Z�'�p���>e���.��#���o��wQ?�I��aQ�,�A�(��K������Da�N!k.���������*΄k����Q%�����'��\O�>���4��;DlLD�C�d�PD�����
d���0�E�
Tc* �y#F=LM�^R��K�!t����ߩU^8�_���ԡ����ld;8��\>���%�\�!CX*�����}��%K���mRd�9��) 3�E|�S����v�1��M�N;���c��Vr�UU�q��X,�5���;bW�Ry�GÇ��XĦ��ZY�p��/D�\�n���|�v�,�3X���e¨�,�3�=H�'�fx�,���5D6�mao��F��xa�1�	x�&˜���%U%�@�8� g J����T ��~ɒ%�DnP�)h8�ԝC����TO�>��< � b +��#@�
"
�a!0���`�0��V}z �Tp>K�K�'��e|�녕��(���'��@���_�2;D���_���R�B�B�<����z4ˠn`�f��lS)��^ �x����\���� ə��y��S��0��<��nm#��`�g��r�,[�凫Yjǖ#`GHP.�.fݲ�	��N����-ā+�D��, ?p�a93��s�B$S�/�؆t� o\C4gd��k�Zok��40av�%�y�V�!�l�Lp���P�9��	���'�S�0D��Y��\���7�'(+�D��C&\N߶���YйY�i�$�Ơ��^��e�{Ǉ��$�Ph��b t��:t]]��t�eG�[��ާ�XE_q]$ٲ�g����6�+���>�H����O���d2"ݫ\&,˖/��"����&��>ș���(	Y����I��y�x%۱	pd�W��C�Ůz����f��ZZZ�U\�hغd�H��I����Y�P�*B[;��0�3AR�Ĩ� !��tS�o�ы!�x���YY'M Y�3*SOa��T����5ϰ�\�g%�@Xr�~�_�A���$��`��uG�����>g���*�L0d?�]7�0���`��o��rx��͡T:N;��T"�æt�#�Y���#��K��]�i�0�> [w��e|q�-9" ��p,�?(��^@%O��6���r��cP�h��%p
3v����I�Eڧ�ƀ	?���rn�AxX��R��јͫ|ȵ����8!vLX"$� F,�	�a��sNd97�w[�P¸zܱhi�����0�$�A���=���mu��5�\���!RF�@tJL+1E��/t8	���<W��\=��l2<8�l������C��R"�A5�1���7�ܴq+�{]��j +�D��^��v�A�|-&%S��{i�^�s?{�u�ԒR"%G��GV��Yl*� ��ñ��U.��LGw��;y���`�K"/q��;!�%�j� �=|���`-��6ᆭ�~��`�X1��fN��]�og\=c:� �taǨ n�Gc]L��ٌX:*�?��;CdU6C�u�P���U�r�0�10"#���zv�bօxqL)!Q@'�|"��s�� �@���A�lbׅ$Y�C��9���h��u��h�ȱԶ����p��jK�l+F�T�b1�J��uS]}Ŧ��9��Z�#5�x�J02���1���3�z/��+�T�!2c��U�F��p��X�N��	~H�S�9�1r� �����B$�,۶��dɒs*΄�un�d,�H&�,G�1T��e���,�+��l]W��eDp��	�ʻ[��u�2V,���2��v�J�V��<���s���:��О�1 #h^��Ndv%��ۯ,��)�) a���L0�%R�t����9��葿���珔L�����*��cQuM�z{6Pu�G��z���C(ѓ�_��z��)�Ĕ��L��uc2Dď�U�����aܕ�`�~�w�ل��	�$4ъe���
ڣ8NESFy:�	��H0a˲lii9�� �sЄe�\Ĭ�c�;N���=�~C��
��8.���d�:�fK0����G/`L�WʔN���!j�,��rv�֡i���Rs��<{�ˬ �UO���"4�B����5�j�אَA��ɁT���>���2S»�1�.��:���9��mS7]��[����J�]1�u��^&��&Ǎ�at�QG͢�.?���g<|���t٥Ki����%��5̂�b� <��S]����aѢ@�\E��6+��ܩ/�2(69^pI�7i���l�I�H��1:f	��94 �V�q�����2�z��{���%2�	x
��ߗ��) ,[���6)�(z��ש������ib�U�4ȕ�`�|���.��v:7Tv�Q���\�$SNc����k�ԇW����g¶��pH=Df͘�}�������"v����?�-]s�w�Pu�Jۈ��{��ldQr���I�g>�x�}�Ewu�袋��G}���*r=�c��k,J$�X��\YP��d�:���-s?F�%�q�m�䵰L�0a/�����#����I����t�@'f:��g�l9R��e�축M���qKȂeY�x�p!���B�uM&�u �6�_#��} ��ʕ�Qo'Bf����=�Q,�_i�r&#)����B��v�w�E����g����R���5�G�̚ <�H���{�5��X�%:`�T�x�G_��{tǏ~C�UM����2c̮���6-���L�5)�s�1�ŋ΢Q��y]��6:����Օ�ɠ:R^�#"��lJ�:��[p(��_1������:�LT�U�~�1��YO��@X>}�\,�N��H��8儹��>;�{ ���/^|vESY"w��0{��ݖ� ��;�@��]�{[0�� ��gJ������Jf�1И�V��#��Y@c���Y�0!�	�����~���e����2�DF��ش�t�Q�i���я?���wQ�WQڱ�@�Z9@��z=�϶�]<����(}���c��x<A���~�ӟ�A�=Y��p�CZt�-�y����g* (���
fFy (H�3�~ f����'�}�, ,�$�o1=#Ć��f�2��R��yB:���+V�8g���{��{ʐ�|#�e��[%�/�T�NF��Jv��F*��a
MES�Ҏ��Q �W����Lt$A��N^�������X�Ɯ��}�Di7����lJ���o��1C�l#�d$)Z�rV��fq��$UW5Q�!rU�s:}��̣����j��t���"��ck�{��0�V�����+G9�g�Ad������* ,�vp��������a�f��'�E$	;��q:���H�l��� �ͪ�m2��
�n����Tt�� ��	O&�°��̒�d�w	�ֽ���v�L�C�꥕+_���8Y`% 1�,8�����<��������_C���҅��4t�8:�������(ք���jiJ�{��;� �I���y����$�4�B�
��;m��! ���]�E� ��C��R2��H,ʻ��%ۈP:��6�Mv����7KLK|b��>�zM�x������;Fk�;�d���S�r������W^ynEA��7j_wkM�{��ә���+�k��#t�~� ���5�	��p�Au���/Ȏ�i<� c�x*�dv�:�7TQ�LJ_-���1�c�Ow��|�^x��`��SQ<��a�r�}@�1�2Ps�4��v��C��I���"� ��ҞK�!�b�h���`��b�����qd9�0�8���L����e�BLX|Stv[�g�.e�\	]�5
�lXo,�dS'�Ax��˖-;w��魃id7�l��zk��5)WtxBu�蚯1��M��5���ܱ�L�|�U��a�r�,���o��+�tI�h�.�a������������
u��N������c1*Ή{�巍~P�m�
��Kv/��f6��������X�gY1�OCԂ5)����Nd������M������0_t �2扦��]a����ئ�{���yf:�f��0a=�ד��L�	���g�BW�w |߲e��ms��Bn�	���N��BŰrl@��)4-�A�s�lp�Ż���� ����~4d���ӊ`�r^�����TXm�r��^87{:�w����6�p�	 �~���ֶ���@��ة�8]�gb`��5�6��$"˦X,B���c>��
̖#5�\_�,$G�kC a>L��$yn��qҰ���Vˢ���F�r�9+d��%s<��[����z��dG� ��,Y�+�rQ`�����I�2��\�U�aܷ|���*�[Zo�IuMB��D<E�U���dG���rF2L9��	�e��$UF�4�lBJ8$F�)�>�隱x�рa(�=�~���2U	kʌȈ���#�wf?�	���ʡd*NQ+ʫ9~ҴȴmjVG�M1\^��0_������`��{$���З,�o[#nu�Y�A��+�-^�'Y��%xj8�1(+���[�`Ov�0�o}�^la�Ul��>#	�		��|�6�%׍S�mQ$bR:��^�8���f�u��B�j^y��yWt7�I���ό��"�r= K��VObf�|��ÑL��,�@�� �x��">�qQV^�~������G��xG��>;g���)��m��.^����3g�L��/G|���M[Zo�%:&!cF��H-�`}M��{:9���C*K ��X�1x8�I<DT@e��ȳ�>�ɑ%яhf"����908�(�
�8O O@X���Y�Z7����]���R*N6�$�IɄK��"v��$�	"�!;
	1j&)ׯ���GG��<����;63ʹɧ���{aq�	 �^�&,;x� ��b�Z�[3�
�w7�zup�{�I�`��L�ӎ�d�d" $n��V��Ӧ��CS�΢�j��E�[�|v�T�([v�f���|���g�������I��?��o�C������f���M�G��yG ��4Y���Y:� l��T��)9,p���x�eݳd	�\Yn���͵i?w����1��������Q�|C:9��|"x�Rا	,�Ǳ�',T�	�׳a	`JN
+��4}��.��z0v6 ��� ����Z[_&�H��ɱH�5���SQr�AV���a6��4��5���;��wH�[by�Aٻ��e��LA��_�`c�`߷PފK	��[a�,�>�Uib� ���-XĤ
$�6* ̣M��/X��*�T
kO)j�4���jklNs���U�`󇣨y�Nd�H(�o��,Iؑeq��
 ��aGu� F=l3����^z)��u�]�dO�S�Dx������ ��^�L��^a
d�Cy�+�c/L�+;6k$ϳm��ŋ_0k֬u�i�E8�޺��LO�TrrG $�����9���7��-F	<��p]�Qd��4 I�![@w������h?�F\5�s` �k��H�P�����w�R0:���^��Y�G)J���ݽ�b1?�r�dU��[hŊ��֭.ّ*�.Ǔqf�G~�=a
��.��ϻ�`���X�B��̪ �U��g�@F(��} �K�g�jx	(@X��更����a�ʻXD�ʤ�S`�!>���Ѻ��ɶS4���>�S�}G�1� �xJQ]�pRf-��DK�UWײ��Na[���i�O~�LĂ�q�㫯��������9s氜�裏���!���?�C��ȓ�2������%��ʲ;������������>C���D~�hѢ���-grOo3a�0nn��It���M��x�Lx2���3B �� %F�5��7��'d��p�@�R��5���������>%Oh ��K"��@��������˒D�;�V��$iܞ�����s3E#u����􉏟O7C��%G�)4g�?�|�(���������Je�ʻ�T�	�re#�j�GH�~N8D++�`�>ɏK���m�4��0�a` @�[��6/ۊ���Nx������G"�륆Z�/�O��9��V�����^j�HS<aP4�@N��>S��z1��� ���G�!|o���1c��y���/2�A������П����7�̒����@`
��P�ꃄ�M�I$P�_�XX|Z�C� ���{�e�����"���-Z��� N��z/>L8��s �O��#�|�?|c�#��9�0ȊC p�]5*��[��Q놁q�:�(:묳x1��s��N6�mI�%+\p.v�����7�N�����:=����F�l�̙{�n���xo�^}i}�c��4���(�d�s��t���e�roO�L�����!�����E.����Y�pL�9����|W�����;����;��Z3��E�E���g>��O���sB�P�+_�_���DnE�]�x>�|ұd��J�ko��g�}�&�=�jFS*aR4VO�
R��sv�0������a	�����?�����3����d�©��������'^ G`ta`
�駟�~l
&,a�����*�u���E��p�������.���-J) �p�*
��˖�	E<"v-��1��<���]�7��Q�b�|������x���l�=�k.�M��\0�O<��xE/��B�
]u�Ulp_���������׼�y�vut��W�ڶ�@sN=�.��T��W^�Dg�u)�kMYu���r��� M����^-�(�����s�����Lh���\c _�/k �K��cy�r�+.3���}5�c8���� {����L��,l 8�;���;n%�레�K�z!���㑏����7�u��]���i��#(��)��D5{^�}*�YL��3 m���C��R�8�́�b��~.�
�|��\�8F�_    IDAT,��<��.B�d����?:�.A�����cG�O�m۾kѢE_�(O9w����kni��T��g1���/Pm]�|������Bb�͊sM �����(�P�d���=v^�f}�H�y晬A��/}�G(� c��C�\�&�r$װ��E�o:�����詧�JӦ��o|s�3~z�����ͣT���	?�
�W`���79����Qc������k�>��+K9V��a@v�eÅk��8�xa}1�3�%E��tr�i9@8��JU�-^|}��'RWw;-�j=���4z��w��4}�!�(Faf重b"�%�����u���>��>�Cd�������±���+H��ԧ�3H�
 �z����(�ɕ�<�(.�!�\lf��������g�毮����}ϙ?s��ͷEz�L�i~�F���g�m�z��'�̎�_q�nZ�P���#`D��3k�,�X 3�%�~�1��7�J��r
_���cP���Q�!1J�%�a3?8���*<iX�����+_Fo��53i�U���L�Wm���9�M 8J
��(F���~���AKB�B .��#����9����b��$1��Co)=����	0�Y��~��[(�襆FE�_�Y:�#�Gt��W�SO�Ұa{З._D�L��'�1���Xq���L;���J���z��N:�N:�L��K/�Dw�qmذ�/^̑7�x#/�8�/q��%��AV=��2�H_��@��������~0H��tJVṑ����._1��ɓ�Ʀy�#&ͻx������${�q�]e��	��=�^~�Ez��g	���� ¸A	'��1�'`(h7�
��2�
`��a��g�i����aA�q<>ñ-Z��� �qMLAp���>�������t啋�����A�^��&Mއ�{�u��GϦD2Fi7J�YEdD��9gp��q!���Ǿ�,  �曯����	�vwSuU�/9�N��<K����7��'��iͿ�2�c�=��7ͬ��N��㽝��C�����А�v/^������s��	'��}��?�}���e���׿��H��={�l:��=��;^� 	Y���υ܀������G�����M]��
Ѝؑ_/Z���Lx�s/�6r�[�ե�3"xISt�!G�	'|�{��f�2]dK�%��������L��w=='�PBBB "Hii�@��҂!�8���w����f�$� ���)�؝QQ�+�9m������OǓĐ'�u�u��������_�~����?DfI'Wp.L�����Z���p�҆��68���"|���P��r̄�6\�n����^��]{�n���q�����[�ՕU��R/��1��� L����,C}��%�9�t�}�*�rjk-k��߫/:5�y��g5��V�Ԫ[n�Co=��`�V��4�<M%��7��d�~����[�DE��6��;묳�S�����'�ֹ�q��8�Xm�|7������8�b�s-�n��N}���3�ל�r7o
�S�V+�T��;�ν���L�8���=fӚ�z:�F.: |��O�y�[?��g�a��s��7AB��:�!�r!�)��@]��Þ�|�K_
�{��;<��0e p^N'�fr8�c�%�s1~�bHV��ٮ�������Z��I����ڔϕ�nMY�w�r���%Ӥ �f�$O~G�?�����k[�e+���^j�&}����E���Ƥr��^zq�~�����7M��_?��_���l0fHS���A�!l��	����)G�ڈ#�y�����?�A0G��7q�y���d			"�t YH#�P���+w�h�r79`���4L��JWM�SO�}�]7�r�)�WE��o9j�����Ӽu�1�1�2�������^�Z*�IPI� ��TX;�� k5�5�����Yp�q@�^y��9���<,+戾��t�؎5��Љ1�=!$-�}�7YU�	�Sz�!l	�U���P�{�K��1�C��ɪTM)�	��4y�t5n���!~m��P��FᕫW�Ա�CMMe�}��5mƹJ���Jjn��[Kڴ9�|>�Lj��R�{�q���tD/%���1�Ad�=��}�X�17`�%�!�c��v�i�q���6��"�O�+����X�ҥ�}>8���Y�|ꩧ�y�ۄ��L���wr��Q��lZ����?��,"	^�a���ks�F}���U[#��W�X\p�/�a�e�sh �EP� :��dђt�+B�q�� 1��s���}��� �j�☳(�����\k���y��[3*��)��kX�H�������ھ����&>��*T�԰W	����vH�	0��s���@�ZHh̨V]u��z׻NR6[V:ԆH�\kTwgM�T����*�Jg*a�Ѱyp*�+~��<�i��aj�[�xm9A�7���G bS�N 68;�u�ĉ/���f�,0	��h�+�=�F�tWOwg2٧�y���0~Ӗ�����yՂ���I�#�Lވ��:u�8t����3*vcG��h,����߀'�^<������9��H?�&��q�{�F�5? 3�����/� ��a���X�`SvP��s�)�8kz��O�k���BO��P�2���k�(E�rج$N��K.�l��UO���x���P;C�/��C=��m�n7ftV�U��[�m�*U���ǝ�7��r� ���BoAz�I�,[�kD0�K���#����B�0���ի��;��N���I<'	Q����w`��8��`����ӟ�e���V�@��s�D�Z%c�s�����xío�i���|׉�d-I-��d���Stҩ'襥��r�������z��:i2:	���Fh/����C��6`�>���SO���]�Vs��	6c��m|7(�F��6M&�N���gU��:gRd�P!��>U�V�V�as�ƍW6C�r�@�Ƽ��kH�%+i���Tʥ�%ns�fʪVzTKBrjjl����Xe�#U-g��ܤ���`��ը�V�K�
[454(�ӼP 8�$���2�!V�����,=a�u�5��H����P�j,�v���k+v�&Rۃ�@���.����j�J)˯͙3gp����_^�pT�<�;ߝhmjU�3�7����2���5��g�5k��ES�ދ 錗f� "��I�-i��	=���3_(ڇf��@TT"`��k,���7�d ��q�۵t�":+��m-( )_`Ś��F���QBS���QGMP:�[����~!�PS�Z1�KOH�FU�Ez�N������6��Qo����ViPKK�����j���z�p>` ;��9	V�z��a��s��F[�3�ӎ�]̙�� v��6mڴ�z&��2�{�F6��ɢ�j���}Y�qސ�k�H���ܹs?4�E��ћ6,l��6)�I&��/Sa��u�X������MZ�|e�`�m:�"�N�0��d�j��x�t1�`r�Y�pZ{?h6�f�-溸� �����v����^\[��|O=�;Ö0�P*�6B�Wo��a[���
A���Pt�^����$`^�v�>���T쪅H���4jX�O�Jgq�Q$�Qg��B�:�ڢR� %;��)U*�@��G# ��w0�����vK�-���~�^"�LxhBÆ�]w��#��v];��@���8���xa���MM ��G[Q�"HP @�v���Lx�A���ͫ4to?���A����2h��*��:�Lw�[C��@��8:�Tm^���/t��? ��cE=���P%��% ��DG`~`9�&ta��"��7�!8�=x��xƌ5�(�R&�m���eU,oWKKB�JR�}~�>��g�eK�������Sg��!~���P�Q�+����ROU�nӬ+/�9�P�,�*�H�FU����u�R���������p?Ha_(>0Z�����?���%�)�6u�z�Hڊx^�s/g�b����Ŧ��z�OT��8�_	_m��QZ�M�6q�������	£6�Z�Z�91�N$�@��F1���+ۘљg���?!�V� 1�s99k�g9�ҀNq&�t �������\G�������;��@��a�$k��w0�2ib
z�ڵe�
e(�פ�/n��ݤ��ʵ�  L���(C�A��C���%�	c��֥�6��;ޫ����/D���`utI��P�I�r���l�`Xg�;|*.��5~3���RO|3���0��~z��:m��!8�� ��?f��W↹ ��~��6 �	��b� ��x�z�Q@�����Y�R�>��J�mI�=eU�5�(W�Ѱ�vM�0Qd�'L� G~��� a�t����g{@�(qu&�
"h�9;��N:�t���(�	;N8~}�a�U*t���򸎞p�N<����Vuu�fUQ^p�*�*ײ�
E|�N�g̑m7��=V5pI� �b��������'t睳t�{NUcSJ=���,ڬ<�k�t�jh�Z5�T�1D �{��f�@�d�x�3�Y5ϛ7/�%����e25�1U0�!|��<G? �|G�	��s8߬����^�S$������O?z��7 VΟ�H�Ά����	�E�a(��÷�'���cJ��@g)��vT#XG8�e1�D@�|�^�z�i�:���	�Q�o�p젣��|�>��U�nҥSߩ�o�'w,]�U�\t��y�8U��as�	1�}4Ǉn��K� �d�KZ��Q���WB��E�X�����O=�mۓ��#Җ��f%�ٰ�'�!2��'���C�U<d�3w�4���js]	���fe������������q�iq���^�Y���+l�؀c�2�5��+�L��a����$%��b���d��锺J��nKSk�xd�@�`��~m����(��L�^��pq�����ý\�Ӷ�s�m���r;8F�U��z���ߵj9�[>�����o~���8L�����qoђ%�4����;�r�A5���h��{A�%�s�9^5oH���r�r-|l�r���f�ϸ��@���������G��YW�_o}�۔���Ɔa�r�y
q�3�	c�c ���A�^ۡ�����&�l�^��`K���ڮ��u|/�
�����*��s eL|o_�K#ĵ���e��|�I�jI�M��娘��R��j�.0�t��i�5���BZ�YPt֬�5�^�g;��m֖|g��� 3���`Ψ	�^-���S�W�Я�S5������'u��oՒ�k4y�U*{A�-ﳚ:�
u�ذ�V�N���e�탩>t��Ua�'L�Rʫ����o��)S���C�S����>����;5~�DQ��'_P6S�=&���B&,)��e0����j�ؗ?���x�k 2��:'�6f��zTŰ��ͦN������Lc&<w�����>$klX�c�$!jDG�Sź�y�j-w6��^P���ef�d�8Y�%����~I�Ҡ]�j5d�}|��ziɯuđc�����z�����+4c�u���ܮD�[��2�2����U�wr(cn_�ܡ{�	$����+ֿ�+���pJK����Y���i��>��Y�>������}�k?Ѩ�o�-~��;A������j� L6m}g�N�c����v�κ��{�|?��jb��cL�ܸM�f���͛w��g�mX�������
q��Aة�����}9�x��������{�Ś�O��������#ںu�f�:O7�0]�����3oԶ��pk�'LL�)�4~JgJa�!ޗow���^{��Y�A}D=]���V�w�O�M?O�B�~������K�])}�c���'ջ�H�B9��-��Y�9
�p�R�o� ��c9D�^��b��A�D�7�HV�fD������AQ;�ڏ�i�5ZK='����� �j�7��� �|�����UԦ�ل���ZY��=���}DUg�}�F�N���G+��t�����=�a�Tk)M�	O�4U����ne��yod0t���0^�|��?����jn���s�Ռ+�W�ԣj%�_ܨ_�b�Ǝ;A#F�JYJ�YU�4S`��r=.��)vְ����4����d���w�}�*w�-o��养ao�=� K�}l+��聾�0Q�'_X���_�����8�Q�G��jQ��ujj��UW\�amݒ	?�Z˾]���
5��-1�;T��OC��Ax��5Z������̪���1W.v��+��ھ���N��ܤ(�re�)�lP�R
;k�����p���S��?N�ʌ�k����o@�}��ڊ�	'2G$E��]Oe�A��(	��q����c���	B����T�յQ���RIjWt���]/<�^s�}Z�0�j�b b@�>�O��q��Z��S!�|H{(�Ϣ����Z�i��.��.�{�ijlH�ɫU2l���SU���^�;���K�P}#�L�Qq��6�U�>X <w���M&�;��S؄w&q@�^�r\_m�?8�b�����*�B�����+�iR:9J��Sc�p�j�&߽�iS��رG���C�O�@=m9�UkW�GV��!ky0�Imm%TV��h�v54���o?M�����&�"��ެ�z</!a����Ef�3G`t�6�[����&��:l_
�6�P��������c����'�DU�D2�B��5�kUw�08�F�*I��Y��H�bHN���X/6=d�ؗox���V�����];b��Ez��G�(ה�+9�J��	Gf\*Ѣ���&s�Z�[U��C"V!_	)�6E���PwQ�cn_DZ�c��L&��3g�����}Q{y���RQ�QwL����C<���ŀ��.��xa�I9lj��m�`�d�lZ_�(4Q��0��,���5hh�	Ke%�)M�6Kcǎ|� \���9b_�١{�{	�/[]�rc��Z���
ʦ��64��O�y�pr�a�XcsV�JU�JZ�dF���1~86�ٲ�������5@��s�̹aPA�^Em��ƞ�I�L2�L��</�&5TC� �ɐ�P��o�+�;x�I!s�d��x@~;��Kg�8l�b����f�~�xPU��������[�D8K��̏�C[7n���w����jZ�jc�u�$`U��-;c�<����b�	�\{���^�������*��C�Ր��!#JE�4�T-ըc�9Aox�[�/���w���Q�=��!i�#�N��3ژ�$V�)��u���%��9B��;l�����z�	�wY��Xs�1���Y�={��&MZ�'�m��	7���Q��>z@�vR�Г`��T�j�j��/�Ԙm
v(�BH��3��������s���:Β3�v�˲c����]?���7[-M�ri_���/&�eIԣ��uИѪ�s!d-�j�ꕝ��;U.7���3�1���)��פq�C�{2��ݟ$�w ���Z��Q%*y�SE���t�{�PKK*�(���`޺5����a'�R1���ȐmZS1wg�1��/~1��Lc�5���ט��Ǽ�{�����=�'��=�s^9������9(F��l^op  ��ٳg�8� <fÆ��ʹI�b.TQ��O�TT��U0ឞ|p�F��|�^.!I�����`r�9��zI��d��C���Y�X��ls���F]uլ���	����Z�ڇ�4rTZ��F�#_]Z����}D[�$U�5�k��ڛ�\��1�����O%�`fL��l�j�_����˦{t���5u��*;B��D�U�JV��m�-*����ԔN�����ZNJ��u�� ���BJR�<x�8��} n���w�뚓K�� �WٜK�`�Sٍ�c �[:ǳ�cP�R��R��x��M�8��=y�d��|����S�7M�6�m8Ԏ�]Y���*�dGӱ��%U��=q���t�P*�S�3f��k    IDAT�6iX�,y���Ջ\���Z���g͚����3`�����n��'���I��q�^wp��wvj�҂.��fuw��Zk
*�	��P:��VJ[ޓ7t��	�q�=�ϪV:�ؘ׽snԥ��T2Q��=�\������c4|䡡VwSӨ����H��|�+�O�	�1��l�%m����:+lr>XCUF���!���� (�&x.�p�����JYj��fJ��ZĤ_���a�fV�v�̘�+�J%�L>����4� <f���M��IM쬑/&�А���V5�4��'��N� �@~��0A�ri��v �E�@�)=���?��E,%8�=,���6wxGf3c�-���؛8b�QJ)ו�,{��t��g��NVk�0-[ܩ�fݦM��� \�ԩ�â�y�:d���+C��	�W�Y���>��6���{�����V�����>���UwwR���7:�ȉ�犪���S2I�r J`U��Ļ�Pj���
PdU�R��}�[21������� �ls��U`|�ƦL�(\�l����2����N�j�
?y����t��n�Y�	{�mG�oZ3���cgQʒ퍊ł�M�)��]��rZ�	S�޻�� W;�EP|:�DA�z�O>�d d�f��jh��m2�T��v���W^yE=@<�x��� kI�[���KK���Ԣ���7:���Ӣ�o��iׅz�;@xGQ�T�h�8�����K:wH���K�X�D�y���m5"������s�Yڶe���S����ZZ�wާ716�0cd��u�H�����  l����/�2�l�.��5��~0�x ��am�q~���N��g� �"�`��^���f�@�� ��`���7���~����^�ʃ>��Ae��m��7�t�H(IC�I��]��&�]�>G�-[��q�lH��C`T8�cMf�(l�6�c��^����4/�v�P��P��[��V�F���"Dvr�:ur�vI�`}fI�ۺ4w��Z��Eez������3V[�t��SU(4�"�	�{�	_��L8קþώo���=q���?J`o
��¼]0�a�6iԨ�n��Z]p��ܾ]w�u���!�����Ə���C��r����|T�/�~������3���g�s�'?�I��:ʁ�������^q-r�6N9��ٟ�Y���e˖ ���`��s��ζiv�`�
̨�<�LX�C�= �H$���'>q�����7to ��ܦbG^�v�ο��=f�^��"�Z����P2�A(�Lh�p1`�!��ݖ���ǵл���`� ��t����p����aՠe{CM6�+��<��CT�@ǖ-���}J���Ot��-z��������/,ѕ�nPG7 gBhM��p/��,�K����N�?E���m��u����Z�r�.�B ᖖ�f���f̸@=]ݺ�������:\7}�M:�4u�t+�a�	".=����6�\����
@���؟P@�`[2�U�\o�����??`&-�9:�@�U�#��3��6p�o~���S/�+'��'|��[���8?�u㉙lJM�-*l���<C���4����Z�z�:;��	@"0���y{Z�����#
+��1� .����f�N�%aI��,0i>f�ZL3g���,�ӯZP��Mw�}�zz6h����ʫ.R���z�՚:�usD�pR�DF��my�8%SDGTT��ل�h���x�D䭵c�ks;gm�w*�\d;6�Hj�kCk+W���gU
ݡ��=��W��|���o���-�'���l��#�Go�t���J�e��2��0vWp��N~��O"Q�!e�(+p
��7�b���WVӧ�v�N>��p� dmN�M�.���:̥�.~�r��`�t0�(���N��<o޼[�&<b������]ԝ�.�l�|���/~���\�� ��h��.�(<���Tl@����~W��կ�0m.0pp/<�쪊M����Z�e�8�aq��;k8��w^�d���o_�!�������MU�	�\֡)�?���&U�TQK�p�@��{��a�)6�;J��1�����"�����|ò��=��(�L�1�Z�?I� �l�r=���Ky��U���/{�e)QYL�w/lҢ7�u��S۰����Cj��ke%��Q'P�	������}V˄��{K��r=�~�<s�k��N�0hB�p�a�4�3�5p��
��/|�g�������o;���
sD*���}��w렂0!jlX�`��'�+EU�5�~̡�����m���_�,DX�,&L��g�5�uv	�H�8r��^�9���P}��![&	���/gZ��bc|l�Ahl���}��f�;c����9"��L����ש��M+�nׅB�E55�L�P;3J*�[O�7����ncfj�J;�vV����WVT|�跗S�����u�ܟ&�P[^��KC5�	ko��=KS���&Xn�r�mڶ������{�3�bK�L��(/W��W׀����0����-�?�;wn����W�vj'� e~c&��=���e�L�6-��f��0�AI���9��7�������L��G[X�s'�Kj�Z9�J}y�A�����ױ��-�Z��;Q3g^��|�b�k�7�~����+* ᥮�6tA�����da�x>R;� ��.�(�{�����6D� 8K^ ,!��$��}�{Ò;���	R�J�Q6-�z��mXV�|I+�n��om��S/e��׉�6u�ƍ=��9� ؄�|�q��+L7���)F�x����7d��p:�$���;���>]��i?���I�$$kZ�j�>:_���F���_���91���
#�+�ʹG�\���L�;bya���as&,��/�g��v�K.�$��(�M��ډ'���ް�x�A� T�;�j�S܇U;�8�29�����=�d�9�;_��v}f���D� |��'��ߣ��ڼu�J�r�	�����j�%9N?��p��A�'M�:Jx�w8����s��9�ӷC3���p�eP��=�RHX>x�/���� ����3�UWG��Ŝ��)<]P*1LK��UCK[HJ񌡨�� �
	��W˄��m6�2���"!N��>�]6Vf�S���
����r�I�^d����	>Ԗ�_�k���{X�BV�ZE�N����o�ӓ+��Cޠ�O����R��U�Pϐ��V�Ř����g�������k � I�*��m�g>��w��L�iچ)@uL���� m̞�1��8D$q˽��1��=��s۠�-�^��ݖ)����E]�����Z�zE0G ¼�����$��!cǍ3T��a�,3(t����2�����-\^�C����͂����aN�EQ/��H���PH$��A�Q�@TG�
�j��ɢ*�h�:Τ��I4�^��L�]~����'���z�:Q%����8+XA`
r.���1+����P�'	�A��%+^�#_���ڕĴPٮD�:UjUe����:b�jic�܆����)��T��ѕӜ��(+��0q�_}��!B��9��SO� �c�k��� p�;S�8c"�i�c��ۨ��<�Wp����q��3��
�ͪ�w��={�-�
�0�Q�V-l�&aFx?J�_>C�-��~���X��P@x�ĉ !a�Ȅ4�S��8?��9����`� ���Z�[Y#P/�]t�!qQq�Hl�@�uf\Q�RԢſז���I���H
xHM�����J� \Ӕ�3��Ã �������~����]B�V>V4f��ӡ�(7!���q��4����ڐ�Axպ���IU�傚�j��u'X�Y�L�&L���*���9�&\VR�>s ����ς��9⪫�
�"A�0����>�g�� <s\�0O=���Kd[3`��ò��y�
@�{::\���b�zI�O�}�݃�#7�\0J���{:��ԪCF����J��.���.؄q��@v��4��q{����YN����l%�&�%�� Ll<�=�%��
�հ���̆�X�����|n�~����ٱ-���
��4;,zi�jlł�!U7GL���^N+E��^�1'-O��񋱩Þ\;�,[�}���^ �d���V�3^S����l�X�f�}d��]R[S�ڇ�Ԑ�&��Ҫ�����>H�}�:�����@��WQ��	��:v��7懛o�9���8��l�Lw����50���
��|�+�r�����(!�S��p9n;4�`�&�����L�"�&�V�~�{�yP�	S�}����O���H�5F��ݺ��[B����%55�v��O%��a�6Nl,��=��H������;��܀V�		AЀ5�<0;��0d�H�6Q~c�L���jG�T
�Aw�>���*�rJe�J%�ܯW�{�B��I�T�M��d�: �y�;�#����8j3[�G3#?�o���f�^p�|lj�o��6d�(0;��"��0#��]���-�J���%����0bs�����Ǳ؁h��a�~|��!�����'c�o�e�p��WHV�nw�3���{�zEc�eD[�N$`~���s8�=��8}�m�A8��Ǟ�O�?/�}̠�7���dM+V���?�\G�=x����<]|񟅚�L�
��R�vmڜS��c�=��R�=�ݳì�L�����7����I�/D"Z��<���{�a���+��2� �I���	�x���L���yLÜ�aA8�o,��p:�~��{��Ƞ�1��Ft�_���v2���������N:F���i�˛T��sw�iϧ�;�&�'8��d b�AS�>Oh���_l�a �����*)q4��>8�x�Ax�ῨJu�F�H�o8D6����Y%z�5e�5�盂3���$l�퍨'����%�`�������	I�\�;u9xI'��~����'��<ϓ؃� ��������!;?׬����:l��\e�fE�wo�j��~��ab��z��������4էhl#7�������0�8��Jn�{B�
.vj���2�ǲ1X��v�ڔ��ξ��&������^���g��n��ݯ�]�A8����ݥ�l�M7O�ԩTQc�5dҊU�U(��N��(-u�&����=F�.�>�\sM`�8�*�[�2�����o�'Vӄ��^����&�6K �=��9��Y�C���>�{s�p*��ڽ��{Ӡ��ȭ�6�t���ܐ��O��:����i�Q�!��~�֯����^BG~tfANU�0�J�޿���&����� �����n#�'��3��L?!z ��z����|�T��%U��o���ƌi�{.<C�-���V,�Ԍ�7��3�J�Y� �鐬1n�X�ӕ`SN�2�k�>sG/H8���qW}�9^5�@h6䕀��`&�I�Ak��{�fñ��@36+<4?�7@���i{2h�1ӴYē�>���ǌ���d�x�?Ã����m��=��$���f� �^_���&O|'�� �qj��L�tr?ڱ���឴��oF��gE�1l`������"�?׫�6� �Y2�e+Vh��_P>ץ���u��v��J%kھ�����J=��M8���%�J7dU,u�S�EdU}{4�.ή�����#��E88
���г����c.��� �ؓ�+�>���w��x����&L;�+˲w�� �9s�|h�A�mÊ����I�R>�Ne'�	�x��B�U+VkѢ�B�bVeA����d<� )��x;��^f�)��{�qR�@h3#�|�|�p���\G��N�Ɋ��-�}�Mںm�.��}�P*����AS'_�Rq��զ�-'�5u��^.�F��pn%l�֎R@�xbz¡L�rI��X�<�e�cv��;E܊�l��f�?�gGGxBs-��خ��������0:�ȸ�eO ���cFƳc`5�5Hr//�<.��v���\�UV�0��0�Y&6�+��9�g3٘�ǀ��C�����y�N(B&1��qR�MQVj;Sd|O]��c��(�X	����7�Y+���.ї��E康����;��5����ݟ�>����6���;u�o�鰠.W�\K)Q��Q��`�a�q�	s����� D�^�+p��j�z�������I#��3���๏A�d�c��ް���|�+�1�|Md��j �{�w�AxĖ�G�J'���)jGx����z���j��	ڴiK��X�[��n�@a��	@�{l+[3{�mz�'OA��9္1Q<�< "�)N=��}���i��c�|�����sp���?������߭�{�3K��U����9������ՠ�U��kRO@�(^@�l�p�h�P�|>������sO��0P<)~����;6�&���`�b��1�`�2-	�=/���6��|h�%��Y%�4�q�������+f�1��;���.blvn6�d�-�U�Q۞m���� ����l�1�s�e+�X�Ǭ�J�כ��m{��?~���to�0�{i�b=����J�iB�c�.��L�x�+}����<\��>W�&�j-�r%/��Jg�D��)��i;~�O}�S�= {�>x@������n<_p�"#c��Am��q�U�My�����}�k}�����d20��	صaarۦ��!j՞��U����9g�+쬁p0�tҚ� ��a9F� F���G��أ� ��3L�a ��uυ��	�e��}ܽS&�H�Еל{n����<8�?q�N9��\�E�ϸ^]]��R�0�z����`U��8ᘭ�^�!����><�]��s��ؽ�I΋Ɔk扣�`�g![��#�0}˃ev��1��ywț��0 t*Ê�u=|-�=<�hǸ'�N��`r�ެrP4g<�Q{�N�dblfMi��oȄ���p<�|�mA���@l;d��o��(װra;|	y1��o@�,�y�6u��ܗ��/m�r���ݦ]�*l��6���KȌ�D_9��pQr���h�s���^5�AZ�)�	/]�D_y��ڼq�:�A��1K_r��nަ믿M�^ت<R��:��	jjlS��W-ݣb1��T�T�;�c�W���r3�3�hcҀ���`EO�\ܝ��=8�Y!#gV|�Ƶ�
�W�}������J�8��MSƠ}�8��6MjimJ��A=�l6�|�G�R^��mz�����x>�T��0����[�D��v
�U0�04��ٌ�k�[x+^��`�;�J����V-Z�s��-#���V�;�`-]�AS�_��δ*U��l�Y�t%d�%zkg�� ��b��&K&�MۘD '��53a\����X�Vf"�6@@��&#�8�}l�o�c�e@��� �k1<���J�����asO�E��,y�|��2�20�7?���L��9^�܋PĘ���'�0�xc��!��u��3q�iE;��ל�In`c�"s+2���Y�Z�f�~�����O����˸�Lm�9!� x  &;r����f���`O�#<�c��2`�{�����{�a��J�+���/�1mݼY�����g���g���C�7��S��TÆ�;�Oo{L�W�T�+�P�,YI�o�p��#���{�+f�?Bvf�V&��.�@lvd��EE5�-�I(`wG��G3o�s3�W��
3����aЙ0�a����*I�9loT��U͔�ΦT.��\*�
��&f��P��섁��!����N,x��`�R�����6U�.>3���F3�@��9o1ס��Y��˺⪋5��B��U��1�P��ZkP��P�rf�m9�
gP�>�cS/����D����xU1���ٖeM��FN0 �6@��D�0�,E �AD�p�m�n��&�FG���w�sv�= 	���� ���$���0(�e��;�0��m����?rR    IDAT� �.5�$@6�H�#�8����D��y�| 2���(@�〓MA�=��g,�8�������_d�,Q���x��w�Mڏ�b����}u�
�!}8��2Gބf��b��ܠD+�FI ��I3n�r��(e���嘕;�2xG�p1���|}��|ɲ���Ǿ������G?6C�/;7���������Rg������c���X�E�=�JT����:���y睁�!8"���0����u�Y�>�!3�nPzȜ1땵��e�x���/��(���J���;w��wܚ=��.�7"Dm�5ZK=')QM��= L	�r�j*��s��t���C�����W���IOL�����}�{�+
�Qs}MlɽA�>���x���0�W����t�k�J�lo���.�x�&L�d��&�t2!�=~�{�K��#a�01� L@��pfr1i�����a�ʀ�=��P���z@���I���	���c�� l6��� Y �s̑h���1 �`E�\�5v(a@�~�=?����o�&�p��$�� 5�gs��0`À KD����r$%� ��XI�=�N����
��K{9ӌ��� "
�����;mQ�\K���w��><��slR���{������	#o���j�%��! >���ڦ������ %B�b��W�����0��	�^�F=�9U��P��;��%�OWc6
�,}iS����o9N��c�N��L֓z�+��z�I �E��<�9�E���>��I�.�߻����~;�/$��܏�?��>�����tz���8�L������}�'+QM�)��� ��Hk3/�c��߱���	 <ӶI����&<Px�[��%)٥C�t������s�\�~��m*�S�8Κt�%S�Ru��;�^F�O�τ��g�2alo�\��Ť�@���yLT&�w ,��e��4|�? �hh� �0T 9�,�̓���n���И��;u}W��r��Afk<&L;�:�-}x +,f<@啓��PZV�6#01Q��s�o�t9x@(7�%���\�yȁ������� ������hh��=q3}����N����ʂsQ��$����F�|�c���W�[���{�3s���y���<�N��������Z�2��� "]�s�ua5�ɒ�ߣ��1��Z�f��ŴZ�G���$��)�TO�g�#Ko��1�)+��aj����x�m������[1 ��}����������9��`mM����- ��=��5�����@U�*=��ڤ�LM-�xZ7��Ѻ�=��޿UWGU�23�P�d��u���J&�}��uڶ�6j�E��<�}g�0������1�cخ�� Y���f�_& ��x���ȅ{���]Lfl���
R��"��59�`E�����1{uH�'6���)}`"��@�z��cF�@?m�� �d�� ��}z�8����N
Ϡ��"`�N� ��?�����x��ov~�^0_�L O�0p���C� 6ރK�"G���PJ���D����w���|'�ŃLQ�(&@�U�G���x������A��B��Y�)�}r�(VS<F�����A��3�/_@�1�R��w�:�4���Q����˵�2�[�U��������>���t�Wʴ�Ǥ�v���-�ܰ"�jثgcW��A>^M�'�ƠD"��x���{��?�=}x�������7�o|yA[���;c��t=: ���K�8|� eM��������G{���L���e��FtC�ح���GZ�jE �r�#T�K&��Ғujn�\��i*ժ�L�,LB�t���m�"G��
/ �2��ق�2Y��a��b�9
 `��Ra;aW�B~LP��L@�8�Cl�+���x �XI�T /�`�8�X"�	@�vp-  �rm��.�o�\ c p�]�`6�➀�}(���>� O��p-��<�L
�8�@�D! s�N����(-��= |��ʓ�Se�/rfL�f�N}��<���Q<�����E?�/Ǒ?�@��q�, �ǽ�@�PĘE����ȇ{�V�y()�j��1���x�L8U��W�s=�J����4���?�!�)�F56��ط���y} a�aja��w�.#[V�����$=�-�=���������|��0�o����W �9b@�p̄-�X(ql�;��`�'��.�53��¬���M�Z����,VO��`#.�XK�VmU2ݢd�Q=łҙ������:z^^R�+�/��b"���y�g��� jdò�A�#��a1�3a�,���d�������^v�"����y�,���4��1�Ñ6�7� ��`Ұl��؃]� F&|O;x>��P"+'� Z��A>�>0=;!�5�{1�A��N��L������	
��<��� ��1�hE�;�g�F��=�����M ��G~8�������v:���
�˸�Ǭ���V,���&���7a���٫f©������W��^SK�Q���U5f����c����C_�lC����+W��)rʦ�;~���66��fKc��{��,����8a[q�����nG����>���'��<ۥc.b�;a�	;��>Y�(�X��,�=i�@�Q��9��5[l�B�U����K�
�'S�+�)6m�-J(�|�T���C� �ђ�/M���T���d��H��l��fb���m�LjX8���o�0N�Cc�����M�q�	� ���
L`'4�&�X�k���8 N� R�t����㏶�0a��&;���P�PnY�6Y�{� p�M�<��w���:~����y> �G�0\��=`�0x�J�N>��c<����L �D��6�˱�$ Y E�B�M��6�/���N�y������$��߀=�����3pl"_��&.�g�=9�ӤdwsowLx��EZ��/�g[U�[ڔ�^�D"��l���V+��c�S&۬D�ݐɈ�nM�R�~
�a��g�8<�]�a ��@H����ڑL&�}���_�'g��5Llnp�t��}a�@�N[� c��Db��B���*�.���׆�W.�`�-R�M�>�LI��
�dB	�K/��	&*��Q�x ��0&'툵:@����6:6�D�c@�L�
83��d� u{G0��� �mj�m��^  �( � m����Y���B��m��eN;`��
����W#V�<`�9,�9F���=����8���;# �6���,w�#'�8������w`�7� � �ڶh34���_�k@���1����]�lA�]L'� xw��w�8oLP����L�h2�{s���=a�ƴ�-�w�wC_ c��M�3C�v혫i��z�G��Y
~��ڪa�KJJ��J%[՝��w�Kc��J-��
�j,��|h?�/+{���x��Zy��Y��g��a_o"��&�zd�Θ�>��^^�Z��it 3aw¬�,ƃ��owfwygߛ}9 ���Rʒ6��h_��Ɔ���-jmI����ư���Et�-��'�T��Q�]M�K/	f�x�v��ba�LL �� ��9*�la4�0,�kP,�c��!�����9:"L��ɲ���.C����� �a��	 A����j�e�Ov�q-��y�U����jh&ǵ�����h�8�u���9�	���̑��> {�Vڂ����v����z�'�B��.�ȹ��YA 3'��S��>��!|���Uy�p�'�w��5��
�}��(+l���A{h�c����Q&N�F1V��`�׮���#��\�*QN*�����/һ�}�ʤ���%57�M[�U��A�0�*0ߔ*�Bؙ�J��V�N$���V��_&>�3G0c�F�h�O�7q���}ʉ�����M8�>�Z+'H[����D^�t"�	aa�6w��Zd��A,6Q�K	w>v8q��߶+٫
��5kV_��_D����R:��a*W�����M�^�Ӫ���K$5u��!YO0[��j$�ι�3 s�D9�1���Q0#'� 8N&�3z8Ppvru(��ISbr��F������@�k�T�}�г�Ӗw��A�w�o�D����>�
��(�X����l�ٽ��x2�o+����J7^aœ<fJÞ��<1��m�W��4��� ��noq���w'�px�ɔ/["�Ւ��N͞}�f�|w����0L�B�::ڴ���̳��z�I�럶ܿm�M�(J��Ϗ�W�摝�~_~W1�M\�E�<_8���=�ұ�7[��7	QTs����W
$k$ʥ��eBD�!c{h��D��~��,�����w�b���$/ `qzk��⥃Y@�]{�}!j��j%�[����[��z����Mo�|��߽�^׾�c��ȆR�,���:uZ��T7��?;���+�y�Xi��/��������7��A.�,��c�B^^��)�tt ���q�Iag�.�R/+�|1 �n����w�;c.���o+���p�T�190��0�K,�e߳���e�6�N�1���_�|��+�݁���k���/H�����{�L͸�\%Sm�Э��vc�KG�=Q�v���X.)��(A��2���!��7��x|���v�ج�I��q��oכ���c"bR�Xi�!?�Ǧ3f�i�`\I�Rߜ7o�5Nػ-7�;��\����p�݉������f� �M1S�Ϗ'M�<��3 ���ۖc���`iG=a�t&�c����G>r�
�����t��h��az��՚5����ި��)M�2]G�K(����5Vvd�ē�6�Y�Ď�ͼ�8�.vDY~��Ks�-2`I����Vlv*�go�Ҳ-��F�d�f�?{g@П���Z���u���?>޷�U�p�~�ցd�������$ f�Ⱥ�.fx�] x�X�N�>��s��Қ�w����g+�N�����>�����ܷ��}�4�t�
ee���)��L��vY;��äͲ�j���z0�8z��m�G^�7����Y�Wp�o�m'�Y3�2�4t�p�o9p��έ��)���90�r��R��J��'qƘm;4par�`��U�i8`�q')xpƬ!��v,��h:�~�q�мf̘�g�'E ��T*���>���~���М�7���&jŲM�r�z�[T���� l��[+m�i��;�ENQ�ض�	�d���,������5��<�cVX0 �M�K���1V�����+v������x�����{P���3���{�t���9�+6������;�>0��uv��l�*=�p��][�>��;f_�K.9C������}���i��7�;�ao�r��a�M*�����r)v\�v�j�oV���@إO�`��ybY1�#�1��<��.��0��8̔k�)1�ơ7op3���ǎ�qՂ�bω�0�R�+J4�B����`� \Xv�� `zY@�܎�t�[&���2O"��]����G���Y.��eĪ��y����Թ�C��{���(� ������g��eK7�]��T�֮j��n��}L�� �΀�ϵ�����x��) ��o�a����l�f��2�HM��g'�#C�K=��\|����"�������s�q�������̹�;���|cv�/e�kNh�������ڦ��U�5{�.��Lm޴I7}�.=��f�s�n��^�w�2#���Xަ�Ɣ�lWQ�9�CD��x��ؔ��31�`�6�`���'59���qm�o\ɐ��T���
ګ�}
��^wۑ�����jI�".������	�1w��G�XK@�Ѩ�P���Ll�r�=���6Qx��tU��Fx�/����ĽB���#x��Ȅ�ӧ�4:��:+��f�}���K1�@}�ԡ��ŋ�k��7����0*(�p�c.TQ�];�\n����M{y����P.��?Nրh`�
��7����6���r]7!vJ�m[C�.�3���.fb��eg�����
��;s,�a�1��@�1���،gv��0�=y�@�����X�Ǿ�@=�4|XBw�}��N=G۶l�'?��?O�B���ןt�&w�����.���T�ϟ�9��V�g�uV�%|��I:�EH�&���*~�6]��
���́6IX������+�x�o
��p��/��?�V:�P̉>�m!:"W�Vsk��1N�&�4������fR#DK.'.�j� ��kw`���s���XQH�#�"�ŕ��������xІ	V+�\���wݬ\n�.�r����^���j��k�+`nQ�<u��7^rPB������`��c>�D�����˯���8^�}�c}_~�
������]:ۋmZ��$��企�lo�lw���-�8raW�tO��33���	{��}q�.A8Y��K5�#*�t�m�t��4m��x<�̏�K���ϫXn�M�Cc�zk��L$ECM�|��ɺc��6�c����o㋽�\�H!| 4c�ӟ�t�W����^�r.�?ĥ�L?��+Lp
�φ(��'��g3o9�5M"&���y���e/�W
'����\S��.��l�1�Mԉo����B3)�1 �d�1��7��v!t��Ht�����������,x��~z��E(������}:ċ���{lی ��u�?����z���*��V�\֦E]p����;kXKk��+u�Q�ao!}�^Lxg`3[�#l�I��[���(�3��Td{q��7��F9:���!�A�n��b�pVK����_A8fJ���f�x��&�3>�M��?�Y�'����p�utDM�V.����/��-�[o�����U[K�:�KZ�l����s:f�)�d����^B�j!�Q�^g#�	�NoBxΛ7/�ѯ��}�帆﮾��0���6[G�x�ސ-I=בI�8Nn�w?����0�܀2��duȜ���w�sO�{ｃ[�}��|��Mk���r`#J���:n�&O�4�5��z�kO\:n��@3]w�F���R�� D��sx	`
�E{}�������*0�_��^�Č���5aK�n�uޑl�7(ky5d����!�Ӷ�5�6�Ce��/m��_�B�AU�Bմ��M�RG�=��~��� ���۫ /�̈��_�r1+f���Px1�s�u.C�����D�_��#ݛ��}![O|�W�Ǡ:��&3Ƹύ��Y2߹nn�t�K��I�q����jǽ����@���Ym��HT�l�-\���;�jx[Vw�y�&O~��U|ERcS�:��Z���9٘!�t&2n�[��l9JYƊͅ�0E�w�y�}B*,w�����׾D�P����c�g�F���1�l�u}�wl� �7���T~��D��H$�Ycp���Gm^;����6��ՊԚn�ȑ#t����[�<\���9mܸ9h :e��
B�|BM��}���q�&�Ɖ��6��\�i�L.l������~��9T���k=>����=��Y+(��Ѷ��LKɜ2e5-_�]���W�6��%K�ӧ\�qc�V:�Pg�$lP�g'!j�����p��
�ūgG1m{���I��]��w���cQ����������TzE�?�0fz1 ǡ��x��α�|g��ګ%?�J!Ί����
�^��db�;�=sĪ%z싏*�ա�mM�|��:��w(�%�?���(�fK�����$�4U�i��0G�2��~�0'xS Lv0YL 8�#�3\��?��`^��	�ZVvA�ۤy�vx��5ϣĀ�R��3�J}u�w[�GoY7�9���D�sò���t����굫�Ң%!D�F0�A9f�Ih1j`�y�駃��n�Pb���g�}v�� S�?�q_	ź)�\��2�X    IDAT@9m&Y`;4z�ZT�ܭ~�_�e��P��L�j%�Jy�֯�R2դr��Z���UM�2K���t2[<�w�;[�ƀ�h�]��}����U�d�oX���۹����-�����@pꩦ�o�ݫ�	�fY��������
�����n���1��Nc6(�~|3�o�
����_Z�HO>�
�|�H8��U�ښU�w���g�E��S4z��T����O��a�k�U��W��v>[a�'<�|�M�b �܀�9+�&H��"Q��b�\l�3�����e��C&|Q����:��>��~ �<\�����}���!j�L�=�#�V�P����r��k+`�%ځAb�o6��/ɻ1���л��J`u�%xY�J�_=N0�jQ�D i@��E�=�b�SJ��[TcC��96m	EH�	v��	�w����
���O���`��'
�=�<���v�>|G�aL^A��v�mF�Ն�ӫ�����A�w��]k��� ��x0���!�mG�kT�p�!ż��n��l���۱+Ξ�#��Z������խ�tF5̉Y�6�R�*j�*V:^�)�*I�%=�L@���U�Ʌ�K��o��P��F�]�>�7laFr��3�-k0�)l��X��vk��W1��躐�ìA(�O>
C�,V�U@��s�νip7�����#7���R�>&�9��чh֬+�S����j����`�A�F4ڱu| �l�6��BC�N��`8��s�	ڎplϘ%0e0�|� �y���A�~~�ew��\T������B��v%��'WS&�Q!׬tf��h��.�eM�
c��1s��s�*��Tcd�l{��cgVe��5��U1��펾��ڸ7���L�;���<ۀ3_��ݫ}��n,�X�Y9%66),��8����O ���Ήw�v��/b������x���{��0s+V걅_R��G�DM��6e3 k��ʨ��j�����<\�dJ�f���3&j�@n.gi�1��v�m_(|�s,��{�E�k E�E&&0�|�6��{G>�]��^��^�3��Z����o}K�j}�@8�zjޜ�T&Nx��� al�8�ƿy����*=����_P��ҫ��p�1`�DZ�P�`ԟ5X8;/��'��h;�'�k��&����%�k�n��>�9�X��oK�͋E�|x�9�C0�Z5�bn�~��h˖5��ra��d�I�|��.ݢ$�Oq�%s�97}�e7�(��^		u����&>>��g�"J;]��Yml汼͢ݦxij��g]�j�h�nWv���y��f�՞cZ��#O Z��Vef��x�j���6  Kq���{��7�
Kwf�**fz�{�$o-_�Z_����uu*�(���M5�;aӃb1����\�g5�ua���sy0}_Q�|�P�����sa�l.K�m��"?�l�!�L���k�{0�T�՜�1�����J��^�rh��v�S�$��ٱZͤ�_���9��[�='��|�	�8�m�2e�~�_?Һ���UQ��8�H��e;q"6	`�A���Ʉ��B������ H�~�,� �ܹs������߅R�/����c�?���h��$s:`L��s�C!�l��_آ�n{@[6W��XJUKV4m��z��`JKb	�e��}���~�~�V`\g���o�|�X=�|����	���N�ݱս��1�}�l+�x%�@�(��\��8��e��M6Sp�:�*���}ضH�0s[��"���2�\}϶a�Ǹ�� c�s�&�zD�����]�)�]�A=���/{g�wU���]g�Lv�UYٷV�E4 	���
QDY�E����Z�B
T�.�V�\�hA\ؗ���$$�}���~�?�p�w&�dk�:וk2��_�y�s��~���tw���m�矡Y'q�`?�g��Ʃ����^R=[��|~�����L2��eW9��,ކ�x#&]�5!��"���� ��c����
pSmyĆ�棵LL���B���;{��%#S�j��$��h4���}W\�ы�����;c�m�۬Yvg{��P�lX���	'�E<|�֭_�j�2��V�a�µ_�:K�P@��\�a���p Z,�����ٳ����a�qx�OX8B(�]���ج��~��5( RR����T�s��պ�y�K��~����������k�<�0 <C�75����k̪���1b3d����1���f�1���m�ɏ���A؆(��l�l�F�G�4p,��F&8%Ly��d� Ą�p�Q�b`Hb�f��6��*� |��q�et���@��������>�a�8��%r�a{fɳ���w�&�e����B��z���n囊�h�:�2Z��/�`�U���Ԩ'��S��L�a�q_�Q�>餓��#E��z�	c+�Py;��
�L��0(�
��, ���W�}�,a�p��kO`��+W=��Q#&|͂�;찱;ވ>۬}a��Ca���3�x�	����*0a�#PBvj�v�Q"��'��}��G��k_��`�m������ �2�����;/�7HUÅ3���s/ ���q�W(���{nծ����9G�e\����^X%�z�T)OR����蜹��mӶ�1��%~5]�6�R3��و��04oAgl1�\��צB�N(�3��C�(��PF���CHG2�i���|�.�B� @�>3�a�� `�=6�iO�@��a#������
8����=ٸ�~���"��T^0�]s-[Ӳ��ۿ�j�&�gt��wi�i'h\���ݫ�>�L?��ot�NҤ�;)6����2�����Q~ I��:�������pe
HiE�+Ű���½������� n�̡d�_�	��˹�������g�;��5�S��V�\��]{��c^�rʺ�'�ˇQ;�z��춗�<�=��
����z�,�a�q-����\�b(
�b/`�-���=��&fl��k�b�$V�1(9+�>�Ɩ9v�`u�����2����e�]�re��~���я�7��=ۥYo;G��dU9�)+�9s� ᰅ.)쾙y�[���� oW�3kq��<q7�.�38b*.�v�7��"
rT<�_���/ڋ~9�;�}f���"�O� ?���7���'��nﲱ��6h�͌��f��\����������s��v@V\����3?��Q}��E�'�/�×�Ws�Y�J�~���u�u�V&;U�/�V�L�_Ŧ�����BzA�L�~D[b���7�����v�ϥ���'�0ǹ����d��0@�X�zꩃ�`�Ƚ�,��(e26�F2*�q�\�*����Ύ�Ps���c
�u��v��q��ÓڟE��v�駩yBQ���*��I#Q���q1�:��RlmF �hX�?��?�O~�q��!�j!t�q��^��,qA��dל'��]c�� �(uU�L^=�}��k��C?��{�����N;３��J��K��UTU�h� �ʑA�<���A�ƌ2�N���%�ڟX��1�C(7�I�7�.^C`�1a�1ۦM}?�^�H��}mⰾ��Ô�P�d��z�Ā�
�����L@L���sx©\�� .�|�O8�g�p|?���>�)�Pr�ʗ�铱yy
��%O�w���f�����|�9�M�бZ��S��7�S;l��.����^*3�5j*���U�JJ_���46��;��oX�SА�7}���?���&������:+�^3ރu���$���+�c<���8$��n��,�J&i��\������c�S֬^�V�=&�f�u��o����/�Z�R))������U`O,'Dc�}4;��VpPRL��ߞ��f)o~�C�0�0
������0�T؋�,:8���Á0���;�OިG��c�Ol�[.�|bX��~�zzra�rEQ.�}�W.07�Gl��ְ�?�{��� ��xO>@ȏ�c�Jf��b ���+ء�g]yW!F�%9}�=%��c��+K���Ϝ�����9�.p�qh&[�z�ސ�5�VZ�jc�}�Ke� 4���Oq1����\!���I�FhP���I�� ��h�%������jG\~�_�z�ŗ\��=��&N�S�_y�v�c/��P}��W�a`ja{3?1[��#�<*(y��ؿ�����%�I���<�`�@'g͚�@>L5�#��F�^��1�`A.���ųY�C��|�� �7�����pјo�s�k�.����������O�v�q��o�;�����Y/��X���
:�%Y�d+ ���"On�<���qز�\C���?�?Z�h� ��� R ���9w�DҮd�)��:_O?���͘��}��`=�||���=O��#� �`�3��HU�6w��O���X���8����钂C,`��Y�</�{�_�Ťe����=�ዑ�a�3#�k���LPқ�2��.3.o}u{��i<D��Bs���t�<�m֍�:���c�f�2 /����\��szn�
ݵx�*}���.]v�;����^����O�G�L��T]����w��P%��l4 /���,r�&�0?�H�͐7օ c�kƌ
��#���w�uW p��6b0W��3�fԮg3`�o"���cH �9������Y�p�c�S:�_���uDH�md�� 4���o9JG��Z�t�{� �X)�rc%�o[d�8�@���.=�oߏ�8��E9��(��Ua�U�e|�M7�ϓ�yIa��03a�>�eg�������J=����y����?+���V�\��k�aa�Nv1��9M�����#�ir�O�Y�Ȍ	c#135h�l֬8��oJq8�L��w���7��>���9�q7w�~t� l&N�!��Y�S�b`��@a����j�fo����6��9�#m�� �������)�I�ce��ιD/�[:C1᜖/[�;�r���^��Vt��gjC!��������SWW���˴�A�+�e��9� ��I55)���E��ǃ�K�/�����
� w�_���<x`�?���y�I���FF�����t��4�����>#���;���f�s�7^0s�̱ˎ &�Æ�wf6�=��OkK��e:٫v�NG�F��k���\��6���n����R�!�3tP�+�TK;��#�p���*��=��u�-����}H�'O8Y L&N�m�?��{�u�&��Q��)T�7i�ҪN�s��;�Tm��N[&;b��M�[�|%����o:Oxs'���u#�Y��8�O#���I�m�q�5f�CńcY86�g�0��O��z9�K��m����7֛8�����/�F�����\됆C^���q���G�����M`םv1 0p���} ��h�.��p�ւ��+V�+�~I�r���}��Ӗ�<VM�eut�����Z��_S��	S�U���,�ǩQφR�6.��4U��m��c�]j|�f��/�8x�dE�u {�Ћ�>{�t4v����"xl~�z�9k�!���b�.19��d�{��7�o�AxʚUw��&�-���}5��4k}�:��N:�-o���3��E�⣋�披EpD�)=Gp�!:��3�;wnȂ`Cq��|�ɧ�ӟ�tp�H�p+�I�r��0�es� ҡwh�6���ӻ\'e��W�ӏw��9�T&�٬Z&	\͙�A�{)�gQ�:���ູ�	�q{af�N���� h ��w�@g]2�3�t@����e6i����~�C#�g86S�-��Ôx�/~����Mq�3o��
d��q,�m�;��o0C~�g��]j>�����=\u���𙋔6%,�nݚQ�0�E�s�����+�>G�N;^��z����Fmmؘ��5%e���/��T��X�J99�֍�a�.eI���O|�t	9��w�������B����c����c�l��Ϙ�a���Y!�l쩠���F����r����d�)f���RO��CY6�N����k�����;�J��7T �Ӗ����i�v־�N�0��(尢�` �Ap�k����i#f�qY�$��u�[Hb�(6��=�"V���cΓ[�0O�֮c�KY�|M���6�j��N}��VwWC���ҬZ��Sg�����G<����H`�%��t��"�}��w!%��x;퉶��f��JG�'�}L,�cc���ص
,�F`K�{O�7^ȏ�]�!@ ���3���6
���33�o�_g
��.�E�c��$F{ i�0�z�F�s�{�k���X����>o
��b[��1̗ԁ�A�ٌ��|^���e�F(�_�k��x���d�IH!,�LP��I���V4i�����!��d���,+bۤ��xi3&�Z04ȋ�g���%F�c��� �C=4Md�z!�qhgz!_�1��p�����0�_,X�1a�&�_�#̄a� av�UJUm�������w���	a�Pv��k7�OO���"[�j�&�$��L���7�'��d��n��"A�ܩ_�Ǐ���uji&e�'1�f=����8�jU���ե9'�����;}�e�-�?���:-9"_� �d��;2f�G�v㝞�1���=:D�p�ͨ�<Zy�G&6��
&,��o�Hy,#/�!?��b��1Nڊ�a��nב���gB�v�����6�@�#��i�`����y�Á�#O=�yµZ��Ld} '�Kjd8ȳI��6���4~�P��y����F]��a2$�!�D(�Fǲ t٬;G�;r�%B�����i�����'�`E~ ��s������l.�8��
�x��ⅹL&�ʂ��p���f�	s�'�lM`�J�w��p�*I�C���� jf΄$��F�q��V��8�Y�cA{Ų�U�B%�Z�[��U.7)�oQ��S��B�Rk�z�f̜�l8i#Y���{F;����GNL�H��zB���8��8�h�06ncNXw�'���X�F�n�J�C��M`�Lf�D�5XY�&=�3ș�%�IL�Ek@� I��A�n{�6�a�� Mϓ��� �/`��C�m�	���%?�qzz��}�=�\ߡI��U+�(ñaY�T!\פ\�5��q:;�7̽z���0���f�p=��|@�= (�A&��K"��9|�3����f!#dF!3���⸱�o&< ��]s�5�9��~�m��#�c��<�1��Yi�K�"����PP*�:l�	%wƅ]���}V����|��SO����5���W_O.�P�\��+e劍~�s�Nꡪ�T8�O���0<n(#��$wZ��*��s=Gۯx>�	0������*�0ڶ�~����	�X����X��۸=��i�=�x���quH���L(�{7 Y8��3&�K0�a�a���c�����f@x�[Lyi~fٳ�����b�Z��U��J���y�T�*[��n;k���z�31�$�!��/��!/���CQ&�$���ymo	9y+�=a�4��������2r�VlD���=�=�rc��o��׭Y�^�=b8&#LO>[y�+�1���H�z>� ̖�.���0���v���K�A>V�F��J�[?�����g4���<M�d��_�bq��J5�
 <�Wف�ԯv���)!gLw�,�r�b��X����)�Ϫ?���c`L��~k�wS@�w,ް��q���F/�ŋ>gB��8��	n�Π����]_<�u�>�B&�P�<�������;�._�ܨ%�̼v�)6Ȏb�˟5�{zU����o���&�+����/���=�~���q� ��,�}��I=��2����EM�1����X.C��-�{�<��X/N�����j��L���P�1�k�\.��k���1e��׼����7��0[Io�$4 ���%3;���@���Yn<��3:O,Ѐ�������ꓢ�#�F���zC%��S�}D-���>E�>ݡ/����    IDATJ��y�W����5�a�����CHt�3����"p�PL��6�CyE[
�ai�	ב�t�K�c�����0D��`��&k�svv�x	��p��U�gx��Yxy>���x�;�`�}�'��X���W�?��7� ��8cǼ ������M��,��dɬs(���ҥ���۔���ڒ��Kޥc��3�l��H��/��Tn����q��T3�e[�� �/�^aQ�� ��`�l��cꐏA��3 �X;]��}޸C�A�`���M8r�ܿ]s�5�" �V�=�U��1�d�cR�Ó�V4IKv���`�.XZ�ce@x�u�Q@��;Pp��k; �"Ύx��������zVi��NRKKU}�u�x�����is/ToO�JՂ
MI���S�j���+��&�{^�1a�U��� @�:f]6�1��R����s�����>�$�[9V`<��3@ ��������	O ��kv�N��]XK������1R�.���j�T���g"//�J 0l��Y�">̵,���!���{��_B�rZ��y}�/*��Qss����<�:�8�8�F�e'��?��ϭS_9���I��,+�mW���z%�}�=x�v���]�*\����c��A<�D^�C�\���z/�ǀ�^�0y���^�ך<nc���l���]t�n۽����K ��J��Ϻ
���՗\[O�TS�x0cv�'pz���y��E̼�!\����f��ٹ'hF�u��O�-�f��:􈽴��U���:����vMF�ZS�X�f�</l��e9$���M��1 �S��
��-��0>��/v���r�7�o1�<����I����c�����h����z���AO`������ ���y&>�矋T1o � �k?��={y���e ��s aV���qX�g��1>���%�>�&�՞�e�� �r�*�~ۗT��W{[Y��;4��7�ؔQ��^������|Z�F��^��]�ϵ�\��X����~6����#[ד�m��蓳Bb05��`�޲u���!�� Ӎc��t��+
�ۮZyW{�/0a�3I�0��3�cf��'��	Sw�k<��'���v���oTQ3x�%�8C}]r�{��������U�/=' �SOn�;Ϟ���R.	�d�Y�}���"Ȏ0�e<6d�ԯK+��(��`4���c,��cθ�~@hF2�c7�^�3�T[2q��1��粓
0!�ҋ��V��d�� J��H����� ����Ʊy�c����r��llr�E���DV�1X��X�c�5^$%"a��8&�iC�ӳO-ӽwߩr�[���v�	�J�O���[�U������aG�H�}��vI!�I_8���k,��	Wz�ƞw�k���C#q8��3����r1�dan0�0L�l�\O�v����t�A��wbS f&�8��<ǩ&���	��H.���C�/�ȫћ��_��~��������w߽�rEI'�:G}�mR�5T|���'���f��ˊ��qrR�; ;����d'�V�t��bH�hDf�V��P 3b�,�|�&쉵5r�{	y���[�E�����D.�8}�3>�6���͡��A/$�� /y� �]rX4��&%�6�� p�(`� !lݛ�_5�L{�U2�rZ�r����ڰq�&���kߧSN>>��-�����2�膅�=����4��3�'dP4B�D� �Y�Fr,�'��=`���A�u ��M��rp�����.}磌�:oLO�skW��^�ga.�?c&�UR;!m=���غѱ8�.fR�	��|}�J������
<��0�E�;�Zx�U��#�W넒�|�Bx��z��:������)�[��S�N'�r�^7� ֆ2��D�)��L�?�{~6l�9�W�c���C�n�l ��Ӌ�2 |f#�1�.���a��O��X����������C����0;�`�;��da��o&?!<@�����=���;@����p�����l$!E�8mlH}dǨrz���oܫ��U�<��˯�K�4�Xm���/�F��2���?�j��?a�J�^U�%������4��Ĺ�c�A�n�����>�(�XZw�=��c]6��׫����1a�-OzaL�s/G�Y���Asw ��y�o
��~9��-��CV�pލ��x#?�e`]/�s]�n��Z=��O�������ߠ=��K��a��>����ʩ��4��P;��SN���,Ւ����WyQw��^�0X��D+}<�caP�X]���+q4C�#f��9O,_?�e���;E&L���a��S����v<�� U��,�x�Ӽ!�qd�7��4%�IZ&�)��8�J�:�@jZ�g+&!6O�>�\�l����E��|^�ƕt��h֬7���G7��	O���>���w����\PWOg�?C�B!�$���nCb�6q�o8=2�ݔ��a3/��ld��%��t��\�y�r��.\���1-e9����x��r�aÁ0�����]��c�A72�'��C����5�\�x��B���3�v�i/�	�n!1�Z���?z�j�U:�o�g��V�g�u�POOa �{>����C����B��"3�E!t<����d�Z������G��ً�+�|�p����Y�B�	�`FmX,����E���/�]�>��t�� ��<p��ɒ��]�B�qo�u���v�����'ǁ�qg5��|aT��w���s�m��oPss����b�|��d������?ޭ��Ї/�V�f�l�(4)�M�- L�i�6<V��i�I@�8{����vl�z�U̃o/\��}cz�F8����{u:V�'LL�ě5L�T3b3��:0T�'�n�y��<���B�e�|O��pD:&��S��>��oi��:�35uj��{���ɲ�<=b�N"��#V�'�3�z&��11f��&�P�nk@m$�{Dą�o'��<��f��'N.[���]b�.a��a����~r�d�m3�r��a@��7�:�d���=�F�v��]�)� 2� �yƄ#	��|��9D��C
��.yN��M�z��Œ���/u�)Ǉm���=��J=��J��4�����96rp"M���|���a�� �##�����66����8��a;�wa*/�zm���#�s�ܷ������9�~�u���!#�0����
��������B���=1���-O��@`B���cP6X�r�7����8;�q�
ɰR�Q�nפ�vjҋ�*��W[�6z���:�����ʐm��:��5t��yz��
��$=-)$���y,�x��A�1 !�ȴ���X��.��G����?ވ3�V۸C�gs�֦&?�u.�=�V�3�+�b�Q�7Ġ�^F�x����D_��ec
�dl���8LF�_�%|P.�n�;�q�pQ߂����K��2��@�*��زH�khժ����I�r�&L(꣗��S�E�:E�
ji��Ξ��[�J�FA�-����W1?Q�|�*��"���\wi|���3��u�{\�1��I���PQ���qaH�C$�W= �ߢ��A�����M��|��g��eԎ8� ��q5�#��~Ǡp�Ր^cpuz���t����W�bBL�=�0�p�����3�(ꌠ��Y�����7[4O9�A���a�TQ&ӭ^xF�dU�_�b�-Z�lI7��yuvV���T�t�����9� e-I�ګ���|c6ʢ'qa&w� ��cm� 	�2i0Ƹ�^�J�Gb�ǵ%�&�W���'�}<�@X�� �	@;Ǖ~`��k���o�8�.�@�g��u���ʞ!l���dC�>�o��!D|V��Yo�c#~�K!�Ax��%�p������>�zӛ�T�ҝę�ֲͪjm��b�8���a3T���ib�I�=�$�h��6'�5�c0�G6)��qp(Ƭ�G�a����wv�;��s�yޥ�N~q�ɍ��=�]a�!�J�,RԪ��fL����>v�hs\T3$ǁ�������Xx
�s=�q�|��'�|������S��T�{����˘�(G����xw��(mz2�uU+�����]}}T���">�RC�R�::9i�|�lO؜2w��|�5a��$�$[�_�?��qYD����4��e�͌f4rQ���opӃKY�
e#`#k�7�`$wכ,�61��G�"�!�`١�a!l��6sX;��l�� SH��������~y����Z:r���;�YI^�p���"}�Q6TQ[�b�����HU�!7�6�O�m_ԥF&�RoQ�ﰫf��&L����B�����dיK�z��c0b����7��x�	�S�X�d��xa�s�%�����H�Er��k��g�End��0�T@�Z`��{3coj����L&�\8�Lxƅ�m�v����(`^�6�s�zM�BU3^��������>!� �ԧ)�H�Bh6�Bz�:��@3�u��t>��yw�q��������PV~��o�&�0�c�9F���g^v�	�cZi�|��!$�У�>�Ro�����^M?I=]R�i�*UJ5�l_X��{�ٚ6m����X쓣�^�?6`���DQ`�;p���w��h�³�*�(�C"f��-�4@��|4��^ރ�xLlBo,|yK7zM��v`��d�9�� ��3���f `��9 �x<��x����`D�`ڃ�nX<�ט�,}��{:2�#�>�;ݭJ_�*�t��U����q�p|Q.7A�}d*�IS&�yCK�=�s�0�I�tE4�O��	�����a̚����� s��� �k��
+�'�`�]�ݞ��u��`$�4���K8 f,h+����˵�^{ј���,j/��p��b�®{����6�Ӳe+B���h�M�K�@�J"4�]g��5 ľ��m�Q�N8!��}�����gs��fፓ5p�-#�;��#f��3U�to���K����~�Ҫի7j¤mU�g9S$Z@x��P|>O�N�}u�178%(�A���j}�������|� �DcB�v4�Ǡ�c��Z��L�/nͻ�r��8%履�#�it]d���iz�d���M�H��C�`��9o� 0I�7��p����w�6��� �P>r�^.�X'�����%����kɲ't��U�mRS��\�W�ҋ��-�*�m����@esM��	ƫ^�"bF�}�P:Y�\�+��8:��@��tµ��r�[�s�}�7�ac���H,3��ZF�6�`��]�1K�����1�e�Y@��c��_�hۜ"��<N�jV��m:a�����{��?@ؕ��xfE^0�$!4�±���㸕'2�b���s���(�u�]����x�_+������ٸofo1��چ�*�6�_�s�:7vJ�����sEe�mz��U��[U�$i4� <}/��Ձ*jM��R&l�4�dl��3�2X�<�1ak@o�{̬�Έ�7���x�I@0���ۣn�;�>�X0�	�9�H��l	t�z�|a����:˖���?�i Y� �ș�p-2�~�=�;w�0�F�VM�
��f��UH/��?����5�vJ�JI;�8A-�R&�d0��8q;�|���m�}T�'������{�9R[ɰ���y1�~;���81���w������'�3�� ֐5� ����*{��g�l�����³����p�C��[�^��r�o.X��c�SV�^4%S �i��9c�~�5�Z�f��z�i��&�B�*!�3�!�V\��N��� �^���{Ă�"�&9K�$.��<�����o���ͼl�`�����o�)_�R6ӣ	��U-w�����{d�.��@�	��4��>��|~@yY�|��YO�f �ǘ$� ?('���΍�lDc��g��@G�0,���Ys��Ѿ{S���KX��3�&��	�sl֠�.X3���C��i���y �s\�g��\W��0b��;�U��)�#1��K��60�'�zT_���j��j*J�;O�f�\�B�v���ꮄ�����h��ev�����)��2����A��L��+d�gȒ�:�$ ���y>��@,���:gW�5��N��^̴�y>�s �{�'`��Q�V�����r�!��D�6��pso�A�����+�SN����_��~ul������r��s�(��M����(X���ٚ̝o�2���!��8���dG���e�	i_Ҷn)�N�nۢ���ɒ;ث���z��:y�{��פ��j �,���|.�W���dDff+�9ed�����-��a�5�y���5�d,y?���y�=*��h�vS�g�qYЁ�B�K��d3��j��/בֆ�9����@�(I��x�f�qxs0�����s�s�E>/p&��49�Zn��g2";��/Q�>M�ׂ�.Ҽ�OT��Rؚ[����auu���P�S����d�l O�s�v�X!/�
#�#p��=a�#�u�r�l����N
�x3�מxD��.��&����7^�䏐���Z�V���},�xLA��)/>������B1�r��ݷ�U�z�;�b�Z=���b�1~i1��Sh��`k'?v]qP*,44�ů��\���Ș �����Ზ��<I�܊��X� n�У�~����L�)sߢq���j�ji���U�o��j ab�a��K��pD±��@�UL>����B��N���l<]d�c�:���3y�R��}���� ���@!䙢��a������:�݇��aa��88�y.a<FdͶh{0~;B��q ����Hy�=���l���m>�b����/�V����u}貳5{����e���o~L<�f�8R�l���
;�Z!�̚
�E�O��zǜ�l,[���!�����!��v�w�y��w�yg��E1�1�d�<`������_��R�����{'��"]]�֢j�|���^���1�k�/������NJ=h�:�y���%O�t�#�0�!�Kh�]4&�Y�Wym� �\-r��c�y����F� /l��o��E��{b�P�L8��V�z�_=�kt�՗��g�N>�X]����5�G���y���E5��x0�/��9]Ӧ�|XGxɅ{��0�J�Γ�c��;��Ŵ�ٶdru�W��Qy�x�:���nh/`mjG�h�e�r�����β��i`�,�՘�S�(�ü��0�a8.i�-�0a�8���c���N:d�35�����d���Z|םa����U}�w�3���?y@��?j���.�kM�v��բ��%�^V6Ǯ��td������aLa���1�<�G�Kb�,ԓ����O�!ț�8)�5�9��)������Ż��l/�﹖�ID t��3ٺ_��j�|��kn������o���ֈ�5&�Z�hJ�q ��t�̃C8��?�ZK�?'��BH�0�
���;n��P����.��� ��[ɉ��x�A�l�@ ���g�pPZ��������p/��@���(p`x����_.�u�]���zXS��붯��^��nz��:�B�F�\K�u��9�����d�k>ʓ5�I`��} ���zP���Xm̈�DF{-�i��88�?�b<��{<�}�A�߱[�^�L�O�����[��v/��3& O�u�sp~�Cc|�gH�&�5`���x����yq=�0��L�|���-c/�� ��X�hb����V��oUϋ�0���^�N�|ʛ��]�5�������4i����G�����U.OvUF�ZU�BN�P'Y셩k�I����J������Z�#;X��?��p�����xA��~ثpx�ޅ�:��K���݌	�;2��}q���E��W]=L����~h�I�W�9��H�VUԎ8�0�t�,���/�n�ZUJ֓�5X,2|2�����ut
A9�������v�m�s^q�3 �-oyK h,��,>���0g���_�u��9vcE�qa�sl���S��c}�n��:=��o5~RC7�C:��Ѿ�q5    IDAT�uݚ5���4����Z�"'���	�MQshd(F2�Lw����l(��y�E]|��~;��+06��\��㉀m�B��G�V�5}��I�3�aY��x?� 8��6Z�M�v�g���.f�<P%��� ���qȇ��0ۀ�� �2�ŋ�[�+᧟Z��~�N�z7h�Ć.��,�tқ�am�.��=���~�}��_��4S��b}	0��/���<�f]���g��n�A.0�P��s�f, Ɛ1Ǔ�]���3�y��X��;�;9���	��������6!W�AX�b��֔����]~��z��m[�#֯�����P�Y�����ЬYoӯ��־�F}=����D��d�B�,OPB,�58l����ɂa��
�����{  ��Ib��(��t=a�3a/,�)�ro�nXx�~�˟��Cv�?|�Z�v�]�?,�9�H��Y5���
�e�� z@���F�1�RR�g��P�?i��f��<�q���s�ꭝd�N߁�X >c��ǘ�۬�qf���f&���K_gC��5{"�`e=�6
�k�x>���c��aWN��"`0��.�,�9�3�7�^�Mf��K�¥��\sD���"+��a�n��~���+��[յ�M����׼S�g�Ύ�n�����>���t�?�LW��)�Y�(�YQ!�{��Oh�e�¬R����w�;�l�r�3�����_���s`��#L�x6^��+��m����Q�QJ��"�E8��R�T-�͎=����ի�l+��R�QML�p��5K��G~7��!�����e�QB6g�BƲ $���_���+�8��ěY���e�vBA�4��+�NU�~��>�7k�LC}]���+�ѹLg��D��]�B�ӧ�\�s���[WW#ۢz-�l�%���
l	0��9�h���Ō��,�-�}a���e�¦fh�@����� l���^�ݢٟ�x8o�+��8�c�h����6Hq�G���{ ���g�5.$c��
=��X@c����3/�CΗ'���x�KtP�}{�<q���sk@���+���;Gtj|{EW]��r��[�������S;3�����}�6>I'$5�yT#S*I5$!T�_W:s�~�h3��
���"}�c҇�c�`��@5A�x+`?f�� /d�����H[�$Ƙ��?���z��"u�\u��fG����z�0����^����[&6���ab���7����<�(n�­ fC$.�LV%�w�:�zK"ʉb��0���IlwvĐ1�lM��F=��/��n�5c�.j���J���/��Yg\���&�5esy͞}�f�<0� �誨�Y�A��O6O���dw�w������k6N�b@J�S��H����i��h(�m�=�Ѽ�F����1� ��?��\�F�UG:/0D� �\m���p���w�AR���zb� p8A��G�M���#��Kw��ԳO讯.��\����L�r���e��k�~=��M�fg5�L
�*��Z��ve�lEO@�m��$-;"��q���n��"�	P�Ff�;l� 6�,R�LҐ��W��8��s#§n߃AMy8����1jGd��o\;�y�1qՊœ���j�Զ�zӛ�ӌ�����Jk_X�r9�c9E�Av�項���a��A�X*�j���b���ISC���$@���Q:3l�-�}��/+xb����j���V�.�L����׺��7��?��9���֯���mV��JnA�O>}�	'y�c�3u&���m�c �Cf�q��,4^�Ќ�6�k�׋v�o`6 ���e8��6�n_ړ�e:�$n}R?$�?cc7b��È!+Μ ~K|���`x '!�+@���6{�{��\�Y�?��p�b�̛0 �}�7�K!=��?[��.}*d'�<R̕t�U��ig�Z���T&�$�V�Xޡ	wUOO]�zN
e��jToY�<��x�7�����S"�����~7l%����L�!�a� T���K�"o��%�>1n�'�
,�X@�@��6n����������������ï������J=���1�L��M�Wo|�B��}B��	%g`mM��v\ǹx(�! ����ʧ+b�Z�LB
�\rIP0@څQ�Id��0�aet\��*�'z:~����R�Ӓ%���)�L��j�S���YU�7�����%G�$ LLx?e2ĞQ�х#b�f�]f�˓� ��.��l3�� �H��u�&�A������4 z�Gz�pߧ�f�N�73��P᝭iG����{b�3��x���a~3����N����u;���E&�8�Cx�� ��P�Dr��)����D���۾"��j�Kg�~��p�~�zT�R��MM�SU-OЄ	����������JT-l
���-s٘apDGX�!�@H��0^��g�&j�xӘ� ;��;����P�u#֙t+ި搩A���	<�ZO�����|.��k\;� �M��řkon)fX�ʔ� �qo=F�gLӒg��s�%q&�h,�`�B�3������2�ʈp�^\CHdF�
z��w�+��Au5,��7�blN%��`N��$���l�G~��֬^���^57eB"�fM���mR8����O �IQ��ד�)UN�3c
pܯ��-����l�l�=q�y�-\1�؜��k�kE����������h͜<C��t��c������
g1�m���/\�3`d>8������8v�wZVl�^���m?�c�2���z5iG���u\U�q���	z�Q'��}�s�������|�/�-�jo���W�#�X|���h����îC�+��G?�YT��a0���q��
u���i!��~�7 �aT���F.��Ƃ�_&<y��w6uo<&�Ԅ�i��l��O�*��]�b�։N؂��C[r�e,
�c(B'��vĖ�g��F ��=B5�5k��G���␄]A��1c�|*K��/�鬫Q�(�k���Y�WooWOR�2�d
�,��Ve0����&��هc��,��@y��o�'^��A(aČΟ{1y�/�,;������K �1�JV L�P����F `�O?�ϙ;��Pf�\k���/f[3�	��e�t�w�^Ω�H!��IA��6�z-��	���λ*_�T�q!Lx/��7��$Ԓ,&����|N��?��C���� C�ϟ���7�8���>��]���ο�R&cY����Nj ��󦒚��s�V�5�-_4���V,n���/d3l[v=�Z������POx��v�c>N���q,��1+�)����)1+����b���w�3�����Rc*y��6�%`pI�q�%��%1SE0��>�J?uA����
;x
M�/T	���Y��e4w�;4m�tr�Qݛ�~c�d�n]ş��nc���$�g�y"�8�~����������@<;�=5��F �����t��t{�S��g2\�m�G���� �t�R�v�"���.���p�Q���zN�B�z��!U���M���ڦJ��l�d�0�6'ٛ��x�,!�]���*��n;��a�=~0��y�w�DMa����xC�C����O�&^a�\�r �X�`�+�m� �dGP�'��ic�z�
Y�f���Î�34����+j! ӫ�\� (���z��ư30l� ��F�\�s���t��H�Â��f��_�������~WϯZ�lnɅ�Z�z�	�k��+��g4m�~*d�����3�<)=����%���qB[e�E�i�,��ʭ���{��i�|����x-ē��[k{w|�%�7Vc���U�v��QS�ګ�v,h�m�T������є)��cުw�C==���A�b����?��N��$d���u��s�v
X�6`^�3`6[�lp2��,�9�����kh�: l��^t�=�1u�w6uw�*jo�7z��ʚ2e�`]���mÎ	z�#P�2�Kl�;Wb��5a�7qa �;e��c��x1�v��n���r�AZY9c�^ߠb�������.��j�z������h��5��B���@8�����[2	�p�7�xW����t�3��dY���n��|�pO�������:	�^�	Cz!6}M����Gb�[�җ�
����������ޖ�{�{�f�~��>1C8Y�V�m4�IjK�I�ĳ�����m�x��/,@�M+�i�r��y�� ˜!��6b���g�p��3�#�Q<_�y6�\6��k�9މ������"�1?Y� ���yD���~Rq�"��gB5��`9X��2�@30�
O�1+-�5`L�^��B��Ya�X�W�z`�@�X(א��A�q��j��B�G--%m�C�
�%��_Tk�=�h�N�w��:��6� a�{���-�� ;�)F|n��q`/��13Jjz1�qrRr,� ?�	���o��1��� �e���L�8���[ߺ��4�|�Y}�+�%�|����/t�;NPw����W�>A�W�k�z��q�_X8�r��y�>��Ǝ9�c��U �f���F�����-��]�q�٤Ћn�1�@��;�I&;�:xŏ�׸�QL|��u�]7�g̑�6>"��5)[&h� �!}lZ(��8o��6Q�v�*fet� �n�]�C�>f̎�2�����ư�gN�I�A�����ߣ�v��c�?D�'��W��%%�q����*��� �p�ys�־�NW~+@��:�	����)1hDS~����7�12�j�1&�+��gZ���u�1�t����X&���Z��}�/�V*�������9��R�K�B�~��r���g5c�#��v{�^o��J�.��pZ)j<&�s&f�7h��Ldg�6�ۺm�p?P��8��Ƅ���B62��z0���]����F�]w�y? �㫥#�1;&Wj�c�=��8�<V�8��t&[*���3��}�N*O�6���1U�����S�A�v 뵒�}��Q_�����t�E�PlҳOm�ɧ�'��Y��Xb�[�^���:{[��e���Id���v_L3�X�̴=F���Gh����J��h�����C��بZO�γ��T�q���;��Wb���K�<���z���;5eJN�~�l�r�q*�K�����>v��Փ�G?z�f�<T�2R� 5�pO� �d�v����������Ƅ�ޞ�c5�r�5evmF�8�1�އÞ��S�����n�a���O�x~q{�/�0g���#��bU=9,�Vāp�q+F�:;ǒ� �w�xq΂��f oK���ټ�L�85 ��1~���V�ʽ������k��L�?|�cz�k_��˻4��w��/�Z8�4�rν�[.~iFb�ܰ1����w�(��!��x�c`��bO����Г�x��	$6��+1����Oa�e����x^��X�����4����X�z�]��٧���ޣ���v�5i��iμ��S�u�~B?���i��]4���{����2A��^g�_�<,5�qK�����):�T33]�nM@Lr�W/��egP������+^5��>�ûW�/��2��|�n���X�%sj���x���'�yaq[����ld�����+�����]c�Ke`J�Y��mS��O+v4������|f�EV�~q�>��k�裿R�(}��u��k��>���3T�4��9r��	N�7ڼ�5�@��̀��`�El�����ld����D����X��(9��]CV��Ɔ�-v�F!fk���EX?ӆ#V�4��;^��3#{Kq�ʆ����3���I��x��A�Y�����8�kƽ���i_3;��`{,c���X���G��sZ�d���vU�]�0��_v�N�}�:6v���\���
m��>��ŗ�W��-iܸ� �l�pQw�0;x��զ�U���Fh�~m���Id�\{%�����#BRvt�m�.�4�7wЇ��wY�Vΐ ��|����{��K^�G�_{﻽��Wk���ԓ���i���R? \�	�dan3JY����q�B�Vi��̛,T���꘻��1���d�=��1�1�z�!FݴR�3��Y|<��p���%6i#3��6ǋ7i���5����-�L�c�g�n����ux��������Põ'f���G[z����%��J����t���ּ�NPWW�>��O�ޯ=��^���ϿR{�}@8���4N� $AMn�W��u���A�����i����:�����%�S��M���'��^:�o8�jaœ4�vK���{�b���S̄c dW�po�.��|��kt�st��ǫPl����Yg_���A�>m&<��s� 3A�v�?n3���bOz����eo�@i���ǆi�g 6%��@�`�4;����wm,�GiZ/�&����u�q��:.���ٰ�š����H��c���4�r׻<"m�Y����f�Eǲ�Y��ѭ�W#ݗ�OCK�-��E�T�/������Ь�oP>W��zH���۵�#��|讀1�p�Q�?���4��$���s��z�`�n$|����0�Ɵ�=��0؀f���&��f��N�'�[��:9�Տ;�g�Q�qU�+aO������~��ϴ��4󀝕-t�l�������Q�:Y��,���ԱH���1� �l>�<.�9�k�� b��y���n=��o�(bvf٥�ᦔ5f�1�ĉ��i��������b&2T;�No�u��Y�~Y�}y="�$�%RiO��c٧��,6�d�I�e������D��!3����1��Z�sҞdl��bj[<��� �|ų����]Մ�y]qջ��YGhܸ�J��V���������M���z{)yYT6_V�ZQ��2�$�K_�� � l����H�X�{�P���5��_�翢 ���r��ń�pD�CVʴ0��ck���1����Daa��V�� \��Զ۶i�]�iC�RU���6^O=�^�x�ձ����/�0�-��>�p��@L|( 5Xx"yU��{贗X>�Ryp���'!���s��k�a?s�v��4��[����e���������:o����>�}�����C�q�؀�k�f�#M����^����Z>������>���Ǜ�x�J���,3��3����� �ٚ��x6�`�Y����>��$E-_(�T�	�w���=ڰ��9Wrr�1���#Y)S+)��6�H�9ֵ�H�H���M��Ga6kLY�zq[����@��t�l�(�$i �d�=#	j���<610��M�tJ�����U���d��Śr�>���[�yd�>��E�x�z��ԏhd5w��6mor��c��L�>�x�P�|S���p���"fαu
�Gb��.i���ń3��3hx �gg`����(1�1�4����)�!p��2`{\b6��}p8Ǚ9��a�5�vJ�A�v �Ά�����:�a挌Y�w���<֩��7��/�W��'�I΅���4i�8͝������Z�̙J�) oK�d��m�f�LQS���J���`��{ｃ�ͦ͞�B�)�wsI�����ޡ�<_w�u�t�Acw�\r�|z��FCeGp�=B�W���c�.���IY<!͔�(����Rw������a�������h�굡�i>WRSsQM-mZ�zcP�z��l]n�5wΙ�6}/re)�	dN_E-f/���7{��pb���}��J3]?�{CM�l}�(i��B�H(Ļ�x�����c���H�����H�7���oo5EnT�Q�:v7�vV���En0v ���N)C�.��i��R@�<Q��=���cEǸ�]����x`���Q����Cޜ�g\�ߴ��
��g�����/*��e�i����	7�b��PO���,5*�8��bSC��^�s�j�U-��:�����k�T���G��H�.��L(?��J���P�O�k��M�{S >�}t�s��B���	Xx�x���E����\6�"@t    IDAT �< .9�03-����SY�z��.yF]��SsSC}}��+W4q�d��Sn���
R�0�����~e�y L��2��� �!�%Č(�$b�|c@
h,���D�aƘ]��9f�~����� "��ras���K��ٟ�/n k�a!ŏ����8�m��|츞�r?p@���� %bx�Ϻݱ��?:D�U =�x�ϊNS��
8s���T���=��C������9I�q�Ɗ���U��<����̌�p��b8oh,w�g% �U�G�r_+��^ݠ��L�I[��TTSk���k5QV��ZhVo/ۍ��q�^�t8�ۃ1>>�}86����M��?��I�qɺ����@8��|���ߘ2a��<��([��B�0���I9A��A�cX
�,�5NQ<��}�׊D�< L^��{�A0����MM	&ŭb���[�1P��(�ٷީ���ڸ�O�Ţ
�R-�\�k\���ԝN��>���S�<R=a�>���A���4x[�.��Z�(iV�sm �ﲑ�Ԅ�a�Y�}1���s�x> F�*��� |�nP��ǹ_���:����� � ���\Y�y�S-p�sJR ���͐�5�w��FJa*ڈs�1l�g��ϸ����������h���Av(�� ������ (T�s"0流��G���m=�n��A3=��3!E����^eգr��9�/kVo_C��O�{�|s�j���M}�l�h�:�3#����/�)�<m���m`��L�^`���p�=2�Tb�|"	��=�^'��z��#�q���4PO���^{�؂���~h�Wߙ�XHKk�jՆ��ݣF��LN�����S�冝�1�E-BA��ꔫ�4%��A�if�Ii��I���B��̘1#��b ����G�v��@>_U�����[]{B�x�����>Y�>�<��7�I9�F1	GL�'�!&A�ˑ@0�2������l �FG�A)��Åtb�3[��5�$	�1�iv�{�:�|���L$�0��z�{ܟx�ĕ������R|�S�gr�����< 퀅`L0t�{�Q��Xo����C��<z	�@��u�6�S ��)�އz(lЁ���^@Ma�C�e��w�>���;E���.^�zU�����Q��K;m?NMM5��!&\�6i��u��ў�LW�RV�*e�.Ԝ
�$�P�` t/��2��#��b�9c@�c\���!��˸!_��(Rp=0�3���f�:��y�K�w#�����W_}��u��#�Lza٢���C�[���+�3�X����*j{�fO|�!m���Aa�f`e�H�d��Ը�>��;�4����5��E8������B���/|!���$�bya�@d��Z@�)_R��1�1ǙX�b5��<��]r�U��ͪJ��=X�=�1����ܟ� \��u�Pc����,���3��k��r�,>��y�G��	3�6�����0^�������� ,�8��(������\�������N1�0
�t�	0ia�0�ab9��w0�i���|Ǆg�>����y>���  @9 ���+���Q�T^�I��6��x �@tC»!����4�q�Y���[�C��p��O=�{�v�*}M�Ь�Ν�N<R���pe.ӦR�E����o_(��VON�A/���`��?��3/��<)g��7�9��c]5/��60Y�������1cl�27T=a��������{ǫ���l@���\sͅc
�3ϻt��/�\4�^9�R-)�ɫ�WSKKs �=�z��>������lM��lN�q>�7��(��Q� 1
- JO=arsY�Eh��T����[B�O������}3��,ۮ���T�8�+���o���M����i���R�@��Cج1�lM�w?�s0��A�ﵑ`���i �;� f��p^��ű������8��V�,�@76ʐ��bHc��Hߨhq��k]q���' $��K��γ�O�-z�'N��st�I�u���Ћ@��v�Oȋv�=��a��-�����29ai > ��_�@�0l�5,��q0��C���v���^r���0
��c�6Ң�Xo���z���s�"u��P{kNW]�>�=��z±�-�m��ڲ�{Z��YW&۬j� :l��K��.�{���M7�<��|�;�O<��`h���y��o�G���u�܏9�0n�/޸��r5�r<�x������"G�����n�馋��o��["�M֎ ��ٰzQ[����R���&���N����4Y�Oy���v=��s���,9�f}�a���Ą�pf��~����N�q,��p�
��<(?J}�y�k�UB�?�Ov,k�<x��y�Vؘ�e35U�6��?���ݮIo��Mݶ5���S�:�̋�ݕS�)�� ��i���*�bx1����
�X�Ǳ\�t�i��q
�9�Q^�H�2R8"�	�����@p&Ɵ~�)����7s�<��\ȡxU +z���5��	��q�y}���C(��`�.��;B��"��<���c��0�	`��:>G/��LpXυu����0fX/s���,��9j<��Ah�?!�{ˑ���� �乧�h�������Iͺ��s��YG����J����f�~q�㚶�Q�i��jd
�د����F������#dƸ^q���Qo�8�s�!��NcG� ���z��y�������8��$���{�a;�������Qq�8 ���~��7`LAxƅ�Mya�����'\)�B)���6���t��o�#�TO>�t��^f�h�]U��R� E�����s0��8��f�p.'fP�߼����x?����)[�8~�������Ї�SO�
�9�x}��sU(4�G�i�T)����0y��%������B�����p��V�����E0*�a�L���c�~�A�r�ӻ�Frg��c�n&LȀ��SB7ƞ� K�i�f�q̍�1	a,��3 {�9��yc ��|H� ����[�c��41���]E���B?�D�k�m������� x'c�w��ť��0n�H���n�ﳑz% vs��x>=��i�s�W��թ�m� �s��Je�~���u��Q�:Q��M:����y@�Y�������R�$��	��� )tQQ:� R�@B�Q�qG�QGfH�
�{g�5�;cEE�����S�~�o��9��rJN`֝�u���[���{?�����u����!G%�R��e���S��e�]�!8�b�40S�Pa���I�A��ڬ�3p}m����@�/�'�6�ߋ���q�8+�J9��>z�=�\7� <nժǫt,��nڬ�u-:����w�Y��z����ٙl�G͆��X�3o�#$�iӂ`~����b
6�Z�`��0ر�! ��1U𽽬�ۢ0p���U)���5���1=����k�F}�>�IS�虧������0�#*�L��-i��Q�'�[e�=�A���o@�
m0�s��km��@�s�n���¶����{2pa~ L�Ś�0��L �Qz}�*�E?-'�況P�3A�����Y�q�#��JPl��͎K<9ޡS.�ͽm��;~g��Y�@p/ƻ��k:r�c���B6��g�s�"��+���e ̭�������K�葇����ujn,k���u�Egk��պ��껏=���?X�}t��r�r� ?t	iJb�y�<�@_��W��6p�g١���?2¼ cb@���l����y7���#ք�X��i����X�ڛc�{�k9�N�:u���Y�|̠������?�е�X���">�g�q���6U?��h���P��0����a8��cDg�Y�`2��.x���E0<�C�0@�{X�:���zo��jG`��li���;tӍ�ʕ������go�[�v������U�U������9������Y7xt�A1��	���OWA��L�׈A86G����x�̭��`7Р�	�g�s,� 6MLV��@�Ƶ�m~q�P�ν���ڒ�	/�q&��;6�p?�1cԑ���dd3�ׄ����9���Q�C/�\�~9���v	 �N{��X��皱���s+C-�C��+��+_�??�U�^���h�7|Pg���ڸ~�n�y�~�����u��kn�aG�R�$�K-�F%�s�r����!?daYǋ-���6;X</��wh�<�gd�Yg�ٓE�9���>Y��+��3���g��= �i���	L8��<r��wlXA���u+LLW���� ��艺����Ц���7!D�d���6?X@�$ L��A�N��P�PW��>еM�	�c;jB���>X��dprj*��#�*��<h��C��RG��ϿI�-�������Kws��v�<�
��Qԝ���t��P%j{KY���0�OD&p���A�,�����bu���|��!е��&llN1��J��6�x������`WM
$9����`���C�T��Y��ǹ����E���W�C�`��_	g�K�����s�Ǝ�n�s�{���U��/�;���Ə?P��Z���jsg���Ň��(���15<���}�� �L/�>�&*k���b�.����p���P��oN��^`?��o`�&���D�Y.�[�VK�l��;��������l�w&:b�����sgiźez�O�14 t\�դ�	 �ax���N
�;2o̚=�	%���k�q���� fT�/���V��t��1gGV�a�WJ*tm֜[?�be��=�T}��3B&Вڃc� ��l����9"��3��cbS��3���O
��|��a`��8���06ؔW�X�1P6Ma�m��?@4`1��ǚi��_��@����w�cb��5�Ʀ����#��tQ��;��+�e�Wj��_W�k��[*�w���5�=*:���	����В%4�_k�}�W.�U��{�|�a��::��
���%�\4.�M�Ih�?��OA1`� D�s�	6\L���ڷA�"䎨�X3�0�e,d����R.���]w�qð��W�t��+��7Wߐs's�N;�T=���kɲ�!l��au�����@��`�ǃ@ '�pBx(؃Kj�4;c�Z=��c����q�Οv�i��.��%�os���-���ҟ�����cu�Q����|OIK_�Ѭs�VG���%�)͜y~a�\���µ c 4����w��?1Ǫ��A�ks/<Vsm�����LX���ju�{8���; �m��N�Ys/�^�G�5���s{�����ׂ�`�>>vG��ζ��8��h�zh��
ɦ�7�tipp74���Ӛ��z�wK��>G��q��ne�Ⱥ���T)�T*&Yq؄!bk^x�L!bD�xnجd�/�;�gy�[���0W��=�v�����0�
3' �{�89�lF���6�';1W��b6���Mw�����&L�ܸ�5��[�'c�舷�&�z������֮_�j�B�b	:wG��xP�^1G�[�����(���
��*��w�}a�
D���g�\/o�9"�x"�S%�/k:M���&˛5z�D���M������`�% L=a2��L��]�]���� �An�!FFqh�@��L��l��M��`�Vk�����^`��MO��$f�Cɥ�����5�m�����p?�9�K�J�ٶ]y���z�٧þp�Bݕ�s���Y�P���U�~��ܬ���^�ƾ.��\����A!�����&-��5���D��BRc��m�D�x<:[��v�����2�L ��	���1�W,���}cre�nظ��rJ��o�}��ӦM�8�P;b�K���g����<��t��g�W��^Z�2�1ǖ���A���#�!�=8Z�.���Y���r�uׅ����}�J��(�m���/�� ��@�-�m_�p�Gi��mzy���Ve2y54)0��Ͼ����_�ё؂�a�C'k���>fr��D� ������13u��P�C�p��X5�Y�ꟁq��
���MW����Ү��L*;bnٕm|-�m^�jY�Z*t��Tt�������fHDO�(��yO55�r�.)ϙ��A!���=}�����`�2����n"�K�1cF0;����{��̙�����:����;�@-��B�YͿy^r<� �p9��磏>����t���΄]E���9��դ5���4s����y=�̟Ö�v��c�p��!AN�Dh��@�`��}p���#,�3+S�Y�3��6�$��1 �U�]:SQ�5������6mH���*��qcv�K/��Z��v3��؄��>s�4�J�ⳳ�~zU��E���t�9��[˫?�i��sG 8�����֪ݖG-�0��YR�:_&�� �Kj��4�������l��*vwh���ҩN)UPW���B��1z�)gj̘�T�Шb1�J)q�Y�1�ݖ�3���μ�|@dy����GG�ܘC�B2'a�c5q �դ��O�+r>�&�{�������.��JB��j���w]���V�؄x�~:��)�(����R��x���6���z�bV���P�6G�9���{:Kܟc�<�b/?̖�!(�:�q��*�h�吨x2yңN��CJj9�wu�I�L�:�Ⱦk�a"��:w�y�<���A �)q�ݸw���1�:��H��;�m~qm�y��1���w��A#��Im;�N�u0������<�%��xQL���j,���ᯠ���W.��a�L�	���\���TW?N�BZ4I�'�|1qd��5&s��^s��z��fln�{�Ø�$1K� ���;���!a�1А�B}��_��0V1� -����&#'�6�J'�!j�̷�c�Ǐ<��u;����-���=E�6jB�	�a���o~��M��c@@x8� ?�,�4�,��:�<~#�{�w��� ���Q3D�I	�A��2��y��8�!���,:�&��B�[�<��
��rlwTج�&���kR���p5�J*���,��w��D���88� b��<f��q�c/���1�m/H�2P˯���}����<����As!��ׄ�ϵ��U�Ȅ������3=�yf�����`���x��C�U�$@K��|!�l�I�N��Ɔ&�����T	W��E�x,|mj8I֠��F�4,�^��l3Z���`8�v���a�0a��!m�9���F��m�Z8!�d��l.�J�\6��=��9���W���4�	7�7��Q�q��3��G+^Z�%/,U{{bǵJl�<�l5��WNm�{-�f5C����k�C���W_�C9��%��	� ݡ-�U���1�[l��Bq�~�����I��Sg��~C�ʩ�ҙ\���3�Sʒ*jea�I����L��sF$�jI��dj�X�g�v��;锖�\�i=���w�j��G+�KJS��U�u�m�}u�1o�GLS{GQ�JJ)�WJ��i��������R��K/�4�p�l�/�	��~!H�9��)���p�{�w(h���66�Ӭ�cC&t�����ߞ;w�u��c��qkV?4���V*�:d�)�������8I�M���Ͻ�ի��q �M ����0`�}̪��V�">���������b��
�*F!l4_��8;�͌�cε���*}:C���*�4zt�Ң�h�2���x���o�jU��� ���0�r��3�Wk��gD�!�W
�.Z�@ULu]~��q�)j�˨��H�Ѫ���^Q*3Fi�V��R%ӭ\:6�����Ct��E4�B�3gN��w�D�>�8߉~ ��sX  c�.�1_��`Ä��DJ���t��Cr�Y2f�6>B    IDAT&��];Y���R��调�����	Kt;k���!��}g���l�֭��}6^Yl�WV= ����P������v�|�PҎ)�1o޼p�PGTH{��߮�|�3!J"V�$f�-Ղ���L���l�F�ɨ��U��l&=��պ䒏�u;4�
��JF�g��)��1W�R�`����pL��k�H`WH����5�������h�u=�3�ÚuJA�,�њ�Z��G�R�Z�^�|-2�����K�Z�,;����>��`������ʃ=���������!`�kӣ͛�/����Ô�(�
^8�ӱ���W 8x��_�"�@�l`�Zeg�]»mX�P�uô�� 8i��V�iJ�I���ScƌN2�÷s���8�֋3&U{,3�_�g�(�DG �ޙ��B��te�`����C�j����L�ݖ7nX�_��:���:��7)�Mj��y�K���Zs��E�% ��1�P�	�����
d��&�W
����}�+�fRjn,覛/���:Y�9�TI뷿y^�<�J|�&N<P�JS�쳱�.D�
�`I�� # �@|�C�8̊��d�'����)TX�.	 g�9��q��sc �?������kሃ0�&*�Q�;�7�R�T`Ι3��ag�ׯ[Tױ��Α��-�C=�jW(�<��#t�'�% H�H-�l���#�P�����s�y�sQ#0�� ���:��x�� a��Pq@s�6��� �J��u�LݫB��>K�&�Ջ���}g~@�B�*���� 3f^��p�3�g�`^�WmF��hD;(�W
�+V,�c�������-��NU:UԿ������Y�^���O��1ǿ9�
W*�����F�f��0�ǹ;b��Թs熞�9����.�x����M� �DcqVᓊ��#ށ����)�@���E��.�qkW/_-�@�#BԚ٪VTH��DB�:��nq��,�S�(BA�t���PT��8�թ�t��2樂d�`�5]@���  �`&�ӏ���s6��hR�ahwΟ�g���&�у��}��[�?�R]xUH֠�O(����3߯)S�Y�M��F@xg����m$�J@���M�ڵ�ScG�t���k��wjs�z͞s�~�K�P��n��Nt�a�(�\}���d��#�a�c��Z�X���wp�S$����q�|r�q0���D(>;m[1����ua��;�Zda��*�e��4�8[N�ӏ͝;��ag�J�
�`��$麥LA��u���ӓlX�-gX�xKE`�-� /�W�w ��~��E�Q�ױz@�v�@¶'ՕԸ�w�������	g��ޭٷܨ^���������c�ЦMy����U.7�,*>�͜y��L9<DRT*���8i��H��p�@��RwG^������Ӧi�����Mw�W��V��s���a�&M>\)j:gɈM���٤�3�"E�Al64��.�|��7�u���8��q�`��7{�p�5Ny�k<�b�`Q����WųV�Ȱt:��.��7�[�n�xbsKc`��1WW�Ls�8��)D@.�B����u��Q�K:㒌��p�w�:�Շ��pC�\[4Ǻ+��&��j�^&�V9ߣٷ^��a��^���M:�Ѓ�l��:��K��7&�,��`��9+1G���4��3S��.x� ����z���RW;󮬹�]��3OQ�{���>}sѯ��}&��+����NRO1��!	_���͈�\a�q���\O��;v��������l��̆�̵��qDD���Ys<��,�h�kJD �zX�����V.j)t��ڹ���	��	������$����N���d������w�WBg��0O�	���3��.�|����k5��k��tj�y�ꃗ����F=��5��k��ѨR�Q)�Bh͌Y�4y2;�ĖOU4�W�17��C�8֫���7*����.��9fq�
�0��5TD�p��p�^�&Z��uX��q�'Em��c�]��>�~��,�=m����N����R�O���~���};�;`�y���qV����{�BZ�u[MB�w��0��'�Sr�!r��Mrh�N[7PL8�6����΂0��d�Z�`�J��ru]�u��������e=����_��^x�U�l��v���^�^9�;���/�����1i��L-���1N5�|l�O�����׋�.Z�ݖ������]�vQK���0��qN����������5�<p��W2l>0aq�m�����3��!��I����qi��vh��]�������Q�JS(>M�f̚��p�'��T+u���A�=q��n�\�Zu)��S��"��p��<�'iF�G�h�������l�LV�8�k�-�1=��Xc��xΈ��#���/0n?�f�p�'�.��@j������g��}�N���~�M�+m����<�6�ݬ*ŋ���ŋB�:�+Axي%!v�T(i�>y�L�q扪���֤��m֓O���_����J�:��C!����I����W��W��ߛT��oG@ئQ����\y��NL,�g��wo���+�u����X��'Z �>�@q�H��^f�NQ68 L��	q��y˽0it����=V�2��mVS�h-{�]g�y���f�������A��)+�)�*L���꓋ۛ�=F�q��/���;9�s=x���:��LĬ$vV8����w��^f���t𻁆�9�����r?��+m�6��?�q^L�P�=Z�4�\����̺�6G���g�jp��o�1�������Ƞͽ}_��>�{�c݋���0ǹ��e����scW��eID���.�4K��r�f��N54�U*d��쮍Kjo/�P��u!A#��͙�b���W��7_���gm<������ZY� cW̼��S�����+�9�U��|�Ec��'_��v_�jѨB�I1a�[8�zŝ��TK���|_���\fC��9�7��p|ߪz��vi�j�H�bSV�j^�BU+���K�/����*U3J��	�8W���5�����d��3�����d�i��'�A����,��!+&���kX����f��z�5�̽�Um���l��p��f}6�����m4�Ƌ���'&��^n69X}�/N����	䁺o3��������`��˱6�Y�f��a�bD�bY[�q����V�I�A�>�Mܖ�����#���bL�Au�4~L�.��]z�U�E�D�R��S}ݨ��y}]������f�&c�d,Jxq��3��qw�ׂv-��u��{o[�?��+vc�Hᜪ�	ׂp̸̰�[���9H�����ʃ�5h��vA ٢�c�~���Ժ5k(�r��r�z�*�S�ohQ)UV*]PEe�
�#�-���(��ʹ�K�<�'񍞔V�a� �����4�&����ӓ�L$��a�-j5׌ˏ��!k�~�y��<d0λ7��b�N�`�um�6�Ӷt����ك\�u���݋�˪���=��1+�6��5G�HUl��d��W;��3}����!O|�u1]��y�~�����k^di�Uk�(l��UL~�?��GWV-�hۨt�]�P;K�6n���{�Oz�v�c/e�.�N��t�Du�)�6���M��˹�������cR�������~@��y�Wu�Q/�H[���c�K[
�0�~A�6�n,>��b���U�xL��~haN�r����sO������IM���F�lV�RU��8�U@�"M����[� ��;k��h3��K�l��$�0Q)��>1	*�!A�	j(a7Ȉ8I�'��_(t�9 $��Z�����'� �qA���d�=U�l��b�]p�N��dbq0x�:��ɉ�Ǝ?ˀ�L~��K6��L{�;X�Z��j=�|Iq �+�^C��I�B;�XDlF�:�[& Km�h�F�i��XB&�.���m�t��yCO��g �\YA&X$y�ĭ"/�̟Y6ϖg��[�ߕ LQ��}�U�lST%^2!r�v��봹�K�:Y�l�r�d�qU*�{���	O��Z��s�x����rCͧ�߇2G��%[1h���]½���΂��
k üϷ����b��̭?&�C%�7[/�淿P��LU�Rw�l�ʤ���5&@�) <�d��a&7���%�� �~3��8��p���0)@��JR 79�8a|��\yw�1�9 ��K� �g�@1񩻊�)�xҖ_���xF�-���m���B �v�`��I��Oo[*Ϙ
ZLt�B�8��}�%�˽�~�\3��~�0� ����CF�G[��"O�I�*�����!��ܗPo��bĽ� M���:,X,T���; ̋E���vȀ?τk"K@��Bv$, /G}�4�+Ax��������J^jl�W�ܦ��M�$ �󅂪鴎<��e��ZM�.���WM5�.y�8d\ׂ�@�n{�����������= <��ˇ�9�Q�)&<��QadC��b����1� �؛��\�kS�j��?�C֭U�ܥ|E�[�M�ղe��kV����J �`���c�2Ø(v%� l�	 ;X�?�,3�aF|���9�&�yp<���
�	l  P� HS^�: nP@���H6��`��I�
�'���Yک���Ϲ ��u�v��~��<ٶy �̖{q-&�h3��Q�q�S�C�],, ��� <��*,<��s/��>Բ939�Ŏ�xN�'σg�,���^ 8l�c i�N_YHXmd�,���`[6�;���b��<{�gjA��^�M����c�}G�.JS�5����&�^T�浹s��~��z�[߭}�>T��U��3���9v�B��l���V���s{M��.B55��Z3���]f&Nx��+5�;O��φd�TgC&$k�����r���<B1(���*n��U:۴�X�G��"����L$۸��Ô��;?<��L�#�>w�)�U���ՓߨƦ������*��Z������Y��z0G�5�bM:�e2d�kA��2�`c�!�~� �l�]�:1��<��L~ؔ��Ӏ�1��<X[G��#�r<�@�8����y����� X�B#{���\� �xN��H�7���q.ㄾ��{����?m`���������S�9`gq��� +�8�|0K(�A.Ț�T�b���A���� �bd�����>g���g��u�xq��;��MH ?�ݶS�a!`Npm�X�I�,c��{7�\�bqp�mZߪ�v��}�l���ǩ���r�G�ι1ڼ9�je���VWwYM�Yu�t�:�����Q���Qf�|�]܋��X,s�`<ύC�)��e����������No�����4�|Otļy����/���ܴza}��̦Hs}5����P���Jp��q��OT�J��{6�L
ob���*��t�Վ������d@�v����������	�Þs�r�z��Z��S]t������^
;̚	���Fv�M� l0 &�6��H>��C��N�(X-�������W�@� ��f���0���G����C��^`ŨͰQ��8R���X8�@���� �˱�����xؓ�aV�7�����X!;=c �9�1ǀ H�1o�BΜ���&���ڮ%���{ ��XlXt�&�&�"�<Y� T�@�]a�L��&���dK�i}@saQ�"_�c¶g�"���ۆx��$ WՒ�/�-Rg[�Ǝ�j�͗�BX�t�ڻ�4n���v�mzmr��Z���U�b�++��w[6C��k��2 �w �,���f���LМ�#憝��a�&*�D�d��D���`G��J%��'|հ�0{��~���ζ��)�TQ��O1�W]CN�<�+%*��� ��#<Ջ��g�B7�5x۩��v�#`;U�jq��"�@�d��!?y�3n�~���j��M�[�:M'��`Vk�t�S�	��JՆ�w���5�� L�"|wu5;��	�2�=� A����dE^  �= fnL| &� 7&7�s`��x��+0cB0�`�� ���po�wHh�L��6/ �q�[�\a�,V�9���l_f�� Ф/����-Σ=��x�^��π0� g�q]Tz��
� ʹ�``�˸����3y.��p��EF�l����2d� [�s.L��3��3�9�;r䙳��o��bf*}�0h�:Ni��%z��_S�R���Ҝ9�駟�;�T����	=��K:d�������Ss�u�t(WGQ�d�O����5s5˷&l<�fc6���M��/�\kb��	��$yZ�&��e�}�	1G��r%��~��{����-�w_�baK���lu"@�R)+�n���'L�-�؀R�H�B�L�o��V{��v��F�� �J8�Sb�39 ہc/*�������)�Թy�����6o^���G���7d��S����_����JҖq(�% <� er�����Ң � Z��3Fd�V@��
�,lK�X�C^PX2e�H��°sO3E �g �ƦG� 610�l�@��!6Q �k���}��2 3�M�8�>9��`˽�D�%@� sM��Eơh��1���P��	�v���B;+���`��]@��J�3����"�2�9y�Ŏ6�Ok�Ȝ��\�5�d��	�̐?��5h� ���y^���?�+�l�KAx�KZ��UK�Jk��Ϳ\�{�z���ӟ�J�7��|OVW^s��8�DeӣT�H�2�T({03���GN��y�hO�ƳD�@V��ĵh<_�<�d��r��q<���D�geG'��:���W*�
Lx�A���n8d��Uǔ�Ǳ�Z!_
�,)��^h|��@M�vb�`GC�\<�a	�AD�a��n�4�z�:������78T�������N;P���f�m<n��ݺ������뀃���7�z���/�×~Lmm�p�Rզ^&|^ �lu
�}v~��&��ʢ�בpV�@�LP~�%�¶+d�JS�=�vu_�l��0��'��sڬ�c��)���ن�p��{  fl<&�:�~�xb0������ar�x�~ Q�f��G����1�Vo���N{i��/:|v�/�O{��H�s�#m������<g��$�����lwx�e�}�䲘�f�5�v����ыK�롅U,nV}]�����f�|�6ml�=wߧ�}�7�m�7�7ݮI�O�]=��R��d�Ą�{ĝv�i����(������a�4.>Ƹ����7� [s�Y�vf�c�@:x�g��&�q�K���{A��ٳgo)K@xb뺅�]m�3�\�	
y������+�q�����eU�����gM�`m04'��@C�`��j�đ�n���\F����g6��Y�A���C~%�|gE�n�E�?�+e�6����[O~��-[����a�{T��$LX͚u�&M:X�\W������=�j7�b�۔c�*�M0�����;	��������68��N�>������v73�Ë���+,3:O�x�q�l~�M��VK�����;'��teU���Y�q�9����30����m��2��W����Am �Z �Uf'����8b����8(�}6�N��6~w�`����#vx�c�˖�������o��	ҭ����N;I�m��9����T��{����M=�(�yerITQ�i�*j�02@���;�`*��8ϕ�Ȍ� ���������52��*�k��XC�q��@��,�D�`�w�5��s��t��a�Y㈫n:t�+d�[��A�!�uww��o�K���m����i���a(m�ST�Xږ��6ͣcѓ� � �O�l��7T9>�+_	v�3�8#�!��F������ǜ��+OG�    IDAT�+ ��ڭO}j���ԏ4i�x��wh����3O��%L���T�և*j��9��!�vN��.6G�m��N�X��@��6{d��r��"��;�œ��s�rA~�4l����s�����3�y&#���ʽ ,��g���|���Ά3�X��Ȃ����U_&�ߛM�U#{�9�?�JdO>�iƖ��N!�B�9����=�!��Ym�4r��zA�>������{YC�Y���SZ�b���Ejoۨ��Nͻ�]p�iڴa�>�/�_�ן�Ҳ����'t�qǆ"�
�d[#�Q�p�9��o���l�v�7�g��}.�5o��0v�����O�<L, ෾����*X���8��X���q�E8"�x���[���r&�}��9w��i�h�G�Z�`�JǱ�g�������t��S��w���Z&(����O���)�L�1���c�;�ٝY	��mo{[��~�{�9`G������������I�A�9��=�R��n�2�c��X�]v�>r�tuw�h��]p�uj�{[M�#f]lI$v�����Q�X�/��<t����'��fu� n���,/��|�sl*�y�A��s4��e�@����ф.d��	�1b0�������@;=�j�7�r���%���k�6��k��rl�����w�s����}N��5,��vm�#�ux�ŋ[��A:�%K^5���E�4�u�-�j�̓�M���_?�O��`�,��Oܦ�'��ik:$h�v�9���S5��1g:V�BB>>�<�����*����
��9�6f������9�@�߇gRL�e��t��;�뺩S�&����4m�L���������:{��Gu��}�;C��~��:;��
�xŬ�3 pf��`KF��>�h`��G��X_�@�%�53 �=�s-<�cV���chS�"���z�ձZ�<�kM:dM:l/��}�z������nVkkZ�*{�I���2:k�E�t(E�]E�]�� ���<�v>���F$�J ᪖�X����ʥ�V���C:�ijl��:�z��.=�41�j�}Qk[���L����جb>1���	���}����H,,���4l�̗���}�-� #�r���hD��W���	<6=،�Eڡh^^4@�4m|S�F'�(���J�J�\��;����
�؄'��]P��z<!j�i�6��N�!S������/�PHV�����%�ۅp<������?6�X��a' �����9�;Ǹ���5����إ����R�s����ܨr�S�GM�_�ިY��PwWV�j�7��f��v|��Z�gϬ��tF����.k��%z��QCz�T�М����oR]}^�tFݝK��W:�"�T�dT�P��v�b���0G`jt$��ؽ���`���7�	0��a��=*�^1{bv�s�5�X��и!�6E�u6h����������RK�l�����#�<rݎ�A�0 <�u͂����c��e�5�y�>��KTɕ�_��Ouw�H<��Vt�^fb���x1n�i�Y��P� gױ���TΪ��w�3���� #�4�#x��n˱3����nuu�V�ؖ�vR$k�U*JK�n�}�}]�6��	�>��532G`~�-�/T�1�����#Ǿ�0���/z����zM��%}����䓧�P���J���,��'�\Ɇ��L�M<��3qj�",�M{�ñ_�)�NҲ�Λ'{/��$�g��@�W��::�� q�|��l�	�����a&���OÄB���e�5o�m�s�1�w�Y	�c7�Z0��}<�ly����^�v�~�įU�%�/Q�a�?²��6A��*d����'}�8<�
v�����á�V'�Թ'������ Y�X��?�ca`Q�uVUPO~�~��k�3�UW�S6�l�Ġ��(�kR�C��I�U6�c;�R|;"x��@����;z��G$�+%`^��y-\�U�Mj۸I���'�|s���+956NдN�!�r%qВ�L)K�r�]3��π���K�%`i���Q4` ����7���XjL�\I�s�CS�l�4��\���8�,<�`|�;�	�'LX�\.�y�n�İ���+>y0��K=�I�8���u�Y�ӟ�{R/,Y6��� &:���!^]Tg� l������P; n:H��?:(������Fx\�$�jbo:�?Ɋ�.E=���*tC��J�;ܷГR:ۨR9�ԎH'�`�	;:"��� �����n���~WN��k�H`g$`~a�sZ�`�*��+$tmV�ԡ�F���PS���>5z|ؓ�2���$�48�z��8��sDQNl� N0�a�~�l'�v����û����\Nہ�>9d]:���o;|a���G`
\��.��A�j�C1��,�3��O+��<q͚���]Ӽ���'�E�z�;�ğ���V�8�L&�c_1�I�\���Kh���C�G��hv�qM �&ah�텈�`�#r�8�/��}�����"�=��p�t��?<�[{���,;T�kP�T�L�)ls��IBj�c.DG$�<Tt�P ;�<��ᶹbg&��9#ؕ�cn��e��N�K!���fحF��:��6�\M눩�(Wר�d߽�IB�P�$��[��Q�t�s��/��hѢ>��a^ޘ��8j₩�G@ؾ!;� r�����7�����IGP ��_Z�d���L�sn���7��M�g�w_�vas�sZ�H��ģ������Ǆ�e��T�0������E1�F�����>��!��f� 0�������#؏|�#�1�;�aV؎�f�i�P����@I�mՏ�oZ�f���;d����Z�d�2��O�	' |a(�CQ� �C8�2+�*�@LyWN��k�H`g$�5s˖�ᇿ�R�K�[�j｛�Ғ�w�[}C�
���<��������8V�=��	�h0G�Qi���cg��~O?��!��㏇�(�*k��8�YH�@(,�3;���9��	>0aGރ)�3�=��Ď�a�|���V������d�}���e�TQ������@xʁ�4s�=��Y=���}U�h(6a�ZbػR����Xe �L���0v!�;��L'�w5�Ky�)���i�Ɲ�e��1ʓ�̹q^TF+�6J�e2��K�K�����/��;�����*��E l��+��#������s^	��a�=�P��.ۭ+������ְMXH��ꐪSO���:5տN��(�kf�C�H�Z�`A o���>")�=d�X�D�M�x���;kҀ-�	�&�i!��%��q��tl
�0�����,�=��#jk߬2���.e�2߸��oVs�ԫ�?p��u���'x�Ͻ�碑.�0����~a.W�b���@��b�;��-dG*+a��=�	�� m�cUB(mm����Җ����%Y#횟}�R��Tvj���l�ޣT�Ki5���/��z��X	�V�	�9����\�{ߎ*j��)�0{�"�O��":��<�F��T�N��~5���=HF��e��B�j�G�M%͛w��>�uv�������+sZ��S��8U+cC��T��7"D-��>�����8I r�c@�;8�����N�ҹ�dġ����8���^1���3|��`@�&� �h.H!ף�z��.es�o�y���k� <f��Ec+�����!jg�}��;d=��ߪ��6��� �� �8V�^J��� ���@h�|�^P�9���w1j���"D����W��+ck\"*�#%,8�8��ؼR?����v�[�v�F�\�Z��[g��A�J�U�6&)�J' <�PeȘ�Q<c�ڀ�� a�;j}pL$���!x�}��#�-%08�Z�R_���*�ݡ���n�w�Σ�p����v���詧�뭚0� 廉��R�+��$Yc06�?~b��� + 's�'~v~,͊���7�9E�0����s�{z�?��ݗ�����	�v&&��`�����^?Tf
)'Y�;�nXA��5ƾ��|�	��LȘS?J�s���������z���a��}U�輙pl�v�\S����&8�!ܦ
۔O�&LX�� ��[�� �̜��Y`�0a�6�A8ؑTR.]��]�������f�#��
B�ٕ��>���T������i��I��5U	�4ү�����������Z�r�82A��#�	����/_JY�-Me͞�A͘�%�����|�a�ZӮ�o�SG���aB6��	c���K5 ���NlvJ��|���aV�h1?��o��0h�o��D��p{G��d�E�l�4a�9�{`��
6d�h�إ�z7	S;"��}���f_7u�Ø���ؽ}ݢ��'����F��رct�ߢ7|`��t���t�@���<w~c#ƏB� 1�%��x �f��}�C
�
��������?ݷ����4�v5���	��@�;���Oݡ�����ܻY_��{t��x�K������NtD�T��a��?t�z�����g�_Џ8�/�3���\t����xG bk�D�����t���K`0���׷���ݝ�R�-�߯3��6m�ܡy�>����/=������:h��*�K�P�.K텭���˂��5�*D�9~�m�з��H��Ox|�B�E�a�(�f��2�_�yET�\����a�r-k�f�0i���&RI�F�%[�Z���G��'��Z���~"L�8a�@���|ԡ:���	��+^�[��h��i>�����go�� 0�r��O�� $�>���"?8�"%� *@��j+�ج�.��,�RU��K��t��y�w;>�z೚z����3.V��S�ڒ�p�N3g\��SV6[��U*8�f��a(���vad�`r�~ ��ih���^Ԯt�.y�����70���Փ� ��Y}��o���U�ZJ�u�t�9����_�u�ݮ_����������?�9T�G���Nl�ٴ�����'l
��
iD*�O�_��onn�-���hB\a��m�Acv��_�4�'��wQ3��b��&,�u*~���e�ד�J]]��[o���iӦ��؄ǯ]M�Ɖ�	��a{�t�t����أ�Ӹq���p1�����?��`�&�a�AG1�s\�+k�1���3�LJYb��f�\�LV�/|�AE@�<Xo�Dz����(��on��j-_�gM�����7j���ֺu�:����z�e5�4��A�����c�)2��ׁ�6��4��]/���D_-�Woҍ�iD���F��|H����TԜy��Y�RG�f}�s���=�55�^�Ι�>$T#ĻB6]xU��}:0�ڍ>�1G=a���-���s�����:��#+�〯Am����C� ��]��%P���� s#đ�9�V>;�ӛ�Q����% <a��cʅ��ޜi�mη�yT��2U�7-��l����S8� V^�upN��f����F$k���7�G��T�{�VI��io�{1�ݖ�b�v�؄�֍��ݬ�z�N��מ��ԟV��SG{��j
�`�9+؄��\�u��N\�W�-R���"��1¶;8ݵ/���`y�H൓�� �l��zh�u�5fTJ��z�f�z�*�.��W�>���I���[u蔣�1M�1��d�^��0�
3�ܹsÜ_�j̀��������ĵ��i �d�;��8잏 ,ٿ /�؜	���L�0�g��qŕJ��9��[o�5Lx\�xb��
�d�D6�mN����1�����B�Pv�(�����xl2 0���#��@�]�B�	cv�m�qp��5�KF�6y`G��υ]<�쬑�1ݐ���_�{B���^G���:��m���s����؄{�VΜqn��H2�
�i+(��A�v�N�	�xG�D���+C���L#!j�4�Ϲ�PL�9-x�A廪7:�o�0�ՒVO��5�
��/��>��Ɩ�JSE��v��U%D-�Y�?f���p;s�p��͋`�
���?>�)��El� 7$�k��t��ǥ-}�XomD�wo���@8��>:w�܏�n�DG�ߴrQK��D�c�ʬZU�2�$[;1����!旕��sgX� \o(	Sv�84�������5RFWWO��^�u�{OOWXA�	'L;a���`�`�-w������Ru���K*�Z��6�;�*��4�PN+���sfhʔI��Q/�=�Q3�H��i*�8|��r/X�����Ȏ�F$��I�NHQY�V.	i�]my�4�u��W��oW:���fG������)��Q���Ja�V�$`�4����,X�Y�%m��k� 1��j���|M��/�7��p��zY�\�;��r��^����o��U�J���I5�;3�8�
��&Pώ����;4������ $�"na�ɞR�0��1���q�^޸B�\Y��V��W�I7h��n�}���^U�RU*KX]Uӧ�*���M���ԃ9���AB�9*����x�����H�l@y�5"��N�0�d����E��OiTSV^��t�a>aehl���T��Ln�R8�S9)ݓ��R��L�1�_ޜ��Wct��I�5�8�y�\�ak�6#�D%�b�͈��7YuXm|_��X�N�ӏ�~���+u����n�b�b�DG�Np��4�g�!W;��ǳw��ةeAqm����������?8��%������P��nP6EUa���F�Z�I�FOT�RV:���Q��;+=a4�8�@v�X�Y<�5�xa�ܯ�$���l	©���X�7*t��l����UU�Š92�w��u:餷j�}V�X�bU�$Ta�`g
"����-�y�0�dk4c��9�j��kƱ�����9��սE�|m�g۲ύ�V|=��L&��m��v�����k�*t�4Ä�ej�T�& 3e�h��r�7�c���ʎ-��8��1��Ât57/tX5SE)�YO?���=�P/���5�K���ZT�H%��Iv��sH[������PL�jmÎD��O~�`Ba��S�Qر�&(����#�m%08��li0!T�%5d�JU;���3� �f�l�0f�z�0�5�Tr|p�=sɅ����1�=c�͵ф�1H:2��ʿ�e��1q���s����L� �N��3����9�U;��M��|�'��}ͪE��0�#P'�
īIl����U��lA��@��<�=okU���!j0�r�]O=��
I��}�
9�ꛓ�wҝsd��8�����O+`LD^Yd��h�XW��f�#{��	��%˗�z�*���*aa�ʅ��Ad)�ޤ�R��@Ө�*���5%��{#h�	Ywwg�Y���f��&s	~$,�6_�q̌�ƌ>���p�&E�|��Zm>&�����;���W�)e���#���|��ի���X�A��qm���Z�N�	�(f۱m(�	W��ݪ����ڸ~�����rwO��+��P+�Q�J:ط���szm��Ʉ=` c��������Ӊ�F�v�,|�q�#��cF$0��&���p�C*vQĦS{���1Y�H��ԩ���1����G�=��W)5(��뫔X,���r98֞|2�Z�����kf��h3&i��c�5�Dc�#f��c��{̒{1m׀�k^Z�R�~�@�T5٢�/��f��+�k�c���%bVBǂ:���!(�f%�  �X�O�sN^]k5z�¾X��Ű��ŭ�m�_��U*��Jg�# <eʔ�6G�]��� Y���:f��w��,RC�p��	��e+_�׿�����7�NW^u����#�V�
Ŋƍ~��;	MjT*�$=�h<��|Ü�gBW�]'�I6>�1��6�������c��ٳA:h���0������y,���k�����Ͽ�Ug������W%pcP�����m�v� QO��X�<<v�&��M�`�<,?�-���J�.���~�(�_�\}�TNk�:w���`a    IDAT���G9�2I���ӧ' �#�����h?�7+��u
pf�%�G��q��w�z��N��A1�/�õ���0|W��Y���>�L�G.��ٙ�vN<v�����/y>���hVIs�\���y�r����FUK{hs[F�7�U(eB\=	��Y���5�xLHb�y%s=a�ۚ	�x{�qb�'� x��s�W~����&ĸ-q|�.aGG�*u��=氉'�l��|H�pt�qg��@v��$aN�p�Z�[���yW��5�2r��q�M%~o
Z˄����Ӫ���{�{���õ�����K+W�5}���jR��S�.'v9�ܙ�2irȶÑ��+MR��zW�����'C���svtt|�dlj��JaG��?�M�TiKIQ����n��ğ����{K_�)���[]��?�;�lyv5��kp�s�U�\|��������;�l���=nG�G������#�RW�f�]��[ޯ���%$cY����?��C&����N��:KeRɶ����Y��ɞn�i�1	ۙ>n��\�w��-��o�I���N�5�����keҙ�ϟ��2���5��d@�=�`K������x��44�w�"���3�p�2 �ٕ��X[��9�v����Z��Ԝ��iݚ?�sO�͟�Z��f=��Z�:�*ut7��\�t]6DI�7s��2E�
ay V@���ϔ���U]�>������|�eb�-R�L�d"ZM��[/r�N�-������F�����{0X��D�Ɇ��ҽ�1����}�xy ���緅�mӇ�a��`�����k8�$)+��|�2-Z�/��lӨ��n���{ީ*���G?����s��P�k>z��:�x��;�9�TnT]&�j%?(�������w��П�o;�I}���n���`���~o�mw_q�qSV�H�����τuk����0�R3a2� u$K$5|c;�iz���I��c�k�٫�s��wtv�Z�+N{�D�퍼l�
f��ک��\0Zw�y��9�h�^եw�~�z�-*T����<g��v�R�l0q*3�{Ad��3�-�[*��>��I�c hIo���m�3h��kGA�(�[��=F�w�~}�m �5���c���0�$S���{�!A8�pU����\m_���f�ܺ7����P18W�t�-\𠺻6ktKU���A���ܺQso����ȟ���[���iǩ��M�l&T%�M��Lp1�ZSA-�>>�d�� k?��$�^`̾��� ��cRi|�%�߻�ۮ�8a����q��Z&ӥ�M���۲WS|;�\/� ;�l��m=��' ^��p͆m��M���%��i�l,�t�N]m=����5a����懪m+W���PGw���z���^s��:[GN=J�䒌�
��w\��cOa�d�0ch���v�z:���Y�1���b��$}
��m���jp3��(ÔR���H���X�v���X�I�h�����HQ��=~{�E��ķ9H�v�r[�U���}���ѮQ�Ӻ��K5}��նi����&�ት:���u�e��ɓ�ΕU���r��j�8$��i7C���\r���;I��w�U����\�w̘Ì�EcsD6���=��s�a�6|�,�ݖc&L5@���\R��*���!�������pd�'*���+5x#(µ;#���|;WܞT�*�L����-�d˪��K�W����?Ձ�ї������?-�E�Fm�)U(:Bzr:2َ9�U��]ׅ��v�����`��̒Wt�P෽ ����''��&�W�����@̴������>��)���`~��]�Y�4i(�p,���� ��m�  �~�˖/��C]��4�Y�e�e:������������i��u�'g��#�R���i�V.���	T�2�؜8T;�s�:�#��c�F���Y&�h؄�Q�����xf0�S�{�����{�U�
�G^v�!�Z�,h��<��-a�N@8�K���[���!����aa�����l��ST&5�N� \���h�|^�öG�ap�a@!�`:�'e�舸T�A����wv���/WJ���+>r��Œ�����>���*����@u��}g���=^�<!4�`��5�9b�I�kn�[�q�$v�����@oi�P l�ؾ�a��Sj`�P�P���^����P6��Ȯ���؄��M@�H���՟\SJ)b�۽0DK�6�C�;��[����2GP[�[�\���657V4�+u�'+��~��g�������h��>v����T��Ov�	�l���0�0°�F��1�M�i͵�(f�: ��h�^��:��E0������7��7�����n�͙3��a-�~�U7�ۆ�{:�c��؄�J��l]F�[���Ïu:YU�0�Pi�0'������c����fwꩧ�z���8���/��{�e9��.�f�\��A�+�VL8SV�g��x�'�<y/u�!��˨�/k�ڂ���~�wfƣ�-�}�{���p�J=IȌm�M�!A2������w[�l���@x�I8�c���?`�j���qt�6����Ȃ��0���j�^-�m�{�/�dk��|3��(��o���n3~mӏ�@���y$�m�0����� z"��3�&�
;T,x��*���PԜ�.׌�*�+�����K��ǧ�h�����_�C4ԏR�@�U.�Sjm�1�����k�;���di�=䍲d����k��%a��l6���v�'�x��8�����${�Q�2�I?v�]s��퍦^��I�oZ�  �� �M� �����~�Lc�� �m*�6��@t��T�uvc����1w������c�=v��&�	so�f΀�%�\���U��Ù)J�M��{�Ǝ͉ݗq�Z�g�yI]x�:�R��T(R�>]o<����	�
��bZ}D��c��VL�wB�fǓ�f�m0�G0���1(hl��k~(��\�õj�G& 80VE��D�b�ۧ1���� ��18ԫv1��0��b^�z���_��ݪ�/��[.�y��b�S�,��ܢ��Ps�x
�r5��b��+µD��?�]�&��5YФ!��*8�\v҆�T�F4z��9��=�zꩾ�,��e���]
»mZ��9�y,NK�I�����3�l���z��a�"i���A�1x�#V����g��q�V/6�H���/���?�τ{�U	[ }�_[� ��N�@��1{7ͬ�w�*�jk_�Ɔ�TI
MW+9��x���o�ӓUUuJg�rw�6Y�nPkx�I�ϖW����n�֞X��)_
�℥;3)`xXM��JbL�H> �x�����g��6Ɩ��P&�>U�8��!V�X�ֲ��VD�1�}��'�%���,�Ύп��+~Nm�ĹB�կ
a�������F�]ñuu9
� �*�ej�x"��{�����I)��λ%� �O� �-�^��ܷ��\��I,ט�$~�$���t~0p��P��$���(̍�8���uu���~��}�qe�%K�����:���IS�0����j�(j���C�\����L�m�R*�jjjs��ȩ2N����\gW�g���ȁ0S�����TfK���Ȅ���P��Nv����ga'��  �`	c��M��p.�I��aA�e���q�]�L�:u�v[>��O��v̓�
��2�Q�(�?z�({�њv��Z�z�V�\h���=z�Z�^i���st�ݖ]�΃��`�l�	�bOfu��y��a~FV��7�����s�;6wl�eu���O��Z�v�Te�����ƌ�C�ֵ�R�*+5�Q=��{ϰ��{���ޤ���'O�؞h[ؾ��l)~@mY�aI:vb�J��!^�.I��e�"���8&nG�����&��+�)t�A�� �j�'wr�d`�a=\{7:L�c;�(��bU
q���`�b��$B���6�j�� Ό3#c��MS��'��"c�&�<b�N�p뢄����2�<qó`!������_�O|��8����6?,5f�-q���/*p/z�L�Ֆ
_�s��U��������=�+��6��o?�Xجa�(�D�ӄ��e���w��ή���Mx�Nz��zݞ�W&S�8��qT,�o	�����K�ro^0Q�a����wt����;� ��Ny�P"ֹ	���Ш�M ��/��!��x1��&X��6��'�%!ʢ��� ¹�G���k��'�]�`K�+0a�C���#���w���`����/���\~X `��:�4���J������}��U��a2�m��0-Pi��b���_���m��<�`Vm �-�R*t�d��*;C y]]�@����=U��/{�'gUvf�i[S6��:1�CH!�PU:�ˇ�AA �PE�E��B	5�Jo"Z�	���u�;��y�ݛ1����_���o7�3o����<�Γ\�e�!1	����Xc���J\�?���V��/�9�M�;G߳EwY)̼6�n�1�YW��ݯ�Ɯ'����8Oĉx�|l���1�
�LB��.��m
����A�o9��Ka�M-�7ӓ�GI�1aס���\���}�SW`��-"��.ס�Y]�J�	Yݫ|\��/.\ǒ�e�� $�]�u%qL�����qt��Ɉ;6@Ι����(�����g���Y�q���f�v������"�#�qEr�������ΊAXI	*r.����f���?s�!, �8�	�-�;�WX�p��o��Ƶ��Vj�7g�IsĀ�"8�����s�_~���٧���H���xI�^x��;��Q��Ր�9�9�?��!+��G�l�3*�E&f�E?��n�����OħL�p�p���[R��Ƅ���1��n�0l��x��iX0!2�\����ׁF��������:o���τe������K�������O-��|4��b��G�i�#� �͍`��)�x�|���4�2���cv��B�"K�@�A�<�aw���d�b�n��i�W(tXk���K;��%׽�Mhg��bN���9q1;���'&�	Xp�l���Ĵ���F��3y�v�r�#7Q��h����u�����x~�)����-��Il��t���p��Y�]���������M\~^��B!�O���g��j^��KznceׇRU<�����a5:�qH<����:	ܦ"�s�p�A`/vk��W��6k1o��;�2�x%A�[�S	�k������\_�by#����o!,��@R�Ϛ���	ekκ/��B�4��phqR��&K=�s��:�����&��_��5�y�d�Č]w�Ç7}VSY	���6,�B5���O�In�$���)S���^��)(�㱻ϟ8�Ǜm���e����[q���o�gќ[	�4��p5���H���^y�v5..�^����T�����e��鲛�c�=��6����(�����o��Ád9�	d�t�qqˣ�����R焍!��k����s�Q���B.��H��#W4d���>Y<G`󻓁v��0���um��i�S�Dt���a�d��N�E&78����Kf#UE�t��X
�{oQw00N)96L6K0��"�O�}3V�\�@�G)��~o9�c��e����<��F������T�0�D��ɘe��N������ۏ6�U�Ϧ❖Y��j�MQ�3�Pf���-�)�h�ùm�<�4U޳���˷��E��7�>�6T�"!�yw�&��O@��κ�g�I�):s��Yleˍ�)���E�`�M±�~�3am���ֱ���e	
�����,(ֆ\˳|�`�e��6Dm-�J�_Ѱ�b�b�$f�6LwL�i��~�3�u�Lc$�<���������_}�J�e�,�����7�4���0ٽF��׿�9�;��8��2�}Sfu��0��X�΋.��na����?����	��m[(9�{�9�s����"2!	�LI��JiBp7�JoaýѣG[�w�)�y�lxI� 566b�ԩ֝�裏ƨQ�p�W�.��ó��egJ�)?X���t��{�>�+�Φm�p��Yh��G��6cCe�![��P^�![be�N�pq�j Д�C��T�0�����C)ӈ�P(f�;{����,Í�kC $��������9b^�!$�Vf<��-����6c<C.H���]��.����\�%Ky��(����N��� eN��D�{<F�Dc�H;�sa���%���P@2�p�8S�MvW���L�������ܡQ4gn�����댚�Mn��p�?O&�+�ȟ��ʲ�9�'.ŀ�Y^?磫0��g�(_3�Y�,��ٹ2�Kõ�2�J�S�'����2i�*Y�Ry8IT"�d�o��ZfcXB,pL���'l}�Q��䇡��m��E,p#d����#95c�2�aS���8����ǒ���޸֙��O���� �,�ʉWd�>� ���_1bw\x��?�V�d�Esn#s�qm3|+|���������3?C�fe�Ձ�d�2�������"���3L�rPi^h�A�t�;�hM29�P���n�B���k�ΐF(���@g>v�<� \D<Z�[��B&�;�4f$@L��bY�$�vg���AT�[��}����t�71�yPd%0ǂ�1�x<06l�/:�� ��W�dO%�l�fs�NB1���f+e\�u;�N�عr�	XB.OO�[5�B�͓��e8qL�\+E˱�%45-� ��<i��5�g���NOfb�����j	dy�sx9&�{w&���
��W�{�F�nFZ�Ӳy�/c�9nv�n��5\:N��-��*��(9& Vŭ�T���?�.L�t:�{~����@'5e��x����:	�1B��M~_,��9G&����|5�<��:�1:ta��� �5(;�wY}���y}��f��,T"�CaB� S����'߷�%����*������q�Ɋ	��gZ��{y=�2���;v�������UЋ��t�I.�L!ي��嗝�X,�h�x��d���z�ͭ��X�.8��n�MN8s��f�V�n��9�6#�a����}�*(��wN�{��9�xѼ!���mg�曩|�4/��n��L -b~�i-�4��N8�{Ԇɐ�ߘ����tP�RϪe������3���O���մߢ9K�vʠ]r�h"�tXz�	:�r}�R������ �@eig�9&�r#��z�������O=b�$R�u�IUaIK��/�ʹl���mns s��4��A%9�ts��qV��%��>������ NĀ>=�@o��M�,Xf�6O+�w�f4�B��%�h��ȤsH�T[��6��Ǥ�Ǆ����K`�����-���X���bsk�ѷ_O��vC�݆C�*E�cP�ˆ�����ظ�D-r�<�j�1|Ӎ�e;�ܷ6�"�!�Gj0o^#>��3����������ݕv<òsѴ�(����·hk�!��6��Z{�(�l�"R��p��7��#H��fb�%��Pz0�76�p]�76�q���Yb�N�)��%����ȜĜیJ�x��У.�|��E��QJE�:�Ut��;g!>����q��O?9���4�ݳ\:��X+��ǐ);;��<�2ea�h<���� 5t�1D����&�u#�Aa�}Y̼:�H����B͗�9s(����H�د�l�N=��M]n��E����N��K~����9�x����;����"
� 2��s�>�[3�X;��ܹ���۷�>�n�b�Q;bܸ]��?^���s�	r�#�!P0v�7����Hy����,й���h��sg�Ճ�Nu�q���������>��c���ꪫ�5�嬑�T9�:��	Z4��	�?*8��꾻�d���i�jg�0S,�A"�g� g��x�5�$c�C47��F��d�+�УgZZr�b����_`��2�L ��{���N�.z��Ҵ��uJ�(|%�d�s5ҙ���V���_,���ev�5�<�$\�\1m��	^������e�����p%��    IDAT���"_�p���}p�٧b�&k"�ʡ� �L��Eʱ�b;jkz�����^�ioʹ��h<�w ;t�egS4�B���w��Ƣ���-x���n��6���@�^Q��D�Һ؜dEz�I��)�t�U���o{��L�Q��Uᢋ�ða�!�����i��"��"JQ�o'0{V+~��3��L]��^=�8��ð��۠��N>��_o�����Ǒ�U�W߄�S���O�9zc�q�ѧ���:���ɍ,�i��X���p�ݏ��߄L��G5���ß��}z�O�!�.搨�E&]v�E��T���᷿�f�Z���1c�G������kY��B9ϹYlPfr�	���^\���ٯM�M:�	´�����YSr�If�8��~{�,Ʉ�|�}�w:�h�I<���>��S�a�� Y����$#vQ�B"�|�9����v�'|����]4kR��y[�4�6�h8=����VA� �L՘i,t��yʓ*p$�e���	~���,(A�7��gJ�
���79�ػ馛:�׃�j~�Xa�:\���,Y��c��V%GÜ�T��gc��F��i�(z�^��۸&�b���j�z�q~�r*f�`A}���8��q⏾�d"�0��L	DB:G��������<Co�5��q�Uȴ-���7�o.;U�EDb$�=Ē`B�:��96���}�M�?�*,\�A�cР^��տ�F@UMK��B���%KZ,?�mB}�����y8�?�g� dM�h�?�;�\#�|����ȤCT��@1�As[�9G�~q�p��Amu�\6�r\���У��E��I�si�riԲWU)@6E����wN�E���b�^�S�������2��t���׺���6Ī��a��-8���֜4pC���y;b,��<��zd3�9]]M��B���5ho���s���}ɮ�6ဃ��ŗ�eV_U5=��҄H����$r�fD#Z�C���_q��? �gDK	��xn��r4� 
�PU� �#yh!�E�Q|2}~���a�Bnp���5�G��/\גDW ����1˰N�3�W�R�+�>�� y�G��Z%0r��QG6K�!A�~+̑�F�ʸ~�Ƈ~ءo���������=�S��;�c�Qq�a��*�-V]*���x|�ĉҭr�	�i�?�:�2B�䌎���:s��?�~�4a: x1��#;�7$�P�T�p8J���@�T��M�j���hq't!1α��\Dw8e�H?s������y1a1hm"b�_�u�)�����z�U#�m�5� ��C*�ܹ�0����޻�n=�[�a�u��̚��u���q�DZZf���cL��.�0�����O����ת�&Ç U�B6��g]�{��+°10z�!��Wg�GC�X���2M��1x���zۍЧo�m%<�ī8�UXҔC6���5{�ګ'bذ5-�z�&L�`f�^�D�
#Gm���kP,�ha��#|:�yV�����ӱ�ޛ��g�t�^|�~2˼�[l5n<��J/'�����Ȁ�m�&���r�� �x}0�0mm-Xc���醨�AP���;����X���q���a�-7B2Z�3fᓏga����Mb�m6Š����=�Y_���C��9!�R=�f��3�����BUUm�Ux���1�3����o���,"h�9g_��S���,��"|{�m���~�T��%L�����4�J	����t�:����}n�4��t��Ym�h����5�ć=���\�Ӧ���K��l3bK����|	�ޞ�SN9��f�h�p=$P��A��Hi�_g������qq�+.~%I�좋.2y��k�5ف�ε��q��g[� �F�>]I���d/2W9��Lc&�Z��������˟~b}�+�P�Z.�b�;'N�����?cH��_L�ɶo�L���܆�=�b�}��A��5.V��r�)���r @48�*��;$w$F;P��K��?C�7��.���p��Q�9?TG;��&�AO'�"�4�d�c1��d$��`.ǃ@8Z
Odp͟.�v#6A.�Ƶ�\�{�z�L�d�l�)�8�x^k >�t6�9�44-�6}-6���N��(~�Y��������-ns�o5��c��^���b�s~~��o�ek�JF��f�����ƚ���������Ghoˡ�z���18���Чa �|�e��G5hM�bР:\s��>|]�����<���hivyc����~�t:�c�>�L_�b���
??�T|��/���)�������K����V������{����������)�DX�>������Ä��_y#^}�V�y͵{c��vŉ'� I�r��8�j�Zcu=�����м�	����x�����j����Gs ��>��Gu*�|�A2Q�T<�?;2֢C�L~7�x7/\dRĺ�Ʃ���ѣ�`�b����	���=���~솸�Hā�>�<~w�x��/�0x@_��q�w�������I��o�F{:@�*�~��4�2�ѯ�f.���G<�̋h��|���Gu �Yo}����ޯ�����t�0�v��#1�n`	K^U/�}#q�V��KVvmq�Rz�߇�0�F��ɻ����DKZ�*�Đ!j<%	&������E-�Y�_�!�.C����'̰XFr1Ȁ�r�H�D���O�֌9���1��ɶ���,̇�S��2�v�c����{���a]���29� xC���!�exژ1c�ǝ�;o������3��Fq��%�s�YҒ�뮻����4Ox<�QҲ+͉;�9��K�Y��zEX�M����&g�:�z�1��`ܸ���k���������j�`޼�h�_��O9�}0�,n����%qsƤ��8��#�����s֯���o�&5������������~���/���Q��ZD#E��.~q�9�7�?.��j\����,�b��=
�����1��٧_'��$�-d���^����0|�zx������}�a1�"Wh�O�8�]c/?������tR�)E��s~�������<s�8ӢX�aqS|o~y�D��q�����?c�� V�&��[�E���e�^�{�~
�4��#�������?���C6ğ�<��ş�̉T]\�s0f�V����qٯ�-K���ޞF���<O��T~���p�yԉX8?�T�^�6�}�I8��=1�Ïq�����g��"��2��k��췿A�Ǚ?�S�>n�z��{l�_]:��/�◗�_0�)�$��x�6��.9l8�L�Ɵ�G�"5���֐�x��̂����p��+P�Ҫ`�q5=����}�݌����s0oN����lQ ԃɄ�E L��ײOθ�y��5��Ck��K/�O<a��.�đb
�$��R�rY����$1��u��� _r�wՖ �&>������z�vN�XG"�0��5q��S��7���k��7������t�Tס�.�_���k�=��:k�i���O]3���y�^Pi�t:q"����d�,ʜ ��3��w5������w_LFN0YCF�������{Ȝ<���X�I�U؂6�Jv&O�d���:�Pl��ڶ�����>���o��C�����h�^W^�'��һ����p�i��\��	S�~�s���`�� ل���;`7�g�~��r/Z��[�������x*�)S��鍨��l�� �G�� �=�������	�͘c�o��:��ʘ��t<����=�V,�U�؊ۭ�]v��By����x��O��=�z���N�ƛ����x�Ǒ�31$Rq̟7]��{wD�$}�9�v�ݦ�&SQ��iss�V���;�'����/2�Y�Яvt�>Xc�@���?pß���y�{��:}q�O�ƀ�x����g_B6�7Y��nɒ�a�15f4��<~y�o���_���Jओ����73g�#�����
�B(�h�B}�*���H$���C��ǟ2���6�}���/r�y�������OQW�a��l��y��X���6�c��������@x���8�'G0���0��� R� �@u7�F��ƌ���M�﫮�'�q9s�1���%��rK��rDe�D��EI %�u
�ZS$I���A�c+�%�����Ep$8��O��"�����~%FWP�,*��H��K�@[�K���~֡!�f�C�|�U$)�b��.���w;�?���\�H:�k�^���*K[�e��H�e0{�\�1�/e�H㵐�04�L���ed����l:?�L�p��Z���~�;�ŸH���5N3�������mI!+zМ.��K,D2JW�+&,JfN' �0Lۍ���ią�[ٌ��̌�\��<둘�a���;�Xlfu*�	'����ej.j-�!��X*ЊR��
�B�5ep�ͷڦ�H�=��[l����e�!��^��
%;�'�mv����cūo��X#Fl�q;�E]}5r�64�����X�Z8Ya�#H0�-���>�*��y�;dm~�Av_�7$��%�d,i�0�!�K�����0��|�-6Gz���~��dN��C1����JAU��Rֱ�\S�����c���a�=v��^
]]�\9�9�k�g��h�T5�z�I<��S(3Xw�5q���G]��7�7��_�A��L������,bL����%QW_�}���bNU�&)�N��u��IV�"��a��&���x���P]�n{C�1p��I�NQ�Gl���N�P�#_hCMm�eT>�̳x�o/x�i��ɣ���י�]}Wk_����(aE������H�3}G5UH���nSK4��G �c�ǣ��r��7�҄�Yeg2i��(7^j�����r�A)�H�}�9���[C�Ȅ�͙�F���ie3y$Kq˲bg��F��vێ�@tj'�%\��+Y�?�+Qb:!���ܝ�\`.vҥi���;��LX���|i���o?|�;߱z�<�@W�&���,'�o��{����|&�0M�]v�	#G���{�P���
�X���1�ic��.7�x�̥���ȣG�:��T;0M���Q���j-0v3Ӟş�x5�45�Yz�!�c�M6�D�D��ô�(�j{{K$��G�0�H�}�Nśo�D��a����hooEmM�|ȸk�YSRr������g�J��Ͼ���z޲��[-x-�r�������L�̤a�X�u�]k}�^=�C�ydŁ�ģU���N�!��1��af.d�����m�[>z�Hs~Qv1'pZ1�L���X2�x�������G�X$e���\3jj"V2'u�z��Z�03���]�[n�dCF�q�!Xk��(�]-�|ԅp�r!Xl(ɢ6��A[&�|���w��=��M7�L���8b�h�)茲�����H%��w�Y�)NX��-����kM-;��s���Zת)�26]���|�2�8~�R�E�$W�B�N}�׵�n%g���H�k��GC����s���;�k�3,�8Gi��^��p2����/>�[���c��Q*o��jy�ąQۍ��oiT��7u]� oȘF�d���E�I��aLa&x���f�>c��-�,���O3qȄ��T����yv�[�ʿWFX���06��λ����0[��w3�ъM�ooO{��2��wϾ8�cгW5r��9IYt�]��ɞdɽ�T��I����Cs���r46�d�����43��h9���&�4���g�ex����B�؆v�	;�ݫ��ێR��[X�n��W���W_�#�<jbk���q�Mb�vc�>�V�%��/:��y�����OV�&!%*��&A��2� ��;�[/&��z��������0v�]Q
�`� 7�(#,��Ӳ�-6�.���yx
�b묵6�8�H�V��4�H�<��}۞�Uch��'0g�b�1�n�e0D�����A�LCfZo�Y�ш���x�Ld`z4"hko�=�M����7��cϽ��[wT^3�>t���8w�RLRJ �i���?�g�}��	slx��#{f_�W���E�$�I�fh]�؈Պ\�s[�1���,�L�Y�$�>�E��A-�?q��@,�:��tApϹ���ne�C�?k�~?�T�ό^[�b,���ײ�gRv��0U<F ��M3Ώ�I�X�U;b%S��)b�0�$�i���IK�`� ���d�(myUO�/s|MM&��Qc��.��B����VኺS�'x�nU>x��0�d����w,�{�P�f��M��S�*���b,�l:���x5��̷B���{6�h0ق)��x3��ƺ\�6,PJ���x�W�۱�.���ݝ? ��5W��^JaWq�����w���GQ,�0x�z��P]Ͱ%��:pP��Jt^:	f�������Q��Q�C=ܬ)�"��X�,�+�t�v�w�]6�8�;�;v�
�@b��<�Fj��]�&^<��sx���a���z8p�Cѳ��B��`	",�hŜ�BM����1k�BL���z$r�Vt��/�"P���]��8u�b`R����<tޚ�������`�-G�gى,q�R�yj��t�C5)�z�	<�<#���)��V7��>h+���X�"C|8J�
  VY�hԞ�"0��S�	��Ĭ}�/�*�Q%r.�2�a�_B�y��R3!3�M2z��/��Ej��E���w1dW�fk����!���x�*�n��\Ԅ�g�6���;Ժr| �������k2'@ǈ#��.;u�׸�0k����\55�V;���>�t&�k�ջh����j���!�Rk��z�e�o�|7�)��X��s�!��Łi�g����E�$&e��5&����:�_�p \(�1v���N�:�-���5�\Y���_���NE.ߊ!��G�J]�BV�rV�c���X91~������N�Z� ��p��n�~J�r��e��E1���]�h)��v�;�0�
Њ0RD�M�D ,3EV���A{�ox��Q���zb�}@C��(�Pv ��v��Jr,�4{�|�1�.4��X����׊�S��2�T�t�rW���@ A�<x7�}w�""�b��lC+�K]�9S���u�ؼe�&"x����⋯�>z�,%s�r��^��u�g-'<׺�[��t�D�H)���"�:�i�������*0}]����~W�2Y�d¿��/~ԭrİ��f��ٓ��i2�@�@���m��紜�dҨ����	\��:�/O���f#���Xd{d����T�e�����oO8�L�%���"";ﴃ��O�r�٬�?�0�'�|��������'N:�x$R���E2�@&�C"Ve��`,w���D�=�o��g�GU���{ ��a)�"� �O�"�Z��=�-�*�?��|�D�El��6�c�q��zư�Te0�����xO<�(ҙfl��z����0�.�qԚ�������Ł�o�h֝���_�>���՚����u�ݹr�1L�4	���9'�����a���23�1�HH	B ��� %��ګx�ѧ,Ds���Ł��L� �M���+0�w�:{�,�:�6��6��G=�w?c`ٴ�$�"f�k5����x�-���{��p��6nl���	+��Jo&aD	�L�ȣTt�V9FO}��K&���bC���~��0֊�$U"\>;����h����ҤŬ�m����9߉1���o�r�y��K.���
~�g�{-�q�@�J�\� a %k�����H%hT�?`�@�Kf��KS������J��C�J�_��<Mؿ7j�����:��KC
������P��*�;�}�|���"��{��O�z,2�8k�DV�>�:چ%.>�����rf�j4)�a~Æu:)��Z�h	�@I�d�-�G{o���Uy1jv�aL�ȶ��:�߲�G]8���7^�3�<��v��z���}͂".]�[k�d�%���0=�}Ѣ���Y���F�:�k1E��[LK3"��P.IF]\��    IDATO�ܴi�%���{�յ(���61i���0.�*av���x���:���?�PTW�L
	�1�y�e.l"����3q뤛��i�1��?C�Ym-��y��PaW��Pb='�����R[U2eN�-�����:qƨc�ni���qh9�C�ԩ���^� a����X��^_���V������'>P�v�S$7?��O��O:�W8��|g�_U��Ap�������[�"+�Za��3&��c�Ǆ�@�L;�����r}g��8�J�
�����:��v$�I+9��c���ϛL���X;c�]�2	���+��և�&�5It����~�L��\CC_k�Ds�Be�.vR���R�|��b�	sF�>�N|1s�1�C:n���0z�XP���ddtƱ6��g����cx���p�[c�]wq H3Z=�:c��;�i�/��"�y�)��6a�����|wo����i�ńs�E	�w:��;&̤��o���fs��0x�Z��v́��`�\j�cA����`�;����v��Q��F�n�:�:4����x�W_S~�tu�Ї|� �ץ�%#N����Ps�����?~��{�/h�Ƞ���m���R��G�U�c�>Kf��1&v�=���!��[��-�ڼ����\��I,��4~
"�pK�>�����_�waiƄ��L�(�b�7 ���^O�����F��'�`�����U�
��b�>�乕����?��n�ދg2Dm c@��� l�˝'*w
޴
t�������BVV�~
�gU�A������u�T���d��׹x"Țcs��#)����@`�<g��aޙ��y띗��o�vۍDM�7�"�;��,یBgqmV$���v����|��6����0�5��$���='im�K$�� |{�[���f���κ�p����$A&�Yh�����:l�����&��ʭe�/F-8J� ��:�!�����|�m�PS�[l6���6p)WsN��~o;Ν�ޙf��'�����:��b���(Wi��R���@&��O>6g(+�54�[lf�4	�iv��|�"�ո���z���4�୷�FS���l�a�ӷ�1ב$�u]Fl�c�W��ioǻ��f��߃�\Á|YEp]��Ȯ�5#n����������ˌ�܃0�,"ʝ}	����}��+�o��6�Ë"�b�>�7������w���>+�\j��	&�ԭ �ى?ԫq��u��1%{���s-�����v���)Mƿ�=Q�j}^Y2~ڡ��ΤA��͔�8�?9:ƃ1�1.�"�S���5��+6�����bE}���L�B�ь�l�����v��&:�Lg�p(&-�>`�VTUV>,A�=SDUu�����QưMҊ)����k[ښ]�*5���3M\' 깱:�cîȓ
�3^����<��	�S�����0��=,�M)�oG,H!
6��Xl����խ���uD��@�E6�⅝%��*�=�v�p��+shl��64�%Y�k�i�a�."t�#y�-WQ~?�X��Y��=;�7Yk4��k�8vڣ����
�	�s9�9�)WX)� mmtF�.��"C�z���;V���Qu��#X�Y������8��J�}�O�ӷ�eY����O������ar6g+��D��Uµ�V
Fu�7����\{#G�+���+e���H��i��X��~�Y	��_���vl�C
�r^}�cuG����r�t�q�c��/��u�y��Gz���g:�4K;j��v�0����`�|�g�H	7�.j�	�e'�R���s���˭(���R��Ҟ;�
�w� P�K�"��pz�����d�K�#W��%���ʛC��7�-US�w1͝��ܚ�l�c[���p|e�	��u-]�}W1��h����z�����]!a
Q(r�3�2��QZ��}�\y߹���y�h4���	N�V&LM��a�X�av��!@��I#S]z�;k,}}�����^Y dE���Ү��U�B,��n�:�@��emB�{>�𿿬��i���X6w�������0�<�\|J���;�ry�]�.!�+3_*�ϲ�>�,Ӻ������蚻����o�g��i��@�oS}~��|�h���g�>��j|�N��RZ���τ�ͼ���:zy L�/\� �O>1_]���R�v�m���[�B�&O,�ں���\+�,|���	��]�ݲ��r2��}���X�;�騩�'��D�s��%�2��د��WW����_����9���|�>�?s��k<T���-P�wĈ�ch��y%�O�c���W�|�&|�y�حs��3o���6���4�r�����)��O o� ���=|�lK��nQ-�~�&�׽��YWLjy��
<W����8�;�oو�빗'��^�2?�u���l(��X�s�Y[%t5?���|C�,�T9����D�#T�M�$�h�?ʟG�/!�X�Y�ڴ?g���R��{�'u+3m��B�	��Z�</��k+5-$1�J�݊��R��`�;�����}C���et$��e��������|Y������q}r�U�Sy���돕�/�[lV?�?��_��+��O�8珈���	l�3�������
9��F��KN��R�,��s��I��֑�a�i%�w�7������.e�q��ޮ�F��Q�
C|����Vf��_���W�����W͕��(��sU]���"��b~0�@T���7���z��������r���խ��g�v�X��q��ܭ=�6��C�/�u{}�u��@�2�XN�P0�d`0�LqxLd��L�L�����Ϝ+M3��W5�W�����Y޽�*��e�mE��U�~oY�te����o�g�.��{�:��M�n�cޏb��STWm��L�+�%�7Wa�:)�H�2���,@ƚ�Y#|Sނ/i�|�b�H&|�E��[Ax��g�װ�Iu��m±�Ӏ���5�ʾ1/~��@i��a�(�]�|��T9〱�o�5e9pl����dG���T0^ނ�	�������u�/ouu��:��]]��t�	��*k��ݿ�wI�Xs�䎅���&��}֩a3O&�̤�^ͻxh?�B�	��|d!%f/�>_�G&P3��UӘ2�^s<��=զ�@x�E]��n�MN8s���f�R�k�jQq��V ��1�����f�a���V{�`�!��y&o�i��Q����,+Ț�
#Q;i�]u��]�۳Xw%V�g7��.��O�0������*�no�����#�F@&?;�����	�lgĵOF��cc�I��8C�&�BE�+,�E�`�`�5��B���bb�AbI<#N�K<�=U�����y ~�\�-�ܲ��<�֎��S7�;o�M=�V�PB*�B1��v�l�]w�Śpr� �U�y�BJxAܱH�Y��Ay��g��B��~rg#��L�gђ�>��w��3����*w)$�������J㑘��v�4��`����X=�� ��{��h�����@J�5u�T�u�YV�N���׋��'���'�"�Na{5Ue�3�?y�-{b� �?Or�k�q��*D��)&L�^v�i�4̟w#��D��
1�1z��ǖ�l�-�9VJY�m?|�]�D.��7�Ϋ�9�2�Ѹ�H�э�{�<�䯹�c���ؓ��m���G�?��J�p�k�M�_;uV�m�����-��.��<�1b�=����=(Y���+�4FK"'�� I�H�j����*J����ĺ�C��J��CI���5�᷑H$O>���O�V&��N:�i������0g=��F��9���z�V�a�м�	o����=�
��0�P?��7�B*d���s��hj3ou����47�ݔ�̎�,���&8���oM���P������zV���~H�Ȅ�;�<�)S���W^1��l�w4)����aGr��[}�X�/�j��v����e�[�8�7��|Q$�$�dƊ.� �A�}���� �gќ��m��Yky�]����i�ѧ���[vA*7I�+�W��5��;1ی����R5xj��A:��#�	Ҫ%L遍?�P�;�\~�pw�����3���#��� ʾ��%�p���Q�$��_�����2�
/��0t�P+JФ�K�!�v�������}=e�w(cЂg�]2r�����ly����� ܻq��#�m�b��Sb������Ǉ��?��#��7�~����y�d�܁�w�d���Ȇ))(�[�+�Ѥ'��l�i��&[%qP���Saq|�����X=��#�g���;�Зv�n�ă���o�%���('���M�GL혟q�Y�
;#vH��(W(m��S^��x6y�d�)|
�0���<��s���[/�2��Bǜi�o�/�o�Z��B	}k�X�چ<�ק�7w+^$���YQyi,�$��N�⋀��3�4�=��y;��q �w+��������d�qJ�)��|��� w���ek�gW����׎ q�k}�]v1ٓ��H���I��7#���0?O�ψ�A��Ad�����^)��O,cH-ϧ�3C�Ȉ� ��N�9A8�M�����#F,�2��%�il�!Ѷh/���N����/��q��oܕ(^��r�� i��	e��)�[�k#G�4`e0��;��q�g1}o<�!��t�I־��=w8�<�����`��Ϫߙ��Y6rU�q�qW���pHA=�@K�E�� ��{v��������"��ȓ-��s��̗���@�Cď�%&n����o�u���������ގ���b�L��s�9��
��ƃ�̽!ֲp;�`���c�=�������g��5O���]���y3r�|. �勃�}�-l� {�-����;������8h4'�B����կ~�O?��cpy����ᦩ�����.���R��Z�l�cA��ˮ30�Ė���x�ڳ�;5�/6h\�� �M���u�*��+CBW6qey��5O���^{YtgX+Ca�W���β�ӧ���B�����a�S��B+�@���
'�J��$~�	�%q��=d��AxqӒr��A4r���N�V9�q���ϻ�>�ގ!jl�2b�m��|���2>���fk����x#�q��͟8��f���r���;:2�)����8�ṣ��[����}_q��q����zt���0�l��;&��^w�H�QvSP1qW�[�r�B��Y/�Q �=%��`�)�篁/7�2�_��LE��s]o��&8ꨣ��&����QF�����]E��u�]�鐣����'Ű5ʜ���v��9AX	�Hi}�w&�͙7���,����Ϛx�O�n9���5�1קq&�5F�!��n��6�g���ן3&LM�J\�㖄A@U��&�@���]L@��ɠiV�'��� ��F�X`f�q0��@�m~���|2a�t�	�Ond�����pvt�X��B�t�DZ����Q	�r6̐����	��-���?wk�OY���������Ĉu�w�u@�r���&h0B���O�x�	�%��\�#\�N^-iʝq%�������!���Cak������9G����.�J�XL�x�ğvktkG�Y<떪�f���^d���18`L��m|:�S�J�1a^w��yy��&rGVlވ#�D�A����$�g��[o�մ���ƍC�^����<�b�<��/1�Ck3S.��q�h�%O��w��d�aW{�͌��	I���6���������_�{)�m97�^^%D}�+�j�U��/���c�=f�!��W�ċ�������R�$�aZ��I	hI iE�	����+�1;�x%�q��M�L���#A>�����v���3�l�s[�y�H��Hk��#�8����7_7&LV��߿Gș�U��w��F
B	��9m�4�9�q?��Qf޸^*�̸=?/��/��$`70}�~�{�i�1���v�i��[	�l]����>i�)�ɰ��Z����uG�g���(�9��Z]�]׷,�^�����ծ���8��LΤ5L��+��{�a�7-d:��������ә���/j�T�A�O�ϑ�1�B �02kFy1e�5��q-D���	�׽!j������ϟs{u{�1a֎�]��~�j����!Ӟ5�w,�0���
j�@J���\m$�=�`�.F���Xڎ��aFI��/A��#$�|P4T�G�+��Z2�=�uK��O������d3���b۩W�2;���_�u��d�����XU#  ����-"K˻>��I ��</�</#�ԉG;��~(�Y��zU�	�0�	Ԏ������<.�%��\"p$yLS�̡R��5�>f��~��b����h$:y���u+fg�>?�T�K�
#a� ��$��;`�m7Ō/>�������f7B�T��2R��<�
��	�a��<yS�y��J���Ȧ�"?�~�̕��#��PcE��j�	���;`e�x���.�l9��٥^�Ć	��Bgw[�-Hf;�կ�#�*G@ �*������Yl�Iv�'d�
����U��N�{�)��}衇h�5~v�t\�W>(���+�e��~��_��&��A\2"���0U�̚�wx<5%�����ǟڭ �s��̺���UB1(��1d�:�k�=PSW������wA`���0��@%�̙!&|��ݎ@;v�X{���u��-z��yY;����2�H�2 ��բ��Z�.�
��9C��|��~�����׊��� ������,���_u~����X�3���yN����ԕ5�c+ոJY��{t�}��Cɒk��	����,"�u^�{&`�ES��ڣ�I����}���x#���)�-w9���\�`�*�^������U�x,�(�B��[�w�}�8o�O��n��!�F�q x�����(Cpp1AmE�9��E��jIȾ��:Қy��c����K.����_<_��@��&P��(˲��(r�J����VԤ�(�ӈ���C	���x4�I��A��kH�CD�Id���X�C�E#�J:3&�/Z�q%��Ǘ�Rc���{��eW^����9D��k���/���l�%���&&?�0C5S��<�N^�B�����ɱ�qP'��b9u�<����9�8Q-:9p�hx,��j���gxG��+IH�m�13gy�^����]�@�/E�_�-eUE"-���|1`ݏ����4oI~�,�"Q�X{�n�߅ߣ��`��c^����sI����4?Ck����� ����Ngc��M�_� N)��=�e	0���%��!G�|S�6�(,Z����<_�a4�<aw;f���|fT�����r�G.�E�=��C1f���drvQ�UGXT "vJ�7Á�.� k�&����R����m�8��=�<���ѣ�L�����"�'k�æ�,(;�J�!�L �s΋du�]{-$�r�6��@��A�G��C,��T, f�='i�a�)`$�L�5(�R#	�"q���b��/���D��q:�GhN;&�tj�9?R�c(p)?���
,����n1��k% ��Zl��$�Ȝ��;H��.�w8�A_תI,�����ܼ_��.��k��<�ǿk����Y�k3X����k�����>��L�x�zx\���������� �����5�s���9�
�d4��|�o���ᤵ�Gh�&'`�>�(mꚣ���_�y:�&L�`>'1k��X��n˪#(��h��}2
�X���#��$�3=�_�Q�xn���11L��1�U�Ԅ�Q�gFK�H�!��fQ��QU�¨�Fc�-���4�$-B�!x��#L &�gf�2�v7�؊���:������.�IC�&�r����	;.�'�MdO����ۻ���^�߷J�,b����kò    IDATA1ӌ�TD,( d+ˠ+ҝ�n4@�!ϱ���g�%̚=O=���'J�gsK'y��X�A���;ݓ��d>;Hs��4bv>��ܠ��yl?Xݟ�Z�:������E�+pҵ�!�ϼ䑖�������siQ�㦅�MC��B �3>ȋ��z�U��[<��z)�Ō���i�����|K���;����9 ������_�;Z�*1@B��?��dA�ei�iMi���~�ZW=?րa8�ψ��+c��\</}G��~�9�YqQo�~�$LY���y�_���)�L���\�VF]�4ymd��+�?��12��f mR�#�s	�t+6�܂�'�ȧG!Z�DJQD����@8Dd�Æmj^Fޤ���<��� ��:�-(�s�%V8�v]NID&e���������gQO��gpZ�2y,d�l/�#UUg�m���5����>j�QD�,b�,g}�|�bD�A�|�-GȀɎ��A1���$�u��{к�*J1̞3�b�h��	�st��\�߹�k���$WcC�6mP81C�r��g��r��4�Z�3��bx��Km��p�	$C��\2�x�ƼV�u���d���g��|����Q�h:�3c]��bi���,&6-0��ߠ���%	F�6�y]<�����1jc�t��_�9I����6$_,_l�1�$22�Y�׿�u�s����Z/��R3�5F���/�[QQ�L�o�]�$���J\�u1����\���c�g���f˵ 4��q�2(1�:9	²��L9&�I��aj�G���ɖA�-�)Gt?�_���5����H��cH����e��0o�L��7����M0	�d�d�
�֮�3�b�.ԎD;���Ŕ�(��w��9��N��"�Cј�-���nM*���$�!baI�?A�u!�p�B>�agA���l4�d}��]��a�D�%��ېˤQW宭-�-gй<<�G���z������)U\��@W�T~���h�*�G�\�W�'�z�o ǌ��.m¾i��A�����'  �3bt�~��Ѧ�"ޛ������R���6+͛J�Gs��)�S�S����޵�h��f�w	��}�XkbYSX?#�Q&�/���;ǘ����܌8b̫��y�U�r�9
@}k��'�+
��:#���ճ��7�a��w�'��K����l��*�Z��z�x�}�!�����ƨʣ�<���K��DC��嚟�&�{Ձ��ųn�J7���g=�"3�J(9�9k�IMX )-�T^��L�@@9�r����Ap�5(��q��C���~�>''���ٺ�I�'"�DY�ǙjټC2ՓN8���,�����y�GrHF��GX�����&E�"U���G��C�A� ���g�m�H.��]{%��i)p�8�b��G1+���.����)9F�?�	j��y�1�D@����5���O�_ % �=��@Z�����{�b��"y�b�bx�C� 4|KJ��a���MJL�x�t�bX:���Jc�U:�ym�E)psSVKG(�')H�բ׳�����32�}��e��� L f��ƘL�a��/��Ȣb� �0?�Dd�g��dº����>����R!�3�j���H����Ot����";ڀ�1K=W�O@��#1�H$r�����n�#�ַq��5��ѥHj�t��sH��h-��J(�d:�db)(wPj��G@�7?5Ȋ��3M��	[��	�<f< _�^:��qmU
'��X���!(��D��>F���R�H�@8w����W�"����*����ǀ����&j0{N����6c�,���uf�UN����1����K���D��4`91�zeJ�C�����O�e-Mx��򀋭qb��3�$h�Y�(�c�͚�D��1�{qI���6�JYC�$�3�g�'SK����(V� �����3�ߡ�Y�RR�\��`l��DF�y/=R�K�b��d����\��~�z˓���x�rF�=锲$%}h}�F7?K}���63�a(�֒,��7�	��#AX�Cf}#2e�u@X���!ه��¼VE�p�@+�����z��X5�-��{�UVI�M��'vo�9�	�
s�)=���9�	�YR[��<a������;b�S�����0�]�L����vP���|M�Mz��vYǜ]�xf���֣�͵����5�Oŀ|R���E�0�m��wA��;s:��F�(
�8r�v �}dP$k���9���;��ڌ�:gfs4��"�ܽ���J(Q�F�C�z��ۏ�������q�@I��u�x�g3>�3}K7�Gm
��٬ed��0rYT���1����v0�e1b�9��tJ���'k����u7���6b���X4[� ���,�5p1hް+�*IKڈb�� t����dN�\�!��y)j@�7��	�f.V�{�Kf�Sg	�Z�҅+Mf�:5S��� ���6TW��*�z��n$6��9�Pda�Mv&���̈� O<��������W����xɊd�e"�2���j`�0&k��W]uUG%2����,��{d��X����ؖ,bޓ�
��0a~VdClT2�oai�hu�)ʗ/���z�Y�֗|�o>i�����]���~���lp�E3o�˷�	3�@XrS����v�x����Â�l3q�0���C]*@�Ў�X4�S�ZQQhkrR�̲� -�56����꾨oX�d҅ �-�-�݄L��h2���3�dA,�W۸HG_A���=)sđ�߷�*W_m)�A����j������'�����Ҏ���(����!�T}�r�T���͆�[v��MNV�z!� N�H��1c�
{~I�P1�
�z�.�b���A'3W��En<b6��8�`Դ�V���E2�� ɾ�D-�gs��|-�s��&��Z�~��YM�m,0Es��O�\9En�ǝD�����;��$�Bi���"�K a>�L��=��ö��6�(#q��Ŧ۳�Ɯ��ᕱ�}�	���4$x�R>[�6
E#�|�w�H�R�u=̲*�3j4��a��>�|�$��lvQ���0:�@�M�ϔ��b�e͊l�֌��"l�IW��V��/�7�,DD�'��}���ϜT�k�b¥0�D�A�(��A��e3EuU-�%uУ�?���H�J��H�rX4�sZQ�(��m�D�\!�=��C�G��ꋆ�� ��H�c��p!n��f��-b�bQ���؋ǋa��ߣ5)d�Z�7Q�z8����t�*M�|�Y1`�Ǥ>�|n}�,nnǀ�^hY��h�X�HU��WU,�����"[4�|��OF��� �����R\�t��i��1�`�c~�,�)�2�|�B�&�P�! H_��%'��㎎��iI ���L�U�L��uP�%8��әK��7�LXlI�?+�t��zv\�L���f]Ǟ�B��g��ڷ�$���<�A	u����l��{��A���� ��mDt�K�|#� S~��6��$KE�	�L��%]��Ra������ޞAX�`�6�bǝw����0;X�`��'�F*)�Q�����t�k���. WFW�� ���u����n-eI&�k����r���'�0�Z�ԆY������^=q�1G����@8^hÒ��5�G2Z@�o��٣c/��(��#F��xOdKI|1n�<	-�f$���������K�!�Q �Hզ��V�������=� �4�d�z��"U��d�C��G>����q�K/�1S@CMo,X� A,�h2@��|ɠ��ȡ�6)Wys����Y��-�J"��$)�D$h�*١X�LaE H�g�"��Tr��tlNx�:�E�����@�lS�"8x���#��1|���^���f>ٰ6 9}V �}�Ii�78I�E	Ѻa�[o�m�#uM%�܎��JX�F��f�=0hض(ī�s��{��A�A8D*��Ի��{o���C�TD!�6&�.R����PʛdUcq	�	l�Ŗ5f4���s����'v��|�F1V�JS��,	��P�Ed,O^&\	�����lwY��}"�췒i/���~��ğ��8wR�c���4&L.�6�:���%�ƀ~8��г�B�b+Z�A�e!⥬1������0̣�h,�S
jM�F�~��C.Z�s�b򔻱�y1��q��gMPR`̲ix�� D)(!oi��tc��>m9$��PM�:,!��S���P�GQ����x�g硵��d=7��\�R�����L{�@cƬO0�� �"$�e�E�i�I��h��?���xb�2��td�<.����c�]���`0=�%���RkQ��x겼F��S��xV�"�&`�$XW:_�=�`��tA����w�I7"t�^�9bz��kT%Sv��=�gϺ�&YK��JƐ�ŰU����2��8���=_���{�m�Y�m?3���G�rS�q�ؒ-۸C�B	�I @�!���mll�d�@(!(�dzI���EN�Ќn�V���g�������[�7�JG���^K:��=3{�-�{?�S�(�jT���$Km0j��;�i���[�����)�T�6��[��p�H��Y�Ѧ�����g�b]r���P4^i��h)��D��d��[�uB�u���2�� ��2��Xnx�b@��k�yӲFG������i�*�:�vڭ�W��s֟e�}=[�	��Qk�LYbL��U�ȲV�*�)���s��Q�������f^�<�ݣcv۷o�Fc�z��g��LN9[ъ�J#�f�Yg���bv�،��Wm�=�b�i���k[�8�Vֲ�8��Z���������3h�S-�F����6�w����A��G[Pl	�n#�G@��U�d�3'�z@C��rm9�4��A?�Ctar#t����hRć�#�ع&Z,q�8��Jb`�S ��B�)E:�9F;8������(L�}Ӗ�V��`'���g�� ?0�,0a��jZ��n3I���m�IgYr��7�1��-+l��JT5k�����'-{�v���oي<�z�9�U䈢�*�~@�RK: \���䣟d���lk6ˆ�d'���|���W�򕞶���G:0񼴷�a�ݖY7��!_Ch�u����1Wh���/��l��B�|0WB���8�p�Y��n��5�-�Yy�~kc�Y�6�Y���L��t�1*'�3Nw]V,��-'\Ӱ�����3]��ZM�R��d �d�֎�Z1!�����۱3��܊�=�vD�� Hcڦ�Bt�U��HR��+�?{�:�o����,�;8;�-b{ۭ���N���;�� D��Г,Sق(�Pk`
���h���*�H:3��}J(@b ��������
`ܔ+�a���(��)����a�Jq3���M�B�V�ݚ0���=�^��ㅯ!�o�z!=7��g���C�����$ɭ�6����R�X}��x��O:�F+��N��.�D@Q�(m[�N�l¢��nw~�VYfլe��3a䈘�R���zo�j��ѶV#��Zݝ�ĭ���XgUl�pᢧ�(����i;���B�*ڡpt�cN�7[�/6��~.�\���^���΄	Q[�}��_d���*hmIl��?�f�Ǌ��Da�y�H�(v�H�R-�E�7��DY�'����L�u3��jQ�|��#�05<|$|�����XEX��]vb��Y�=y來��l7��6�YEC�]S�Z���^9l��%vOOb�굶s|����h6�T��λ��{���#�p<@IX ��*��2ay�(̯�7��	��pi�������*��sТU�[�\�ܫ��Z(X8�)�DV2!ll�%�P����c�=�x�M�h+ŢsM�?2Lx� $wռ����m�1e�(�f޲��^Kk6�w����*ǜbc�A�`���|D����ylڶ�ل%?�7���;�*ʭ�6�ؔ�@��U�"�u��Z�8��k7���h�V�pPJ꡽�H>�l�E�Z�X��������ąLx6P�n���ƈ�,#c�s��m�4�r&�_��w&��*M�1�8H �JR-k����{�e��A���L���DE��Jkd�W ���L�[9[掙��s^l$
S�xm�E=l��;)��I#��rb��Yê��f&XےV��%�Ț�������M�׬���S^��E�Iu0�T���������1v����Ģ>�X&�H)��b�ۉj"t�AP;���0����~Z�q �$�0^U��>�~Ђq��P�ó�F�@E�1E^���LZ (|�@ AX��3�p��IN`�y�驤XSN�p(�~�?�Y~���
�iN�L�p�n���F���;��;�b@8�f�j�[W�9�@)��M;,����̏�k+Y��/�ʢ(6v�a�FMw�E�;D K��$�Z��l,����Z	�G8�e���(Е�p  <���3�X�@k܆��{A*A���|�;ߴ~���K����}��lot�����=zzk�6C�Ll��aI5�v���bbk2���H0A�x�Ҥ�t:�I���8K����7e 1��/ ��F��bma,�B�Q�g����N�%xiB�Q������#�2��ʽ����,.7 �m�V���p��y .�//�<�xFb�7���qd�8��$���#v�Lj�b����641i�ֲUa�7�'�nq���m]�Ҿ>��ݽUk�$����ε������w�i���@'��{r	��")�[��_K�l�?l��
�(YCq���tb")���&�⌹&�Z��(B_J�XA�@k��8�c��rM ��"3���9' V�c�.����yV:9��]�Ŝ��z��"���r��s: <>1j	�0��hV�]�j;��-;���[#!�0r���"����#�~�&���3ូe��I�Va������=:ك�� B�<=ȭ���hi�b�J��M�҂$�J'�g���CR\C����!g>�J��`J�	�G����u�	VI�48�8�q�g����3g$_��$�ʢ(���W_��e��󪧮ڽsc}rt�(;k��d�U��i���� �9kPiL�T��=��T:���PcQ��������I�p���|抛�(�,Ei�����\��+C�<.0-�u0�D^����ck�2S	05�`_��L,C;�K������+>i�+^]�ZϮ���ɦ������)[1=i})Y�5K���"P뵑�j[�ٿ��vgod��56�hYk
�m���A��������1��O��b�J &}�s���9C_P�A@XrD��uX'ז<!ǜ��ø���}#9���o��J�a�B
��@Mǜ����M9���&�x��yf��*�IG�� |��g��������y��Ƭ�vTV�aϾ��Gg�!�b�UXЋ�9���r��|��;�a�w�����YA�R��m�3_�԰�,C+d��� S��?~�l�+Q�#�t�<�,|���|�����2q 2.�����bb���"s�EZ a�2<��5TIN�͵��+�w��qM�cT�L� PO�37�|�O>��=Ky�y������ؽe㊬qN��0vֈ��5��&�њ���!;�<`g�X7!���r?���`N��w�k���^��luM]O�Nb;4��ϺW�����S������ߙ�Ej(N�"5����e��bLg��'~��LlX	&3�h�L-A���Ľ�!Qɬe6\1��kϜl؉��Sǧluc��r���qݲ4�
��R����=X��=�5KW���f��F�z*U��11:fqT�;����n�>icͻ԰e�#0py���{��/�jCK��`<�s��ń2�=d�jG}�~���u
�	b� �r�s�	k�Q<2 ��&��Zs�ZLx)Z�Ϊ眹��䞞>K�G4��k��7�m�ն��Z�l�>h≉� B�*x[Lzs�ik�qK������_�a�+B    IDAT:ά�Lx���.�
��y�c�ѕ�(�q���\"�]�2���L�tiG�!]Gc8�e����g��RҖ�<�'��3���G��0Bf#�r��ƪ+�xU�6,��kHW"��-�c� ��`�9�.Ϫ�'�_Z��o-+��Ʒ<}�ևoYg�4[3��*mt��ƛ�6�r�w�8��}��	D�p��aC�J(�W�dV0������En>��shl�I��ƕ'�c�NM8�����:&�âZ���2��yf5�s-�w�Ee�����8�/@�-k��������<�j�bY��n6�Iw@�՛X�J��C1j�6�vB���	[9M_��Yw�fy�I�j���j�eՐ}�?���m�g��pD��(���^�!;K#��]w�=�����!��Ć���;��X`X�'lsZ:�"#�%-�0�r����s/��:�/9��o�y��&�D�$��!˓#�+:Bm��<����WY:�p�U+�r�M�ŝ��l��$���yVԥ��=QݶWW��g�o���6�5��}�0�p��r&����6v׷mMlVO�	�V�p��I�ZRK<��,I��9B�/fZ��j8�$H,�I����T���F�2��!��31z��1NȘ�KV�|f,���
��(8¸;t,Ϣ�x��1a�; ��8�.�A���1w�7��ۧ�z��B�~>/�Wmߺq�=s6�%Ӫ)�vf���ο�v��s<�3�"N:_� �י�Hc0�y��MHb8:^�N ��_�r_� 0�I�ɤB��%��ΗY�Ux�FaPc��i� �@z��ib|��ꕒ�Y��u ` 0�zp��9���{ՙ�0/t0IRL!�D=P���P�E�q�Z�e���(�ά��6����q��N�b;zt�V����ܹ7��"u��V�j#q����G��p����nzl)1�+�\~ ����羻|��.3�A�5�e�p�$=�A�R&�,�V�VR���h�0i~�@!�HÄ�@Ӷ���9�c! sK�~�P�8TB	Yk��X�@DdA�SCLXKOq�L`b��)��n�f�Ln����B�Z�z�e͆ō�����ڨUmGm��~�y�>�D��;�x����<ށZH������6qwᘫ�g<:u)��@f#���d��#3>oD���n���]�նZ��8u��\%iHㆶ
��5O��c��}�o_��/~���\���}�+_��~����N�*���T����¤.R�T$���*�B�,�|��jn�xd���7�p��.+?��o�ڑG6V���'���i�0L��S��_~�m|t���>/����>���19�ƈ��Y��>`U�+�6(c/zы�)��G��e�]�E]�������*3J%�h4�<��I^�:#�2׿�,*?�9l�� ���֜�4K�V�&�jN�X��
Ḻϕ܁עj'�|�#�^�Ɏ�[���n�z�)�@A�Z�;J(��<@��8��Jl��{�Ln��96i�hR|���fI'�8��Zݶ��m�����F��A�k�SO_�;����B���N�Lfm��b���e *���{���߀%�(*|M�H *G�E�����9��9��7,,-Қ�_�V&�駟�u�x|�,&l��(�M ��ϸw@�	��Z���!'�8�:���d��C�Y�6rWR$k G��i�*��k5��-����xT��a[s�k��X��P��RƓWHB��2[�OYv���]�)@8���̤3�F;wn7��q*�t�Z�f��Z�W�#���!�VO[sjW����_���ojk��f����ox�k� -5G Vj���L����m޼�ﻛ ҟl��6i�3@��f�ݒ��?�	x^���Y�X�p�e��n��e�5����[��
��v�QG���?r���w��o-��{;,��W?5�UޏI�C���(���(]��X�^���yN;�E4>�b&�����B���U0�7�Zq�p�6B�2�bxp��^�[�j��֌բ�Fwo�tf�z��5S�	(N��׏�#��_�j�U{V�>s�nY\�ѱ	V�zO�)�ӍbK���8d�,��
�+�<ڵ۞2cvR�׎�lZ}|�b�����H4-gq���ց��f2������Bz{|_;j�o������% ���X��i����l8F82���Ԏ��+��\e�J_�0�BU��b.���{ca��6kr��z�#��Jh�,�b9>a���l �ǜ�qó;#$��i�B�pʚyX�ӟq��F�аM�O�Ӭ(�Z�I�؞dȎ:�\��z�M��m
*��E�G�,JS�6m�w�n{��^'� \DG����r멱04,�&V���i��}���<��x6��H��L��]N�l�7~�7|�-��E�J@ZEj�[,��_z�.�^1�A�w�ĩ�'`c��������Y0CkJV��Kƍ�+�2�@̳R���"�Jy�EѦ���=oYv^���[VX�l�S��s�s�=�%��w��_���Y���		�0��L+���xp@g
��AC2�1���a�����}��C��9��h����Š��`>��a�l�]z��G���/�'���&���q�͌�X_5���������C�En��cK�VZ�w��9�ҨϲJ�mٺ��vl��`ș�4�d� �}a@ވ�	��;fϬ���k���������ӹ��"���Jl�(��������^m;v�q�kR;��f�w//L�'֣	"�U�}'���[d�hb��É&&$`���'��	�д-�v�0�K��5fd��J�P�eq]�h!���a|1>���&���Ҹ!I�()|d^����p�96^�hj�8��{��W�cםg���)���L�2�"�-�2�[v�7��v��CF�JɄ��[����'���S�̼��I��r���g{�lUʣ�� J �:�SI��A������O(,���bA�ve�/��kQ`�,���2!�n�G�w��#����y�+�����uñ/i�-��<��[n�ſ;��Zqo��޺� �&�r�#W歳(̀���+m`u�}�;���W��a��d����Lh|4���Я�6��)��P��.�*�'�U��?�4���ц��|zp̙��:�T�V%޹�Y++6���^i�}��OY_���b���ZV#<��"��`E�,i�YT�V�g���6t�S�	�}�m�۴i�kp}�U?�A�>��ĥ�I8{ r#ʭ��cy�i�Ql�񫯲��,I3�խ�h�C��FaS��Ib?ٺ�>�7_�Q�SkuOÆ�T������r�䢋��O����ov�e�+>@S&?�$&JOz˖�v�Z5!�N�<���Pp=��U_jr�R�0��~ ���|.0��%	�����31D{hR
�%o�����H��zv�AD�_��0{�|��S�*���l�ն.��N9�,�)� �@�"k٪,��އ�����o��ﱆR�0�"�O��S�b�؉	vN<�?��Y������7�f.���~�ɳ�|��ޞ�J�ô/ɋ7ݏ@=��5��7J�^y�΀a���W� _|����Ӯ3|���4��}��?A�+-6�2��"b9���X�`��?g�@�Y�J*�[n|���� L��ac[7�&F�A�t�;�^��+m��#��;~�����(:����3(L7U�X��ѐ8�ІE�FD�{��^��0� ����]t�ׇ����+71�@b&ZqC����o�Z'�b���H���׾�56�_��9a�q�vo�w[o԰zJ�Vj-*�Q!")UL�v\���[uh��}�5}��^{x�N���M���E,1��AQ��zl�G��qbc���]��W�ꕫ��V�p_m�\�E�-����s���s_��MLO���a��ٕ!q�6��"��9���?�R�ir1�Y@5�Hb�$��N���`�i	`��@��� �P؟�����LL@���/�R��f�x���*$�iBr�7�����P�ǽh�`�`�!��E@4S�5�,��Tg�����}bi��.���l��ô�
Ql��X�S�ǿ������bl�n���.��-X|faYF\w!�M8&^�s�C��������r) �͸a�9�?2�{ �ō>`<�7�^��=��p���M>%�@�s�0�9xE8.��x�,li!4�j喛��ۖ�׌nEv&c�Y�<�^���m߻�v�O��-�='��	;
C�ԑ|���ʢ�����'?�4�������C����װ㗼�%�z�������WZ�
�I� �k_w���,jOZ_Դ�[���3�,oY���WN����.�78�i֎�����m㭛mz.kΖ �a�Ԟ-ct�I�{ѡQ��e/��׮-*��5o�^ �ÌjUkf�=�Ӈ���w�w|�������0��OHL@&b�F���߀_ ,p-ڭH�`p�4%��Ľ�ó^��	�Ra.��0����ώ]+�HzF]G��k3I s�0�j�r4�Pa�R�`�O���-a#���cR}�A�>i�ܷ&9@����������j��6�(,��Ͽ��F��`X����	5qa*;[����}�KvםŶS|�K!!x��$��\ �yC�Qʲ[�AX}�O1ae>���L�s���H�ā�ik�,������Ɲ�7c#S�`���i�a<�	��5|�w3oX�q�M�ZZ�$���׽{y�0s�[޴*J�z�}v�ΰ�/��~t������Z��0/V,4��ix
@�B+6�0 h:�������h<4�0e�yp&:�R�Ť�o
KÀ<ڠ�-��R��e��j'�NF;0�g���W��@ݬ1a}����齖M���j��r�mO)�=��Mm�aFT��/v[>�ֈ������#�3�.G(O$�lM����	�31�/8�<[�r�O�Z\+��)Mo�x5Ҷm۹�n���695U��E������	�~'�|��4O7(3��7���a��'&$읶���/Vǳq-�$\[{d�v����=�هLD�Tߊ� ��������sM�	��XV���Ua���!2�CV��@ L��D���}�z�^CB �~�m�u*���*#�������I�:ŭ
^$���ʨ�<���۾ioy���2�C�`6f�O1aL�n�%��d.�{@��B9��º�����M>!��,�ZHO�Ї܊�8=;�#9��4Db��z����g�a�ϸg�k����/
�ݺ}���fd��w����6,_��#�<�ЦU�n�iLu@��+.�0��V`1at~W�Q8x�O|��	 k�Ya	�E`R���/v�ba1���\@��]8K�9�8����u���V�,jLXo���	WҦ�F�+��<59��F��_���Ҹ�ޱ�6}�3%Sͪ��@��͂	�l���SE�U+�}�+
Lګ�� �9,j�T
5���ωC�V�l=�pk��*q��Ԏ\SN�d����3�8Ma�:`T&c��,_z):.\��59��2F�L��Ư��1�c���Ɛ@T��1S����!��$�;iC�_1M}�x�Ox_YWb��a|b��O	-D��g��j��	Ÿ2&t�.��-��νV��-C�_	w[V�H���ń�����aڌ���:Y�a�� �d\ >K�v�%k��
4��|�!t|���j/@�fQ�V|/�@���c�nYv>��p�ѣ�l���l ��pʱ'��_�2�#��.�?ǔ�I��!�#@�ae�sF�&���ԧ>�lW&.ǱZ��ot�x��������W���>A?򑏸�,P�х �s9�y��)X�<4�o�{�ڪ�ׄ{��3a4as��Äٷ���គ�c.��n����mőO��#;v��[?�ż)��p�	�Lt��� �Yy�Y�t~�@���s\j�r^4�g\s�]p�|�l9�rϚ�j��ݤ���`j�#�qM�E}*kF�mh���� �q�Z�E
�C���|��o�/���5���u���$����p����I�P��2?�ǋ���g�M]HZ�
��X�0�Xp��pұ�R"U��+3]V���@x�L�@@X}���0a����|��@D% �<#�'�g8�y�(EhgA�|<�5\�4� 9c69B�E�!�q��!�@(G�yފ���_w�ۗU����wl����+��1k�d�yͫ��[�{?�ow̱Zs�au�&��V"����F 5zaj����@f%�-˩�b���qڠ��Z�tP>+�+��a��q���Wmh��)뭴lǖ�,)@��o�ʆ�"��� 4r� �n=��Ӭ���D�u��u�glz� 5��o8��{ͤSYɒ��{�ܑ操h�>~�E���K'���U��W�(4dXb���sorӳ0����Ҁ;�rɆ�������^}�1��NOw�:�Ȕ���p�$	z-�2C��!h3f����P:�:z6@͙f�8$���P���"8� ѢP��]G���i�Lu"��!)��j�7�T���(U4bҘ���q�X��E;������4a->r��Mń���&y?�#�����4a-���M=����N�ue�9�܀#֢ȹC�~%>WʱH
 ��S�� i���p� �D��=�E�d�j�z˲���+޲y���%D��=C��W��z�k�����5�a�@�ۈF��Qd:��P��TMڏwS��u�Nۮ5��q<l�kʘ�M@ŵ�4[r��pֲ��~{��^cCu���V�R�������Z-J���A#1�%�=�Ȟ�,�)�^���a�ꈧZ�j�Zݶ���L� �g�h�ζJ��:@�v"�j[S��平&K�X�5Q	.c��}�q1MڃDwv� �C"C;�m!���dR��@N]�),g��_��~
� B�T��7�K'��hu�"#6%G��s����X��� 8�F�PH�>K��؇7��ߴ�X��D@���;�̘�Á^�<"����zO����e5�m	������3��� X�c.4�Ŧ�A����|�#ǜ@X�,
]{� ��[__gh�n�ǰ/%)��V������lN.�u����P��~�2qÅ����>��4M�7�x�[���O���C�����t 4�f�yϻ�.�������'k���e�,/nN�U7@� 4���̀&��<MT~�L���|Ql�L��W���Nȑ:[����V���?蓂���<�.��|{�S��;ئ�I�ڻ�c7L�R�<|�)\���Fq͒Z�E�~[uؓ��/{��s��w�u��~�h��v�ffx�a@T��$|��#T�M �-)����ZB�u2���\���y�P:'dܳ�е:��s��_��^/��K�!����Z����Y��X�B��sHz��bބ㑬:K�`�ra^J:�3@�^�x�����U�_h�.�M
g�B$��H�S"��o@����c �*�\��9�ƊC�6`�UeG�\IE�0E���A��_�Ӑߡ,�馛n�j�Ax�O7�Ό#GD��TQ;��g�%�t��{����;;���sS�):A+4��F6��j�@k�db<�[���T��*���H����>����B ��Ť݉�ʊ]*�w<I����nN[N	 1kY�R8S�{.�+�����Ψ��Z;K�V�əF�h�P����1E=� �uO�0���J�G.y���o���ŒP�����<��7N��~ ��|-|�\�o#��ZES.����4�	���_$:��%�%q��x���g�TVQ!��3��z��\t�ԅ�d_�H��/D551}q�N��L1S�E�EDa��3�2)e=��+W�k�cX�<#�O.T֕�E�7�����e-�^�w�����s��{�����U����֝b�^~�mߺ����d�bt;*$�����y���`�$|�< �)�H���f(z��>�1�
�g�h5J�����&���)_���l�AW~�`    IDAT�d����j������JU����b��)Oi��B�����1�Ez�I͊�d�N4ݟ����췀S����r~��&�;�ׇ��������Z~��@�쁞?_�?>+,����H����^���C e�IǗ�S@�q�����G��F-0���_j�b��f�V� �A��3��y�	��_��_v���)A�$~!�D��z�~$e*� قci^�K8���H!�'B��k���S�_�� ·�����ea��_�{��3��R� M8����	§�r����}���ǃ�)�W�It,l��A��8�b`��e����ωF���O�,2������ � (�=��P9w:�
��^Zi��%[8QO�}�<5�C�e�d�:�_�}���iR g� �׃vH�E����g��dL����u�`;b:� �{|vG�(�н�K a�L����?t��h���<�s���s��/����|����)��s5�B��W��.�[> �:�^�+�� E�=
�7rȨ%;Y��U|HDE��983'e�s����j����M%9���sN�#����i'ji!LӂT�1w�5�\�;g�yfQ�j��y�	;��~�P{fC�5ת=.GP_��5�~�Q���s�SN�`����U$��A��4
� N
'��F�q��ly�a�46���פ���~�������=��"��wz��4
����=e�I��*kC{s�����Yg��"[V[����)}0��m�`�Ԙ��n�b����� \<�����QW �>&�;&٣��r�	;_݈E��C��X�a怀Q��T�m�C�C�P�_�'s��v�ii�w��4����&���,���Y0V�b?���|���T� �H�BG� ϊ�8cpGa�r�GH�X�+"4��p���:�)�~P@x�����ҙeI���@��Ɔeնo8<��AX���(L�7�,K����1JĔ�C�`�rX����Z�ل�:�94���C������i�-d��oy�T�V��L3��)w�%X+��v �b�{^x�=�+���
zSP��3 �`,>��q�k=tt2i��7T��ھ. `>J��ޢ�K()�ό������<O����y���@X��,kS�$cO&{�a���V�I|̓Ї�9�<�$�9;[�-L����-���:\,n�Lt^x�����l->
���/JI��K ��C)�R���s�vl���t�<��O��]���eg����4М:�ZK��L����#���# �f��:�02�r��� ��G���W�)�Rv��,�.	 �zj�)�� �`�P�J@)�X��\��xY��öju׆�S�ʫP�����͢�O���J�I��;�*k(��������-��d('�&��i'C�ܩYϠ�JY:KgW�y����`0����"x0�m�k��[���~�Y�k��֣#gB�f��s�CPS"�%�N���;�$tg�q�:��clUa���w�+ic!'�AH��W_�q *�P�x�F����|� ý��k.�� ��Y`�V(�
CS vpK�=�Vj��<��������:�n�kL<7���w�(k6����^kΰ�4���*�m�i:��������H���@�@N=u�_ܯ)yL9&�]ך��\۵ȣ<`-�+O�(Aد�2��������F��)���:c`�e/!YDphq�-h\�-�/�z6քS�5��ɚ���kM�\k�I�x�n��~ޅ@b��Y~���х�ʅw��ShZ7!q?F�-T/�c���V��\Q��0T�g%��:�LXm�X�:�[ S�B1�Pn��h�\.�2,�S�V�d����"<�,�k��J��x��#��d"��)�
���kkY�������5;�nn�<9B�y1�=��|p_��lN@��Z!�٭�vj�e� u\��l:�R��_;OMݹ�N�n�u�ɱ�{�u��E�t���@��������r����5�">��н`jᙏHB	�ٚ�\��	�J9����hC��)� Kh����Gֵ�g;t�8��n�� ԭ�@�����T�� ̖��\s͛��	�����z�C���3�/Ą���k�-t�RL�C�Pj�'V�5�Ckx.��^;�����>Gy�X&\�T>{��W�� ����ڍ��U�L:��"���֥�n�^��r�C�j�C-��jEO��s���BdO�5�nv<_��:I��]{�o:�3v.����?����U��mj�\81���\�B��9���>t̡8�O�Av!@},�.�J��k���7� \*���U$���5��n��bq!yb1�8t̡8�O��Ɠ�������#� ����Aᕻ��2�:����l���2�����x\��C�j�C-���c)g.Ĥg#��ß;�r�� <��vk-!�.���5�!Mx)C�б�Z������n�Z�.�Z�Ơŀ}x�0C7I��_{�o\V9�舵;��35vA�'TMLZԂ�X3���D���d��nN�<�VP��UP�c�����	���-�U%I�|�z��}��Đ'�P\���L�ӱ9�%jf���ۻ�W�����Sx�f��y�����w�p�({��4�J;����u]�s���m�v;���<݁F/i�+����Z܇>���ؗ�Z$�����X��<%�h�������V8ǦiJ��篹�7.ktsk~pc�����6����ay�0����w	h�:;'(B�1��<��=kH���X�Ұd�i�p���� �G��8O�ε�����jd�a������S�49B���Q���I��2E��$J�����!lS��HR�}j�nֱ��:�¸P�(G�����*�	STM���+m��?�P�z�i���3�ɭ�.k��'�ND��Ͼ��|Ӳ��\�cۦ��q�AiF���3���yl5�ޥ�Q���\@W�Ȁ$����	�_����Tǆ)�4�R�<�&F����C��Ɂ0���r63.�䳁����ͬT} �0�N-c���Rjm7�	t�b��\��Z���|L����3��c�2�4�*L�Vv,��wҭ��®�WY�*��(�X5�9�td!/��|�6����иA(�!���~�0{�� <q�EY�VD���KYR����P��njS.��ԏ��7LcQ���q_�ܥ���k�K��򷵚u�
���TUb����m.���}���w��!����R��{������)�R�J8�BY��e�،,�pﱥ����X��݄�6`Nt��`57���X�Z���2a6V��v<P&���*�V���9,F��z/Q�)T$i�e�$�Q;�RQ0��ƠԢ ����UyOڳ�:[�eY�$��馛޼������9f���[�ugsa/e	�5��&\Mjv�	'y�3�+�h�Q���:p�S)e,yHm����:�i�IA �F����W\��Qb�F���O�a�}�3X~Q�	'�lZ�B�;�.!�����􋙨2�Y�a23�AX ���,Qas��i=�PLU����'��)|ń�
�<,��f-��+sB�E0lc��B�R��\����s�����t[=(�h\h�ƾ�����,p��z�v䡶�dRmH�ߜ/��a�����K.q�e)i�7�|�o-+����{��-mN"��f�3�4m{���/�~�g�����������F�K=8�9پ���x0X�W+KI��^��Wzaw�
�u��h��?��?�5!l^TB�^l��"�ʂ�	�Xf,p R45��-�P��<��� �S�Zf����*D�E�� I�~�U�:;Gk�w��$�¶�%2�(��%�} ��Rd�g�x�>v�ئ��`��!�9q�I��/��S�}˖-N� �b�c�	
�����n�+�qmI����R�禛n��e�ön�4؜��eq��5�v�e�k��ēO����η�Gn�X; ̍�TXj��P����#O�` �V&�����~�zc�e���0c���a0����9�r<�
����O�	=׽w�2Q�Ye�a��	���4������K���^ĀB=����c�'�"+�;�B@���b��H��ؖ���v�0�  aɀn���l�k(��K�K�'�`�<'8"�J�jW9� i��9��]��0hD[i�����Gb� �oj�K,�v	¿�� |�o^���M���Rl�C�ZGv�i��/�ܲvn<��x���29U�Rab�00d�*�.+<��/~�M/��<�����њ�~ɁƋ�n�wgl7�=��-e��e-N�(*�jgb��ahW/�ζ�8���Ga䅊sk[�wo�7��"�p_1���bcQ�����W���Q�Z�F�� ����9�m�v3"iv2��eIKܩX?_�I��g�1t�! L��"�0��7�W��fN!��ga�Ȭ ����Q�I[�I��֡���6\��5{�o���k1��"a�C;�l`�!��De�7��,���� �]t�c��,���.�j�	8H��l��?��[c��ҡ�<o�q|��7�������9/� y>��ڵ��K_�[�z����?��[������&+�#�ѓ���D������V/�3Iit��Fg�O9���/������c����ڹ�^���l7,Kؠ(�8�,ɫS'9N,�k�N�V��_�E��/F��,�V��hP��;)�^l���Y��>�������J�e��[�1ױѴ�Z���zll�iQ��r�FjOY���le688�+8���B�Q&S���;��X� �U̖��3������|��*}�]R�F��u�O9>�n��\�(��Śb5�0��{-{��?V��BKAE�`xX~�0m.F�lS�������}!?	�ɑ��o 5��O�=�k�����~�U<����E�����pa]*s.;���u�s��8������}C����|�+�|����d�&�gc4 T_�9�[q��
sN>�dg����q=��q��c��o�j�A��m��	;W��k��֝e�{��ܽ���~���*6�,�]���[f+���I�1!Y��h�dx(�>�����4 �\���x�w��M��{��^�A 4�Y8:"��͞�YO�~B�z6�h�������f��a��Z�����e6lY�kI\3��i�a�5��a�Yb�%Va�O���l�;.ge�b����Gj'��am�f�eyϰ�6sKz��m��3V�V��L-����me�ϵ�a�X��ڛ�u���y��Ō$7	D���x�ٖ��arL46�\�������w�f��ª�������Ҕ!&��K.�ĉ�fѣ?'�����I���/�r�s.s�c�$,��ER���/Ӿ[c^�G[0v���7� �@���`�� ��	�8�GO�,#k�~9W�5I"�"��M�[`�ӱC�g?�Y�GinEQԊ�x�7���SO=ud����6��8��<�ЦYk{��f`�����?m��v�~Ӧ'g|�L^�'l�':�	��ɁHs�I'������}��a�	X���Vt�� bP�����X��Ă�[y�jQ��<��x��8q�L:I(l�Z֞�a��ڶ�/����G�bGyӲxڢ�U���ȗ��;9�EHiɄ�J�;�K�]�YT+wp�,NSk�UK����F4dI��%�j��Q{�I��'��| �PA�.E�ȡ!�L:$MS�R%�cذa�O\,��ǒ�<�����k��a�/"�"�gԜa�/�C&.��s�)M�A��4a���:�|ļ��gø�a��Q����a�.spbΪ��	�L 9N}"�N?�tw�}���������5�\�D?c�FB��� �Cb�8�5H m#�!��̡{�<�c�����]�& |�5׼���~��e�y�sS�3����f�x��m�5f߸�߭VA̮�ꊼ�nv�VEn�P2�:O��@`�������?��yq ��
�x=�Cg3�B��x���0{�r׮7�*���XiIT)w��,�&�'��<֞s�����tݢ�bI��X\mZ�'���w�d�	}cP�� �Q,X9{����\��l��&����V����rа�9�k�������oج�Y� Xd,�tJ@�6�G�,Ą������A{k��<y�e"��_�җ<tJ`�6 �r�).p�o~��@g�}�?; Ä5��k@�� uM�����jC9 ��cN��\r�ƽ��Z �|G�N��W��Ua2��|��׿��w�
�q��	'�`�_~yg�^���9���'�"�n���e�6����9����	(�T;��L𓍇_��W��iG�{L��5��`�sЀ5Ƙ[�c�e��������V�Z�Ե�^�{�
�a�p�^q>�����Ͽ��z��y��=c��o��v\�E�C�����n'��X��:�,w�}�_p@�e aJ��c�a�p [@����$Q�\�.�b�f��Ȧ�Ik�T���m��
���X%���l������c�lz�NK'
�7A��,�iY�`Ū�Ŷ���<~�[�ю����۶�ڝc҈ݛ娋͢�5�A�6�o���-�eo͒��f�8lV3��C���x~&m*�!dG�i���g�s�1�MXk)�MLv �2�9�Iʀ���w0Pq��9��#�}^���o�������	�L�߹��s~@X���Ó�1��&���#X��� E�m�{X�|�V�d9���-&�pB���SR	�ym�� 2t LX�ĵ�8�3�]v�[ь�?��?��(9N>(�	��/~�k��E�v΃ �lն�Ap��6�m�G`Hj��ԧlb���J��'�s��o_V9^�{Ǧ���s�� c���^l�}�y����۶<�S�Z���+��C�0aq ����!�����eT�kݺu��7���$�$���4 �Xߩ pX��l²Jd�z�=�����ZOo��m�Ѵ�c�p�����Ǝ�Vi�]�h5'-%���e}+�ĖEm�-�=��� ��P�x� a�$��u�2��5sL�Ul:^a3=O����f��Y;^m֬����Ծ�w_qYFN-|b�1a&&�����ĵCY)���B��cp"-�ޘ��������W��c]ˮ�5���������7��#cx� ,тL���1��$'�m��r�s�m�	�9b�!�s>}���w+����˄�L��/���}z��9c��b���+�饗:s_�YI�	$M���h���cq��8H#��c�>>�<o�qr����o۰aÞ�X[���>y��G64��E&*��u���_d���o�O~��U��E�1�r��蚼2_���,ei|��4�-���%F������J�ַ��l���R#�CL�*+W|��
p-�Y�ֶ,�,�*����v�ŗ���g-��m0�a���,�u�ٞ]MU,��Fl�hOZ�3c����-�"l� ��ٝ� a�+�S�*�-ɩ��g�����E=6��ht����Y���hX-��*�c�6����_g���X�&�b�0Z;�-�`��F�H�?�2���!ib��hh�qMm)�?�'V�&�R���X��Zlh'_����Br����Tp b.(K�$�D�Lr_h)Ѿ�'��C�"�\���C��9�(��a��ǜ��"�@�`�,��]���Iý �<�^��Q�;�ڗş�Xg�{���CF�P��p�m߹C�ҵ�(���k������]Kc��ʇ�l^i�s	�":��O����W�w���>K[ W⃆���$E�<�< Ecȁ�g���̅�i0���I�~�s��f��s_:�L	9����5
 ��v �����s
�)���9b��N�O�g���X2�ǲ1<f�j�5�զ�oUb����q�2L��H���V8�J�!�'{��t�&z�x�{l��j���#,<����md���zWZ�ƶm�öi�-�Js��2���N�ðhO��2@��(�+�n��̄�[̈́T�<��O}JP��d���?}�R@�c�J�pѓ����R�,�қ5OȒ��EVćc`��0����&/?O� }�3oC�l    IDAT|�j�p��a���_��_qf/�<c0&�a�������>5�Y�9+�Ϲ9�p>bi�=��},�x�y�Ґ,­۷�5�$i%�ʧ����߾�䓗�	�����գ[nퟙ<��nX_������Wٖ����A��乯PԐ�a���D&l�N�� ^:�ق�K���t:�@��y0)^���q���| �55�+�eI�</��9�γ�/�Ģ���̢�n��X��n����{���VV��U��5,�N��a5��Z֎�;��!I�j�p�� �e���{F�<�i"��L���DGZ:t�eC�ۤYd5��j;vm��}�c>xh7M"9xfs̩M�,&#�KE1����4�n��IqL(h҇�-�&� +[I�|6'�OZ�9�&r��������=�dԢ���#�����R����ʜV"�/�*�G��:�#s&�~+*�>Ww{� �w�Gڡ|:��=��7֏�p�6�关��q� �w������cz3DNl��E/z�;���	<P;s/$v�`c��"cY�q�ߐF�S�Y>g����_�ӟ��M�L�m�I�r����v�o����G��:�Μ�8�U}+�5�y��+���g�j4Z�P�xb�$�j���x0Y���á�`��������x�
N�����c�G3ؔ%#`�SsLK3��YVi9�ҺmX��.��R�)�Jjq{��{,�����Z6�����*�%V�v:cV���ê�ͨQ������ a_�<��@���C����fU��W�Ht����[{�6c��y�؎];PX,�����^����!:�1x?X �-������\d!���A,	-��_AցE�,��O A��<���m�8�o �v��x���с������~�/H z@�����':��G���x���G?��Ge�2��_���:I@� 7�����d	@�R�3�����I!�$�3Y��8N6�|�o]�d@xŎ��4��#�VWM{���8�t��o����5� ,�S���LQ�w��*i�����/ o�V8��I"a �)���/t3X�k� 7��!��{��k�P���t'-���ε�/��(Z�T2��^�w[4z��'�u&� �V���X;�*@xM͢����aq5�v	��Q�`����펼*���DByP�ØV���Z��K�i����Q�,J|�	�s�T�ik@�I:��B5���̈́+z�@�����2�q�2a`8|��$�[lsR����
��b�k�qA*��s ��b�1�áDԊ<�rl��cɄCfͽu3aƗ�Z�Ҧ��7��1�7n��G;]u�U��}���Xrh ���'���'|&'��QV���NEf���yqέ��Z�ǝ]N�8�6���w^��������j��;o�=�R�#�Fn�x����r��{k��ۿc{��u�T��<�FiHҠ��cN|�;���d^�9A#6��/��l����'��AJ�22�^ �=�q��(`^;����n�;�.-A8F1Ha»-�{��L�rĄYҮX-��c�%�yâZD?��@�9Ⱥ�� �Y+�!�c.+�
��ؒw�5�NV�H�p6�D�]{v;v��qhƲ�	�	��e�jA{����-
c��o��+�`EL�4j�έ��q  YʄY걡�p+�S�E���X�򗐀�sa��_���X�ɯ盭m�N?/9B�7�q� �u�n��O���6,�$0��?�tX+�p�X����q��״��44?���tb�C_@���/��R�7iǟ���w��noodsc�<@���e�{7<�l���n����L1xJ�`Ő�%�=7Xw�q^ד�)�ê"ݏ��Ӈ?�Y�t�M�'�h�l�'g _��>�B�T�%B��l(����S�f�����B��jn��a�#��,۽���أ#`�E%Nz� Ѱ
L8M]�)4�"Y�x�Cj0����d�I9��������׃ӡg�4 l5��9��>�яt������t>��оfa�c�	˯�s�Q��I$����d�md<���BR	��c	�|� J���XwH�[�O?��uc*S����Eb���ǚ	�ϸ�L������w�	kH�j�P��i+B\�z/�g�+	��"��t/�"p�9VQ"�M�0�JQRT9�r��]{���}��q��y���Q���P�jN3���U���/�c��ۻw�'+��t`~j��0����d��<���48C� F������Tx	�F�����A<���`Z��c��#�~~5�ن��y(�9@8j�#��{��=�-3���,A����6c+V�XқZ�Z�	�{Z2�C�ps����,f�T�פ��4�Y#^i{��>��Ԧ��1%�k�}���T�͹Js1a@9��	?� ̽�AĠ'.���������cG�C��c`���`�9�T��}|��G�3�I8�]8� a�5!�<�����_�LD%�������!��� bƳkLз|/Y� #sN�j�n k�L�B!���q"|�aI�\�q���u�D��Dj���y�F�����~k�Ax՞�n�Z�o�Y�*_�o�y��G�e�\nO}��;&<������(�a�_q�����XB�-��D�������;5�u�D�|�΄��S��>�U�2�(����b� �ǹE0�ֈ�,Ax`�f��[2n�kWc���ZeƆ��&��N����v�.�o=羞�QTS#"���URSw	WJM�hOk�LM��Շ>��t�9��҄CGR8�5��ßgt����,�)�i�L�C,1$
�0�1@VĠ���9� 	�Ysį��x.2�p��_p����/�Y]�7>X�9�[��$k��m�I{i�S,�p�=�UD6�X�)�X�)�_�D�(� ���H��e�b���gL%I�믿�ͧ�vZ�f��W.B���?3���6��!k����#���ϿЫ�T�&	Ńk�X�y`�[<�8�4�@�QQvV:�A�7�/`��8��C�r����}��sˑ����9b�q�!e0W�#.��b7�Jdyk�V$;�2r��>`�.�plQV�V%����:m+�L�A&L�Kg�D�)mY@[�����F%6�䊈	��	Q��m$:ڲAs'�t6XD]X�Μ}�`�s9$�c�b����v�-Ą�cN��B��h�D_�rR�����B�L=͇n=u!Ki��h���}bZ�З��u2��C�gZ$�Gat�Ƶȅ���d�z���&|�SV��WI�q��9a���r��>�`҄2L� Ua�*����5�/�o��^K�\ߛ$��������SNپ�q� ÄZS�Z�EloT�F���N��Xjδl��՝���Nx34�J#�aa-���.�ք'U�X��Z�X͘��A�j*�.!}�L8�T-w/<�#S�p�:���+<�"�T��{lE���?���,ߵ�*�5/{�&�5r�iZ�cվ��6eq�>w��Җ�+�sA��je��q\��OY��cʆlĞb6|���������d������G?�1DZ�d��jr�=4i�R���sK�q:<<f���Xf�&�)m��	� e*�1�m�p�R3��g�1ǘ����l8)�pqYʄY�cgc�ZS��-+�]�q��r̅���sR>�;��?m���e�"�[9k�gQ�V���\EbѶS�1�P{�f��o�qE��0[,&$Q�^�B �(�`�~`A��$�Y��9�ƊA��P�?n�⁤�J4g���r6h@i i ���x脜�/%L$��#�4�(���iIԴ���%�\ayT�(�ytĊ������F�|�KƫV�H�Ȭ�p�C�*}��(�S�"G[^��K[�E�(k\�#��&Q$8Sʒz*�3���3,>�Z}'8[Y�~ddrY@�I���c�Q�θO0 ���zʹ�@�u�j�Q	a�j�j�9M�p⨏%K�\_s,�� ����{����\�x�ɿ\�/'��_��x
�R���n܇�Q���e���A���b�b�ݖ ��/�
#���f9ڰ���-�p��И�Y��H��2�3����2���~�-��/��/����u�-���	�\c�2�wZI�h�������Ԑ���JիÀT!l��,J�Q�7��}V�����l�����c@���V&�,��c�}�l�N�Ɖ����0��,A�m�h�ab�Ҕyw��>\�1��uΫ�!�"��|���3,[>ѦmЬҶ<�ld�1a&��61dEcU�"\h{+����<�ؔ���K�FAh:s]9ESE�/���1�!�-3�X�/��J�S,5��D���̧��a�@�9����zDu&�8�� _��cT֡p!|v���/��4~��y�RP}�ꫯ~���)���d����<�4�pjUY�����%J�����>���2�H9v� lYW-&D-�a�L���"D-�A��ȧ-�4l�0�p� Wr��,�Ȏ+�E˨A�����Sт���F�ϩ���^{�e+N�f߉6� �~��ޑ�b¬����M�y'����j cn�?Ŵ���9� �|���2���=F�_�R�Z��.�*G�sD ��e��|�X��
L����+��\[	�}��jĜ�[���	/�8�!�MC��M��h,�3�|�mY�a�yI��tssi�����v����F�đ�NTCΦ	k%�3��.�@���>$I�˄�j�~h"9� �K/�ܓ!�J��ֈ��wX4r������[gUK) ��XTi� L�ܴ���R@�eׅzV�q&iCr��QA�cW\`�$ =Ͳ�S����0���yj���oM&�IF�$t2���>X�ژ��!kcV�_&��JJç_ m�C%� F�T(1i��g��Q�D���	/��1�YHHr^��#Nrڗ>�?#�x����A����1"���>d���"�K�-/dg;&���tȴ�H�� �CK�G�<z-(:����&_z�;����g���W"��	��6�&�Tc���� �!�sp���39��%GT]�hg0��ˊ�JdI9b�%#�Z������'2KҚeq�Y�� �#T�_���˗6��w6�$�W�k�gЩ��d���FO�lų��m� �,�ѽ{��f���^�2�F�T{j�G���)9�|E�p����`�&6!�h� �����7�^�0a?���>Iԑ�|���x�\�+���0a�@E�f tZ�	i�(���8"p��
�|���x��F��6n�ܦϥ�ӧH�:Sd��R���$-��]J_���l�fr�"fb�]-�"�)ZV[qLX$ܢMU0���f�{m�j?�Q��kU	�y��р�*�P�;�,11�Q���B :"�+%gv��뼞0�I%�>+���z��l�6�ɖUҊ��m�M�jᘫ�1iqMv[TM+��[��Ow�#.�Kf�;YSLq�&�a�c,_y������h��fY��Q@���̈́e�2Y����U���r�i��M�|���5�b�3i�Ì�WIH Oz��)r  `X8p�!�(*JYv;�y��(�N��@����!X`�B`����I�� QO�0���F3>�Ѩ���o�)���`GG,��"',V�~�n��cDFĞ�\Z��`�>�/_}�տ�sg��u5��թ[��i���!u�:�������D���`��SO��CmR�G�����.����]���c[,ݽ�l��!jq^5j-��=V#m9���kl Zh�*a��j�o���L�D̡^���m��\0e���h�'Z��X���Q�3��>����4X%�҃Bט�r|Jv�x&.Z;(8^+�ˎXv�Ez�yU��3R���1�n���:Ąa�%bQdn E��`� ���N�d�J^�| Y���IW�{J�R�������S���g���.�Wu;5�ĈC|���*`�v�q^����C��F�`�c���}q�u�V��&�LZ�S����aM g�e�p]S��YAè�j���|v ���m|z�*=��f�%qfg�;�֟��B���6PkXOk���wZ��Vk�|��vj=l5?M��*=��V�ޟ[�PԽ�l7.����
�}#ϝ+I�>���~��UkE+m�~���Zk՟b�jeв��G?���zM��[�_��~�U\���M:Ҡ�6���H�..���Ċò��$�����������c.�ﰟ�]
�׸�<~��)r!F�x�<dRr|jQ�I;�a����J7�}��-����B������=Q1�$%-���{~�%�cMDI�����g�kt��>�YdOq3ܛ�l�w�Eڂ�BB�=��Ӓ��x�oX�d���4Ԟq���nMb���g�S@��0Uוϙ�ܸ�e���A\#��al����X�a����^22'.��g�L����f$��@�������ZW�hU��b��"�!�	�[���ZwHXk�U�j���T��ֺ#n,!�(��v��������͏;s���0A�>�<�ν����y��|��}�{�ѓ�jé6<���+͟�gޞW���J�f�ғ?2�������4t�})�R����fͭ��Y�)U�2���Ŏ��O��;͍.a.�p��G�s�A�[ޏTSo�i`d��뻺ӷ~�5���z�>4+oo�?0��fW�wݞ��pΧn�b�A����ٌ�Dd��@ϧ�R����ar �5�/R>s@ǙT�d��B:K�C����&N��O�y�:���s1�`��1�J�@X������0�H��m� `��;֔���˾k�5LG]���0<�L<rue�jo
ޭ�8+�3 �A9�� |�����-����h���8k�O�B5�.� ��wDo
���W�s�_5�5���R�|�Bc5>!����T��I��q@`7�����Cs����ݝ���Ҳ�H�<|ߔ�ߛ��G<YB�!
����9]����b1Fa T�h��l�+q��k:X�\�J��4R�3m������Mw����4�wn���<��I�Q�� ����YC9n2�e����HhG���mTpqq�!m�̲��g2cLؕN���;qO����xV�F�q5�u,�8(f[��j��X����`A�v�(Q�6����x�5�hg�qħRg���{%�8��?JأP�K��w�H'���1w����Q&��'�y3�ޡ	+�\\P�a�N/bt�9�����gܪ�q����1A8�Sȫt��z-k��*}i�V�	�{�7�=u�t�K�z��<�r��Й�׺rv}v���~�#�d�����0[�0.rDd�ݨî��H��oY�(r���M��J��3+�5��`eϼ�ܬ��42ܕzq*��	��;��ul;D`G������y���'׍S:�����ц�e9��x�x?l�)5�F�|����e;D�}�m�q��� %��I�siyd��c�D;����+��}G ��y����Ĉ�v�s��&��vm��x���0ʛ�m0JL>�q���:����3����4ox�ɀ0�0;k�	Ä��p�O;�y���J��p1���r�Ƒ�ϲ G%��wݑۥ�+˶L� ~��s�B��,Fm���C�eO�>�����Z���	*Sw_ޝch�Z=/ި�i��)'ú&\�z�����	�yϏTEbIi`h0�V� y,�����ޑ�T�w��=�RmhG�&�N=�p��:C��� ,��ь�6|Ɏ�%�C���dJ���#(	XN!a�q#˩v��:_)I���"HH$�t:j�x#��b�`Tn�g@��8˱�c[ęQ��9�_���t�o�{�A][�;,'��4ͥr���qF�����ׯ?���,:�m݂&��2תEn�rr ��I��ȍ��J�NI�C�C��	�����F�GϽz�w�0�#�E��0�X�Z-��HwW��3�D���ONVv�����W��9�C��v�V�'��x+���H�N��ùJ��m    IDAT�r�E<p��Q�w�``뮧
@?RO}LS=�{G�}��4������ԗ�#�4<8��K}�l4�8��٥��LB���k�Q�ߨ;�3؟�E��i���kp�ZN�}6ʍ�ow��S5`m[���R81,�6�2M���(�U������	�n�1��o,�1�Y�`�-r�a�ܡ�R�Xvن<�P4%1��` g{5�0�I��� �c �V�����	FA���W�[����a��{��-7]6���ı@�o�G�$��RHC������O������
�����n�ǘ{�D�q�T5=�c�
��@h �f�uో\�Y�������Z����,��\�I�������`���2-'>���`��]����袌"�ew���ݬLN�Yը���]i�p�W�){�9���T�	�y9��3E�����4_s��؉4���O4����S:�:8���I|ﾲAX��Fg4�Eu�������v1����m�]��x Xx%)�7�x�V�C���f�Q��Ⱥc�&[�c1me�Y6:g�D��O����a N�û��㽭�Z�FR�O�]����not�)o|̂[}ټၣ��#�,MG�<O{`�,�t)0@L�#��,����H����F� ك�կ~uf�9²��_�%}����F�lC��:t\l0�����@�DO7aa���RO_5m��K�>��ޮB��W
�2�YlW^��f��sNI9�0����bۣ"�;�,3Lf�gw�kp�t���*��ix`8�)���]��h��3Ə�k QFh�c�'W�;DD�O��9U�N�DԣǺo�X˯3���d��8/- ���h)A"z�%b���l���9^�ԁz,`�H}4c�9?ړ��l��J�2�";��C`x�@\߈+���X2L���$�'F]���稍�GA�̎���3�}�­7_6����f���������@魥�G��z���ܹ{��}�ĎJ�!���cB� 8a���I@dtTSw�[������8 ����,6d�Ҙ��[��e 娅��JA���ʷ��b��w(ݦ ���FW�!d�P���G&��.'|gq�+��n�1�sfj`���8#V��oH��t�Ȍ�-��/�F8P�q�gnԈ� �0Y��y����q222R�V�W�^����������qo��eF�����>�ꛛ����%��}.�g�����<3Z ��;zEu鄃�`h2 7	?H�c�Q�6��F$������Pl�Ɉ��h��2��t|���f6S������j@)�߉�!18@�~&���0�S��3���v�Q��0��7�*gI�3GI$��N�Wv�t�pT��U��O�Y��� |���{���n�t�T[>8ԟ*�=iN����כ�?���'<6���?L7�pS~xG&
�X�W��2��T�ёyg��I�u��(lEr�gf����hv��yի^�+��@�0vT<��L�����=k �����/��>�����ӟ�tƒ�N;-�ڏ}�c�8i��'P�p�	YZ��%��o����p���*P�o�t_&<��U*��֬Y���2a@x��o�t��m˙2�T����ZZ�|Yz����n�rC����#�2Y�:#�9�@N [�8!��lO�6��xE��9�5�C�1B>�y��K:/���V��{�}��5S�����V5 ��߮]�6˖��H(Dn����gdݖ���o�L\b��g>��!���Ȑ�W�z��椁�q-�y3 PwvF�X�j���޹��9��d�	���+_yR���M_��������<t�=��fu9�0�0
�;R@�'��e:�ta� ����f$#/8�{���8H��V=��L����Y�k�o�ƍ9���?������s�T�d��ߌp@�$�j�9���~��8j���c�0��Db!��?��$����3�Wz���z}���s�ʋ.:�裏�c"�9��Fh���vå��+�g����:��?O��vk���'��0� -q�)����lt_""m[��]ՠ��b�w[#7�|]2��f�੠�,6.��d��D*v�ؙ����� }��~�Yge�ǌ�+_�J��t�Iy{�ؗ�����~p�햸; �n�`~#���J S@��	�u$�Fd�w�'�
}�=ц��ow1�p��犕o��G�a^t+ <�"�k�w�#Z�^�����~�����s�c3� � �a6�y�o��%nh��~�s�˕�s���>7ꄓ2�u�ע!�hB��͵�1�i�0s������	�N=���p�%�4��������H� "���,�e��A3k�M+k"}�S�p�br� �W\qE�>�ឞ��^|�9aC�fo�gEo_5uwU�҃O/|����?��t�/�z�}�
�ٳ�l�~�2@�QG����k�"F/�7�q%
�d���'���m�љy��)���vr/�s��㙹�L����k��f��0�8q�� ��_�H ]�3��
p� +�~�QGe�fd�=@��dʞK@ 8�}�o����+�+֯[wnGW̱Xc��o�l������R�қ���)�9�yv���+;���B~ (M�e��Z����<������+���Y��-�tR��Db�Y0�py'ͭ����L�&w��؀+4[�4�+O�r �剋����&w���fj`�5�bR'���$�����~&h��)�a�G� 4Y��~����Z��֍�pI7�s�x��g~��[2^�j���+6���Yf��n�l~}��=��'�bɲt�q�������0�,a m�/�1!F�&L��f5���e�\�E�`ʡW�� Yco���Lu�Nfq��IE�+��d���yqE���������@���g����]Q�#��������P15Z�hq��C� +�lGb{��h����a���+s_��/��8�8�.�i�;�w�i��V*�׬^s^g�#N;瀇ܺu��{�Ȋ���i�cN'��������?�M{Ι�����a��v|+���n�v������O~2��6c�,��F$e�mres'�s��
�h���I���,Nڽ�T����u�KY16�nq��<�{Ϝ;SS���J,0��MDF�Y��=&�r��/� 4�4\���0�p�o�;���D]�w�e��&������^A�V�t_�f՚s:
¤�|ح[7Ww�Є�ki���N:���Gw��7�=�Tzs�'t���&Y�s#���k|!�Þ��?�3�ۿ�[�B ��s��:(k8� F�1`׀.e� e�;�	�G��Bx>���j��:�����['N��aДGО�#vU��\�� ��^t�EY����?�#�d����?���o0�Q b��׾6�� ��nr�{��9���H$Տ�vf��)��ȘE��QЮuww]�~��7tT&����o��{��O�ф�Y��c��yp����t�w���"��K��� OY+� A��d��J�2�&¡�4�!`�nXhs�4䪫�ʂ��J���54f hW��PN��N��v���� >S�������������vjv�]Y0^�[VŲ�����l�1c�g�}v�	�����Fg�`;��&�� ��A	��s b���I�93(�b�.�Q��bnÆgw4�;�Ϳ��s��S�v�sC���_�����$n^�|���
Q(u�Ȯ���p<������ׄ�?�ъQ��/̕�bt^� �ד��f�\	CÙpyW3�VH���it��1���u&�{̲�5�z�_��;`\^54�	O��g��d�G 
o�۳�K�6������R�>��<�Ɩe�XDz��$n �a����q�]�'�;,��C̈́�%��G��q���wt{�%����o�_�JN-�F�J�?���)G�'�����~�n�qK�XP��S��0.� ��̱_#�3� \��9DE�(X�3�1�?'��	9do�����a��"G��-o,�I�mv���D��`���@t�KYC��e���L�`�Vlذ!K���Ӻ�;F��ۿ���س)���! ( 6�G��G紤���lj�#G
������>s����y��כ�=�,jh��g�K۶ݗ�~��t�I/O{�~��~��F!e�N	F�_�# ��K:K����_�r��-�y�a�/x�r���5k�Ne��LN<��� �o�FFD0�.ӦL�>��g���ەe�i�d�Tˍ ����͙����Uf��n(��L]���`R&'��7~��,`��'V�� 1��b�[臨�p.�{ Q��#����(�����ի�\�b��v����]�����7e9��-��3��N��f��K�����G�I}�~���0��.tH�V�e)!���qn�"�������z0Ss
��%q�X 6���#x�r:$y~�ɑ�ӌ�q0������kT��1F�-����5���
����=^Wϲﭞo"���xl9,��R��~��(�Y�гo䑳��F���{�R �v1f<ΞʳJ�#H��m�M"��%쬁4qd�da��^�)���8��� *)FGv�Z�z�ʕ� ��nټ��}�u�����#��?-YrDη�*5m5��Ί
�~K�(}�m7�V��^���F�wݷ��T������Z���t�TA�rǎZ�.Q'�Af���!vJG�<��&�',؄�+!ŭ���k��xJ����ࢮ6è[[����8��Ȩ_��ٞv����a�!�dL��nx�mI��6NV�QB�OJ�F�����$���	[X� ��.���?���!��f�h�h��F��.ᅷlټ���c���]��7¦��4��������ex yHqTعy�^m�(�Ȥb��=���P1�Л�q�2Io�6IT6��ow0���pd�J�*x���A�E0��z.l��L�S��1F��-��'	S:;*���L$�re3Ze�����|Yg?��>��ːe_q`��9 ��Vl�����,��
�'���q�v�ߝ��g��]�������h6�C��|����E��o��	Q[x�-���C*���Hv�U*�y{��jW�>��R��E?!�������Kv+iTP��9��ў�q�^+�����Kc廨�L��L�}��F�)�O��m_|n;��c,c�0{����k�S+CZ�aꋲ.�tNɇ6a��3Jmۖ���3r��V'����2U�Ҏ_f��]<�w#����A�ߔ�l/�]�����S��о֭����)H&�G��ܡ3�BWRg{Q�Q��l>�jժ3:�	��޼i�4�CԈ���P��+�y�{k�l���
��x��70�w
^��G�|���]��q^�{E��4��=;�Qv�^\�5c�.q�ȭC�7"�����ĥ�tv��#�N�G:A�rQkC�f���#{��Ap:۾�{��r�38I����?���U�5/�}N-Y�ٶ�ɸ��rRԊ��(��ygJ�_�g��c�?S�֫�R��D2��,�D$���J��yΎ��[6�ڞ�p��I�ၴ=��k��OIc�Ԝ�8*;hQ�N�Ai�\S/��0��זEG`�#�*ǎ�N�@�B.�� �p3:��Og�dY�I&�(�jL��п�y������~G��҉��`��N�M�{J:t�Z��$5��Q7XW��������՚�f5�2�*)	��a����˱�M��Hg�;�	��y�������@x��n!w�15�UO��	���L8�q����O�n��4����5Em3o��:�h���ָ��8�
�ց�6�8pJ���{ �a��>��G��� ��.f�����	�'L ��� z���Q����v�{�ʜ�҇�oY�ˀ mI�	��� Sf�T�s��>��������Y�ǎ\�GR�wfBq�Jh)�%�ҁywg0�팜:�e�\g�b�����,������R���U�N�a�ڞ�ێ��Ɏ9�-��	�h��6,&��,I#��� !�Ƒ:N)��N:�1�?Fi����S��`t*HG"� ̋�ynS|�8�!lQ9��Y6��g=+k��I%�&uFAX=��pʱ��N$�)��κ0�[��e�W2 J���?=�����G�đJh&Z%[��,D`�5�g�����Z��c���S��T��0��ݩ#R�������X��uhc���|NyIሳJIbw�g�$1���sٯ��R������Z�~n�ʕ���7�ߐ#p�EM�|�lo4�+�k��>t�si�udgN�v�!��=Ǻ� [�3Q$n���;K��q�-��]�/����A\ո(&L�PLØ�u �h�>#I���eS�9"o�z�U�]7��8c�{�'rvz���������%3b��SN������75�K�_���e��o~s[^d#�"	�7� 6��~X��C�^p���X*�c�2��h��I'�@rg��g<�`Vf���vlD"!��>�6���[��OG��U0�@�ddƞ�3�,����V�^=} �(:�*v�8-K�h�3���\�� 0�����j����@
`	[24�����v��rm3�3	�x)FX��&d��> �&�S�k�0a�2jSiߩ���p~��|֡e��$a�h��?;ǰ��$A9L�A�#�Hc� [����`�.�k�\���xΣ=a��S�^�}h{ڗ�|�0�^�r�=ǐ��킢��l�ϱQ,��V}��~����ҁA����l6bV�Si�f��e����իW�:mL��
��-m���:[�L8���P��u���a�9�IX���z0 ������d(LU�6�9:*�ҹC;q䍨r�B�AnP^���7\[�w=�s�<e��� S��v����ߣגf�J��A� I�=�i���h����m~Е9����r-]~�3�%�����n�àMx"�Jy�=8�<����L���9���� 2�2�;x5g�o����,"�h�e�Fn�Kwww�A8�	�~��yC�O6:b,9����� qA�U#8����\!��P�*6B+&���Q^�̹���	�+�|yǠ	�1 c��YB�Ш�{����q a�q�kP�g̯@�W]	�DD����Sov���:�6�kE���I=�qw���EG��Xe���}۔��3 /�~�����3�5ϋ���V��
�9β웂0ύ�20�~?Q�PD[�n� �#����s<�Y�/�p3v@��rI�m�i���O���'�v�~q����oy ���*�,NכU\������@/w�����l��tZ-/?�n���~�ba6����Ɂ�@�5�N���AE9�c����܁t��=\�)@������O[I��TR��xw� �m���$�h�q���b���؆�q���oAK-U�Zߋ�t�ǁA��;�C��bߚ.K��-Gr6D��3;�)Y��r��>��������_|�i΢v����qæy��O���}F�q��fc5c�>���]��@��)_�ȷ*�n��ǁ��bGta�L��b4�XSFt?e@�Fa���D��q�n>˰"s��щ��g;gy���;�d������:���d�N�e�����`���]�F=��D�1��vv�qê<��8+⻸�7��LT0���#���a����P�Ѫ��V<>2kYh�-b��e��s�7�'~�Z�Hi�	��&|�ƍO�hRw6�\��f����@��M.�"D��м�HV���)T��+O#�M��݊I�j��{3@m��~�!�r5�������}���L�-�h�YM����0��b�ttbK��[Z�N�k��5T�G�=ֽ�S
�D@�H;�>�0m�2X�����]��\�/PF����w�j�\י�������ϙ��Ug0�%�����=Nn�k    IDAT�˃4��Y��"�Ł���@O=(��V��2�6�y�#&�Z�8j�J{�E$�M@x�T�6l8�� ���s�ϖ-�������Ã�T��Ô AB��s��E��e�cQ}��Z� ���S�����"��G��x�؋����	s0ؘ��%�t^�&E=��3�Y����&�-���=��*I����M�������E0�Q3L����zR���U�V�߸�	��d�q���UG�{��j��G�$c4���pu`y/��t�U@�r�dAXP4N�ε]`�w���l�W�tf�5�_�ڙE���c�g� Bd��PgQV��������������s���?��-�����"�����ܞ=ROO5�n���7�7!G,\�o"'3��놝�)5H2e2��a���9u4�3��!5 8�xVxq/��˼;��G��`�>\d���
�W����FA"{�f�jO��k45�hxh��>u�P��������G�Y�L�����APo0Z��9c���(/�e�갲R�h���9�&S�>���;�G�)�DBP�=p�	^���:�̤�}�M#A��z��.3β�j{�g���@}�x�xԩ9���I��a��=���l�H*��%: Z�>��o;]s�5��2(��� B�����3��DT8�44���^,V©N��"���y�Z�>
�gv�;���������I�#��R��''�a�2��k#�i����'=�������
��蘌^T&�H��*/=�N��n�R��SO͙�	��J��\���.��q=;�#����jw�N���-�>RhIN�uVݷ� AxpT
�1ֆ��p����k��f�ޣu@i���Z�:.ue�.��Da��brωr��Q��q��q��u1­�b�AX-���]���h�/�}��
^��"(:+��	�Ԗ������@��B����#N��lZ���S�X'�����@�5V�Z��г��5�yM^<"	S�i��#yP���0K��4��[���wY��XZ��KRJ$�v���C�$�[B������n�|����f�\��g�s�q�\Cs�[jw�"4����?�fAt���gW<iߘvqϬE&��<��('��Â4���"B�Y��#o�02Ȕ|.='�(��]5�I��J��n�E+Р�˿� �IK	E����!E���s]ų\�&�}Gu��q��|W�6��a���;��&�Wgk���=��C��S�B2����燫�U��+���t���SdZV`�l�O�}���$E;߯�SA�A!�gGi���f^��G�AEY]B�8���w�Z����6���;V���@����pҧ��ȭE=Iۍ��;d�1���	\�E
o������.��]_��ɾT���᯻x^��ԽO��@�1��<�n�����xĥ�D��k�ߴ6+���,���@�a�8��7�4Qf[��|~x�J�2���e �4�g��ѩ�]g[Z����K܅��C�A��W���'[�� \e��@��G��r?Ti��~�D�;[�ǆ�|�̻��	�!�L��m<���P,�ǈt⺪u�_t�D|�d�>���[M���@g`;�/U�:���6�zs������z�r#K���cq(���`p5jG[�
HJTS����b�z�$%��-4��6t��J�������#�m���
������B��5�C!��A���2-D�V	��/��߯q�0Wo7*"����?r�oi|��x0l�����v+g����gd�0�E5.�(�U�Y��6A�z���卣��pBq�[�eF4Q�Kv[Un�D8�;T �����,�X Ti!�#HZ�&,�K�<�u0J"���K�� c�v�!����y��!E��W�m��|5mA�𝌸Z]}ʺ*1~b Q��	�Sv�]�F%�Ҩ4���/�q ��R�8
��Al�M�#�7a���0�Ã�ɑ�>�+~���~�0�����������9���i�<dF|�)c��R���f����s��q���G$־�ݙD%!I�l�or�&b��i-9��D��?�{����I8]�����h�&�H?������ 4c��~��j`壬����+Yݴ��z�lL	8|�SLT��}�'���H��������9|V����鳯L�! ��{��������Mϡ`
*�e��V$8�O7�=�g=3W;���Q�M���3��o�R�,�>p�;�xS*��g�^�j�g?���ѹϰ�0�ik���O��p����]��f�V�ǃU��'sD���{�=����Ue�±���-�2{�^H��� ۆo[���m�����+�_��EAA^�U
�����!(ĿBӯF@^��?*��紉�P��:)��/�� ~����n���N����öQ�*�H�_F��}��!,���bw��Wۖy��}deQ��\C�`h��(���+���_l�N8w�Sد��E�6��%�6�e�§#���_K��R�v�O|��Or�?���7�-�a�*�z<GĹ |�BL3��D���c[��0�u��#�������!2��J�G{\\\GYY�ί�.�
T>}�lE�F�Iʷ?�M�N�o������$���ةA��E�f;��L)Y�O�a9�6}w�,��on#�\�P���;P���x�����/�u;O��ZC}�&�~�������;ym=YHZU@
��y���NOG���2: ���̴}�v�6��7���"d�(#���h�&Z0)�X�_��v|؄�N���|q0�T�P���A'`��0z_Sɻ�X���C�f�m�����
Y븀<��̠n���t%�	���d�A���)/ e
�US��������nMYz��v���Zf�D���s �*p܆�n��]�N��p<��� �����]�Y16�OpQ���.OIl�sM����п=7R����g�iv.�o����}b�gr��M����>��C�i�mq��6�: "�ɢM�jVH��,�}&�f�H��	U���q�]-���͉��70s8�%�dq�+ű�j�XY�x/��5m��;�����8���������?��B�ѝأ�yI����"�m�y�r{G{�?A��N��}��^3eR��"q�(t���?hP�U��a�&Q#3Ħ���E�nN�x��'v�&U�۬#W�Ϧ�\o�sa(�k�Gh�O�T�QWS2�Eb�zB��c#��$C/����(�v=v=9���u�Z1���G�Znj�G\�Yp΁��wT��U�H���:�#�BP̟����C�D�����u�׿v9���F��G�U x���HV���j\WM��a�-��G�I��Ԙ��-m��/m���UP0v�,z��>a^��Ⱦ�z?ز��S��e��Ci�ĜK�4p%]�N!�d�Ϩ�BW ��k�����(_�V3G܄)��5�Yj���!�b|"ѳ#���UTTދ1��r��2��kP��N�i޾�$�I��^�A좰�.rf��`��8i�*!0�y�?X|q��6�IɲV3��{��O�������y���x�Y%���=����FoZd?K�~��
�����C�����{A~+���5ӂRw�ٸ*�F�o4�7'�{ �{�N���Y����O�4D�^��c�y���"�Ju9%W��ra)��]2���z�!��D��Я0���<�x-�ݷ
�3zܐ|����Wh�x��\����D���J��AyEx�1@�(�q�c�1�C�[!V OK �C���*����P��И���z�� >.�ht��R���%^�@ no >LE%��d��wx��<�)N�y�04>®�|q..E�I*6`�����(�Z��^k����w:�Yج�o���KF��-���GP�X�uM�c����39@b�����=��� ~M��G3�l�?�
JX����"��5��ʡ�w�vC�&!�2��Yu�����wһ���j�ޥMoy�/�� O*J��ts�x^���(l�������k���.��������Z�ގ���M�%4�3�p�+����c����}��8�����µ������l�q����Y#�z�X�������T6��1S�������g^�u��j״�a�_i2�5&Ry b8�?���i���QLݡqn	D�/mZ&�3eS�zJ������;7�<x�N4�Bj�b�w����|
`�Y򐆈~�!T{�i��{��]D��.ɼɹ�zZ+���!�"aJfQ�}��/Gc�lAP����Fc��%���y�ڀ�����ii��l�7���SE��;T��Z��N��p_ޟC����x�hg���J��m٥�;�qr�R��e-%���xO�Y17"h\�F&����:�.yT�?���Я-�K�S��'�7��
 PQ����#�Ty�9���5PJ(� �TF�����F{p���x���M�[D37~�i&��'��Mrnʫ�v��B��7I��c�ޒ���_����j��j��F����}1�`�x�'�v8W>��j���2F�?
����
FR���h;bo3ڀ ���wjh�m@�yS��qV�k�;��2�m��1���W1�p�����7�����8�K�۴���&�O6�/��h�f�����<����}Np��N�yh���9~7
y�nM��.��K4�Cc��_F��Å;���(*m�^|�}���2��;A>Ç�,�t�a�s�WD�EB<�� $�(��^c2lyD��5�U�5��fW y���"�quޯ�+s<���A/W��֝��3ٔ�5���p��Ev�ߌ�^�TD�-&=��+%"�k..�Q{/��B�� .	���"��˰�D�һ5�W�1��Bbn��u���{X���rD��o$�t64I
�pV
5��ж���Ñb�
�_��'}�vd_��2��|<S�Bg��>�HV#���4�v"s2�g}�xu���Q�,;+�<5X����ż-2�* �jܒ�Xy�zff�v�v.B�>��3Z�}o{���*��8�z���eі��ڙ՗[��8�h��	@�@� ЙI]]�!�����A�g޽�c��#����#����z���VBՒ��]h�n��//��	>7�+(w6���ƣACcu$'=j��V0����&��'Q��)��"��6��0XP����D{��ǤrQ���QX��n��g����e�{%`?<+E�	������ID.+D�,d���պ�TF�^L~�^~�A��^�#�^=ZV�	O��pS�=j�DF���-�1X�H�I����#�W��PS1�����z��.��a�a]u�h�@���;i�.P�<Rx�>c�<rr���19EGu�l��X:Q�d���� ��'�Z��t�g��'1��?.T<��X�V��T&&�2�t����?W��kȬ܈�K�n�S�;y��>N�%��R�N�[�eL&�|�H�O���{�t�D�h��H��wyZ�6���T�)l8e�ǭ�v�ʂA|�&���Do@0�juʠhI�y}fja� G��a_@��^��Q�����M����E&}R��T��7�,L�pS����l�c}r+u�r�{�{�]�5������(.�&�ޯ�	�M`<f����A���Z����~{c�������	"'ᬳ}���67���L��g��ɋ�ɩ���%��Q֝�&;/��eb�m͎���ެ�WZ�5��?�7���|y����HFF ���>�Nm7μ�a�`z|GB�J��v��7�$3-�i�����m�4!�2��\�O��x� Aq�J�m��$ͻ"��+��f|'�u�
�6QH#j�r�QM>jV�m� �<f�b�w~.e�ёލ �j��*�5-.g�1��ss\:�3�+O�|����!L��K?�m��
��毉��׮1�q4_/�1
	�&���yN�,�%C�F#/b��;�b�`��X����I���֣���0SK�b6�p��a��0�8�/����w~��wL�y��5�Rgo��^^�(ѹ���:��I�[@��Ո�a�[�I�ZӨ������j*�|/��x�\�+׺^O�雏'���dф��ao�^� ��T۽%��An�������oS]�el���}����~9�s�f����!�F5t|x�RI��L�F��O%c(`��A�O��|:\ɸH���7�&�X�z5�R�di�$��>�6j�������s��A�$ه�J�{������1�<�N���O��2�J��Z�6u��񱝟׉�OA9��Z�����|��lط3S�(��ӲK�NMem�ƅG ���=�jX|�URr�r8�"�&K��\oU���XU�O!���u��(~p�PH�|V���T�s�ƚ?>����A�)w#����nԭ5����LW���z0�0�"�8{X!~35�����~"%��ӕZbU��.��3���eKC�Ro��/s�i��zA��j�]?�Z�� %eX&�b�
�֗�����8�6l��J��� %��R31a��֞�N���IT`��]��Ĭ�H��W�j�2�V���n�h+�.���7)�ғ!�3���4AT����&.�7��9����~�װ�Y��ʢ���ќ�Ƥ�B�,ee��@lWHj��mE�	��G��3�.���\��EG�'�w�o9-�0��s��{Z[��C�jh�w���K����S�>��an���3��o�o� �fW�^�	��d�V����R���<��P�C'S�߇B�lBV�p�� �:֗���V%or���mݥ9�]�h�y��2�G]qndBs��L�FO�p�G"*���5ǝ����M-��W�|S������\�'�u�BQ���t��8���pu���˽&S����q&5�v�����Y�]�'��Є�w�ʒ��l�L�Ge�S�����m ���[$�K1��X�Vu�ϖ�Q2�R�g�F�ކC�ّ���_> x�Y�p��ͽO����ș_���fLUhfH;V#I��[1�(���IM��˽��B���*��C����߄z�� 4D�葳���q��]G����z�;�'���.ݼ���ⰰ�HT ,M���`����O�f�V�寍h�6^A����(���t+2h�b
�"����_�!�h�JYx��W�ϵNyo�C�nu��>B,ۤ6,~;t`?���]����M@M]P���"x��ۯʏ�� t���T�o�P���3�����掟��0�1���tK�[�۶�Yr��D�~-B�&�T�%�u�k����l���IO�VA��6T��:H��	�?l�$x+Ov���e�S����g.Mt�3��K`ͥ��J�/�4�N��}0�{S��n�/��YR����� ��^���@��7y'��Q�T!��o���HU���3}A��d���y��K&�l�/��s�������5w@�[i���~�A��� ��,�3݄���	�6�f�M��ק�X<��m���~�~��X0J�{3�D�|� t��H�������)e����P��H?��O�$���g�>��o�oa��s���I���h��#��|��v�)1�,������;c~�Yj��}b�N���vK3��0�O[?��l,�v�T�|�sy�x���G"7�5)X�O��jf*W�y���ﭫ�.������t�Aliҭ+�&j)��1NB��((��=q=��nR�ɦI���2�rȲ��j&����I߸2gc	���������H�y4bY9�����(��w�˾�t��j���;�k�`dx+���{M�JT�������Z�l�t���|��t��\��&��}�i,w3]�c+��?l%���m�b���9g?%Yv������LV�Z�HϬ�^	d��������j�J��k��x]�E�n�X�E&6c������DRZ�i�B��S5���ug��Z��'h�NN�0����4$����\.�{ށb�i���h��
�Y�2��Wr6뎥$��M�0�7"Z��Rs4� ��Z���O�88%�ʫ:�����4� �g�g#-��ڎrӳܾn�Bax�iȷ����`H���ϓ��b��׷�7�J"+/0�O���N���AQ5j-�ž4��y��xQ	���$)��.�?�b<�2$�>a[g�s�����_��:���zZ+�8��g~k+�X!�*�_;��\������	�B/ �&��ө"���ZۂGנk�0��ڦ�_�KSM�`�>�n\�A$�mH��.�ؗO�C#.�AQ��Y��ZX��ug�<[;�ʴ+�?�Ow�x�O��VaH��u���⽈8 [觙�&F\JO��-�I��TӔ�[���E*�z��C @�	3K�>
�g��;AA�����\/�eԶt���F ���PmO�;�?�e�9A���o�ݣ��'rw�(�bA�֨<���Ű��	T���Tշ�sv"�x�UE��t�=�f\?N���KJ`�2�,5?���9������e)�7���P]�z��S���TAe{���>�{[�NYi��^�;8��D&��!���K���X�p_)����^��U|B��P�8�4��HڄT$��^�)<a]!A�7�QC6�������M�f���t�O	ib<�����?�6U���KѸ�t�k���`�%1+E3�`+1��+�d��xu���}��j���$�L��
lwH��IH�������5�=aݻYH�W� U���;�ꆾ�PE>%�*�hV��"L��L�K�!���3�}�C_��7]P�L�E����D4<+�Q��0�^yX�Un/��e@y͟o�B��V@���k�6�t��c�4�S�_� �!���(V�<��Mhh<s�!�t����$��6�L�¬34��$���!�'P�D��nm�Y�|׎h>��9��ƣ�Q	���5l�^͝˝n����*���M��s�y�Ț�<��JA���zKP"M�Mm���z�7��8�tA),@'S%ѕ��,*f�����^�����Xz�2�P�DT����.7(����e!X��ā����h��&S�����@m��Ra`����G4��	X�����썶p��[��ZQ�0�^G�l�E�����Xi6���Ե��a�"A�t!?���y���C�M��T2�]�6��"z��9�	xA��F��lq �Xx��X��2l�c�Hkƣ����5��3���.�J4��u�Z�����i�����]���e�`�*���A)/�@B;���H��9���9�L+�o�T�����B�f�^~W�I��M2��CZ�L� �U��E���dqM�&4	Ln=W`̮>/[鿜��2uqHQX��=����'�3����#WV���p��Q.���0�c����f�L׆�)ɗ�qv�70-ND����?_���oc�������+�D�5��'����V/��=�ً8��xy�=	ĿY�4S��Iω�ױ[�?��BY7�-�~6��n�lyv�Bc�pȹ�S�W=����t2	����hQ�0�S0�[U$�\���V+����Ի1�`��/�,y�y��,�.}b�ߴ��6e�@����%ˌ\n���,�~��a9ޙ]Ow�!�l1jN'}F6%ڿ�6�M��/��XU����Q��ʸ��\�8r�z݆�?Ӓ��R��k��3R�h>��'�N'�~26P���d�5�t���nL�uj�$g�q����0����E��]LȰjF�X��_dB�����K�w0�Q�(���/�m��y�uQ��V���M��Ѡ`-�1̏��/:��"c1n!K8�I��*�	5U�����l�L��w��x�u�Ug��v���VZQ]\'DgK�]���$�T܏��Zfh��U·�L�E���\����M,-�HӡtǱ��2c3O>�*5}t�SL0��'<s�hB���>H����%ѷ(�H�V�7l}n��XE<����~mx�n!�&��Nc��7����s�b]#_��m`���J�����(�{K�����6p�F����zv�������a������t�l�9�ǍͤUԺB�d��U��G@�s�h�6�����4� y��H��6��Iȓ}��ލMN�95��Qұ,\�]���fY�yA�������zB�I�b&v]k�=5�[�#,�^�(=IjjSd6��:�b�^S�RR����D	�~|��l�* ��!pB��h��9��A�ԗ���E{S��E�Y.lZj�H��-o;�8J� )��gL��$�8���D� ���X��o�?�?�����XL9�����'���Ŷ�S�5i��Ki?�b�ZʑV�Ϣ|�t�4N�<��z�|G�����'ex]&�V��C��#�t���;W1�a��֎�ݝg�/6�[O���}/�_�<
.�1�җ���H)P����i��-��t��Uf���t���.��9t�J������`8)X�i��F�џ����Ki��{�P<��o��@E�' B�H�k�|�?Fp�B�a!���鏟�1ǆ�{O����\�~��K��=E��B�AǑ��]Æ�=u9K��Ǵ�x�3�?y�3(�4�,��B��!H����H�I1�I����r���L��ڙh@��9�	�g�A!:ӱ�]E���"�����)FeTdZ`����d���xR:�\��me2��g�h/���^%�A�Vpu�"o���䉈�][4����X�l��ѕ7��qG�T�zd�$��|4="�wR6K��T.�c���&;�Y��xb��&*����ĸ��1:g>_O��K����?pg������'��:���x	�{���z��Ͻ䃎J,��\Ř�ңp�UL(v���j���7���$;[�/w1/�A3�lQx��������`%�<�/ey��C��_�� ���]r{�!ou���bM�%�Fx+�+��8�K�3�ML��S������h���c��?Ѭ�:�[�7�s�P��Bw�a�I���g������>c籋(tl��W��x�5�^��M����r2�Wm/ @�EU�-1��܂�r�ՐM}�v}9l�iB�P�1_^�ȥ�j�Z��+8�5�kW�5f���!����l�վ�ǃwZwY�eB���GH�%���A�#�<X�s~Os�s�E�Hf�!cL����l_8���
���ƒ.T�p̶����͹��UN�}�gߚy�&���%�F����Ұ^�Q@7̸�����u�X�Y����Ũ�y�T_�(R�TD���)u��t�!���	v�9��HZ\e����c[��>����uq��|(��iO!�R���8%�	[^���C�B&H��H/T��&[�/��Gmk�s��w}�N:�c����� �fIrZ͟�X��S�˫x��Fep��'�� ��r$�#��H���Lt�MI����r�ػ�l	���bl昳\�y�.��s��%��a�젾!�s^/�J�V�ݜoZ'
�;o�{��a�!(�MN��I�;J�u�X*$S��#�/BF-��t���˂��cg̽4�y�d����9F��2[_�N�j����c�ź��' �k�EN+:���v b΃��ƞ��,��C��䧺���bR)����]:��DV�2��<j�3+�}��V�/���.�)NpW�����y��G�|��kևю^���jj����"���!y��h&N�T�A��aL����Д��E�M��k�Q�	�ma���ȷ<Hm7ٛ��Oܨ�R��w`��D�yF��מU��X�2ig,5B���Rۓ:e���3p�װ�y	�TFC�otJ���D(Cu������`��6Ԩ6��w~Ϧ���\W{�IT�|�5$\�֜�x����%�l����3n�9]�B�/�[�au�����G��W28ԝ:P��􀲿��dv=	(Q]ˆ�̥�|;#ЛG�t-hw����"�,��ؗ���Y�!��(�+�Y�O/T��Td�c�����V|M�*^�Z�OcJSNo~i�'>��;T��;�ؿ<BF��j�@��.�1,�������l۫��2��w)k�jٿ����Mg�7VOX�)_R�p�<q*��۽��K�������:v�댍>�%)s{��8R����א�
��R㫕�Ɲ,��.��!��t$yfI��y�)�ϧd����H5� y�/��"pN2�z�jF�D�^,���;�G��#�|Z/��q�Y���U����8"���ЩA_E�Vʄ0I��ʡ��V!����c�h^��������9"�1�NS���Rʤ�Fqُ�� �����b'[T�W�)��ʢ_� Ӏ#)щ<�:G7 '|�����&�T)�G(c��nZ|�����w���g�o��T�6�~X##�3�A"�ԣ����%�W4�/���E4Zwa3*�� �T$I@)}s?��_��h�/y�(HߍOq���6V4����r}`m)v���$�j����f,�z��؟�ǲ�XYm�y�est�oLdq��%����x�˿!�Ϗ�h��E��ͣ�B11�&Fء�i��O�%��]����R3�
	�<T{�k���ȭ)Y���%�l!]�-|W�"p�{�AL,~��_�s�\~4���e����{��m��-#v�!����Y�!��{�(��|��&�� W�U�I�nZ�� ����;�������~#i�Mϵi��bfl�-o�>K?)���$�n+��䅴������X	��L���A���nޙ��Ɓ�i��N�X�mk�X<���+��v�;b���4����S��>�����=0��I��@H?K�D��#,,���T�TSe��m�[e:`HX9��E�<�K�@ĭ⅋O�[�FJF�Yp_!I���E���i}d
���qd ��MSD4c��<	eT\*�
<��qC(�I�6��(�R8Ii<�S���w�|8Hi}
sA�CF�|ü��j����_��ܣ��A,��]�O��*gJ_������b@N�5��1d�e�+���M����1/!��f���O8h�)�G�N�n4Θ��.^�tVԬ��C�p�~�>�b��ewK��mL^��Eﳆ�~̺W7��o��j�?� o�F�q�^Q�P)G�=��X.��<� ^C94�5:)�*g�s ������ Kx�X�e0��XH��!e�j4�߶퀐�����Z�ttt]3JfSi�+���V/?��tq���	[&��.6��:��_��o'��->�3	E����N�e�ϫ�S;O��ܕ�ʰ�K�|5�b���P3��rGB_���W�&���o�r$�\!��]���kF�&&�%�'2`��5j�4���E���à���K/di3-N!�'�i�nRaf�;��/���;p��}�����^SU.�6���:v"�p-p��%�I�x\g��Q���G-�eb.�M�Y�'q,���wj�Nb�9il���W����8�1�G�V��].�_��mSs���h~$��+����BS� ����٣���u��uY����@ $j�N����R� �c�\�ϙA3r�/Bv���(��p�d.~���l�Hd���*�?��l<\���?��:4�k��'�[�t
N�����!k�9�`��Bԋ�E�NZS��Z��
�Q��0ey��]�n�UQC]I��~�Y�:���Z�e+���G�z{��BA���x�%a-�����7�,�-{�����>�Sс����@.OQ���"�ߪ��GL�V��Q.X�6,H�E1:�,��?�]��n̔�R�SP �H%vˆ6��eF^����=��W�m��*{#�I�Xb��>�|ĭ����wa����ED�ȫu[\����*G�Gv%*mkΕ���O��z[9���h���tFHy]U�=#ַ�Zg���mVW2�A��Bر4�)��W�tUH =�:vGySd�d�8*� �bb;��;��]���!�6þN�m�D��U���T>�ƃu�	魖�.H)nF��)_�x6���3�
�ztu��vq�(�΅�Y��^Uf�g���o��L����5�����
�{6Y@0��WKc'�sE{�%�s�������� :d�]���P[ύ��\�R�M��-�Y�2	y�/u���D�Q�hW������_�J���bF{�]���>'\��5`���&9)Z�f:�?a����������5C��D��A`2��&������R+qki���/j	�b-��/R�\1�O��m1:����'\YH�>ݑH���͸x�K%��ȴN���pI�khW�Ib�O��"̺�E�_��kG�k�%�����Ô��b�Cz���1J�:z��3N�h��w�{��N.�̮��>%6���(�k��p�HK����ƜgR��gZ�x�)����(�fy��/������T,���e�Nm�|p�v��9Gz���DW;�T΃.R��	feNp�2��N�Mt��\�"���[�����X�"M���Z�BZD�pe�sm �"}�j]6���|�IJ8�:/��t2�ϝ@Ԁ���6�p��@��G[@x�b��FEO�����lo��ϒ(���ۖ�ޡ��զ�ºoNcޓSS���WW����wȧ���Q�F�����⨲���7�����̽꽗E|�bbyxsH��wZ��J���̐�(�O�ͼ����`��]�en#f'J[.v�l���XZ�4:u{Td�8%����ɪ-�-~������]�dLo���2�D���/�B�����E_c4n}b_�=�����,��mw�!�����D=Tob��kj�-�|�>�>j�c��M�d���^r7��b<K<�$���N�p>��3�|�6#� b՜��yጘ��oj��pu���'�DmP�)�<�|i_V<K� C��M�����-F75��3[AC7�%����L=��p��1~��s.4�۴��2��~�'�Jw�$���S��.��E���W�NJE�1L�=��l�x('j�FD�w2d�����`�]\�9��bAg�*z{.���JA�Y�%v�mk��-�w��J�ۚ4Ka�
��y�7���z��[��R_$�s�T]�.1�{��kKZ���{cq�r<�KC���(�.����A�F�`ơ`Q`�7�A�z�+g����H}Q�G��* t����6�R1��(8�~d��������@�@�$���B��q?��7Ñ+{#}�s��+� ��И/�7���������/8q��=Ƃp��u|�.�i����.���#��Z�f�9�@E>ȗ9Z��;W��	
�&Qx]@��΄���<�]�!��,X+{҃(eS+�l~?�y�1�rGEW݆^�??�@cLLP�0$"ҷ�?nrDML��H��e.�A���W!�%�	k������Oc	�x�B�u6���3��k��f�m~�[��'�9�",�x,�����v�q�.-��g�_�c��~��k�"��g�l�}�a����Nqh�x�g4Й@����v+�p���q2VJ����y�<�~�3��ѫ�pM+w�p�B��_^��Ā)WK����MI��I�>�"��⅛���׵$P�>�4*Bc���nL�̎�t�F3�6*@(��C���� ���䍞�|��7Ѳ�1ZԂ�[�_�B8�I%j��*�&���P?YT\��e�L�u�Ϫ��7+P|"�Y���W�v���zx+]�W)�h[�1��ܕ"�����(=��L%����y�ɀA]�OM8�	%q��b2�i)��
����8R���m�V�@=��z�:b��=�s����@lY�
�TR��<�K�`�����`�h6�]�	|Y��|�0�?�V��!
��$n��n{��P���4�㌐X4��R�o�*}WLT�>[�����ۤ����%5 �21�v7�;Y�k�f��@`�J�9�d�Ǆ.��|x����s�7�Z	J�t=fV��5b�;��(Fn��v�;g�@��0qݤ��Bd��;�M����|�c�O��֑� U�@�\,V�d��������A6�z��Q|�ڪN�(9�f�Im�Nk�j7�X�g��M����B�
��ڠ�"�7b��:��J�AB�{�=���ǉ�ݵq����c�$V/��J�pŇL�琖o���$C��s.
�ۨҩo6@�4����sY�Y�2�笭������.w�)��ꍦ@Jl�ݮT�M���ݣ�n��	b�p����t�nt���>��R���.n�U�� �l7�A��a�`I>Č�˻Cέ�2�n@�o�H
���|��Lk)�8Κ��"��}Mڬٵy�1�~�S7��{���\���w��������,4NM�_qm��^>_�U�Z�Y�X��l��~�d��tL_�iUW��w��U`9F�6�����qݨ�BaG��ғ��d�u�3�C����P�6��J�k j����ȓ�kg�����8,�Rx;� BG�������R���B�hm�nE| /���.��SSSN=$��_�b߹w�
~Y)�M�B�κ��ܨ��?/�O�S�s�oZ��AO���W�^#ܒU��3��:������G�fUQ�M\��,I�������-y���%���?�N-Tnj��7+7�T�7�\�v"d�ʊ
1f��v��uS,f��2�o�.;��͠`0L]2���+3����.�B����L��J>i,�U�����/dKA-�v�����B�I��
�1<�^S~��N��=�/à�#��N����O�\����Ь ��xb�܂�٥xP�{V������I��������SZI�g+n��1϶
kҠ�)q֙�]�p4��-Wf�o}ī!��WEs��֌sLE���L���2A�FD�ٿQ�O45���^�Q�L��i9� \Baޤ8uW��L�s�d��qNUS6�JiTgT�ܓ"sa-XTOˠj�L�@l1�VH��	)�W�ΦD۔�/�lu�U���i��"4���SB2})`y�Hl���Bc^V�<�cpJݩ�`���}� c��c˚��7�S�BI��"NU�G�\�VQ�E+��C��D�e%�qz	�^;[v�3��I�L�C�q�YHf��rQj�`���z?,���T$&�M^{���n����s���E���B�]e]��/��}i��\��[\����*kE���B�mcG>��D\.s�H�����P����u��q�mAܵ���)q����-պ�M�����q���TP�;���ʝ�;~���)1��)�%������3o�֐m��}����#wO�L��� �vT�~���		��? ���l'7�W��2 9f� �4[b�z���)%ԣ�{I)����� �@]��#������!�-���J��c�+�%:�m��f�(ez�ߜc�YвV+>���s�u�fn������I���Ul�P�)�ǋW��賰_�2L)ʵ��Q6�Ax���gw�	/���M���C�ݓz�L�S�'�x\r����×f�9�a �Q������FC"A�N�b{�=��M��`�_*�eD�[J�S��Ԁ�Vdg��9) �EG�C�ފ	w��eAF�a�I��!��� k��35c������D�k8՗	R��;�.��b�ڊ+rrl�Р�
	8?��g����x�@�)Bl�S�N8!�?Lѕ�0C�Ĺ>�KN<����x| �� �+^������g���6�M�Y��0Q�����we�Z�@�0�
�yӛޔ�w���纍���u��s�'�9�~���W�����`�����1xŊ<��L��9�Z�^~�Eu���r��}��Ҽ]O�/���ݕz�V�wݞC����Q�kH�@먭�FO+�� �#������/~q�n��D��Q�
XVҳo�]��Z]�r�E= zjq��1��@N+c�� `F�S�=u���q9��Zt�����O�Ld*uۉs%^�v��d���Tb�Mh�Ü�!q��Q ��m�C��0$Y�\88����~zf�_|q>�{�J����ʤ�Y& C?D&|��_����Ȁ� �q��B��b� k�<Ϣ�Qv: �C����_�>K�<����`�1�'�@�K�ӷD]�<�(�L�����!v�$ �Fθ%R��aׁ0Lx����h��=5�gR�#*=ݩ�ڗ�w[c�*��2r1mrT� ܞ�KePpב�ȱ��S#6#��T�
fZO�0�3U��t�i*���L	�Q*�ؐ�T��
�#3U�3�2��Vj�v�H;Lq��Id7|����wU��{�Ȅ�n�^�|�3�fˆ�@��9�����$�=Lլ�� ��3����͟�ɟd��������h7���p�'?��p L������
�I��rl���r��Z~ٯDCv\�HƫK�2+�`�H��"F�dR4���Mg��9ޕq|���s�,77���'<;�Bݩ��|ڴZ�.�#��~��[7ϫ��ݖ��&s[ޏ�]�)I�49NOdU�21�����kF[��h�TH%`d :�"L�LQ��Y�:���0�9��t<^GpSs�7�8E��c]�n�Yb�f�L�>��U9Ǻ�םj�Z�2�O��3�,��M ��h!.���`��:�b�s��p�3����&�L�Q�����.���Mٜ�s> eyZ�O$��K� E�J6:�@���;R�%��Y�83^)��Z:�xvC������F����\���rD; �9G6ie�����t�v�:0S%�6�{��QV���e���eW�C{b���vU���d:Ʈ.S��og:��:y\��V��} 2��ѣde�X�W�.d��	q;˽L��i��_@f��l<�3��,��9ޫl��g����8������Єa�0�hw6gu���~�j�e��z���-�	�@�=���.�&6�@]M�c��ϻ�p�C��e����jh�:�D��||+�����j�[��s��Ϧ�(�	�o���|*m�
ǲ4�5<���'\�����#9R*3ǃ�d�ѡ�wesmw}q�pDs�����ɮ��+����eH"�>��@x�W�Y�欎�������m7]�J�`ٲ�/?p4��4V�9 ���ifG�*owꠑ��iL+�a<m�	��ɴ��9����R�w�39��X���Fd����9��3�@����+��e�Ɠ�{v�Fv����b-����J���m��I9n,���~�}Fg,W�]����I�^$�)^�N/PD�HA�qz'���1����=��bW�^f��ٛiVciP�-_��h���>���y噒}(Cd��i[ATPҾs�/�jH��r�w�R�Rc9d����}#�R&%>�,6J;��V��?��q��LR��Y����O�]���p�#�n�|�p^���1'Ǉ��3�&G��:T՝V��S�q	�g����f�i�H�S��2�3�g��_�~��h�ZM�:y�v�S>��?���.�I�2�`�{3p�vY�q���t^�R��ؗ���<I��x	 �|Wէl<�|,K`��͑��s���f�`�mF0zw�R�̺u�N?��#o�H}��ʲF�	�� �մ��E��)�^RW���E��hd��v��Y�x�*�����r�:�SnU�~ou�V�G0j����X���#j�婴���-@Ff��;2j���Z�M��yO��+���X�0������3<�(�,ʤ�2�7��U�� (�-�c��s��n�|�p��ㅨ��2>��SfZ��y+�G�h�܋�1LE)BQ>j]�u�V�G���j��"�+�ɛx�`��f�
|Zw�f�<������FS����Rw*l��L���7��T�]�����D@x�:δ���f�QS��E�7c��]��}z���-���c�N�X����""A���N�v`�ʲ�x���׬YsZG��	/������/oo��;;��c��Z��<FR��]5`����`#����>d&��d!w���ޛ�Kz�����=�<d&$@�à>8]8W88!��H!�	(I��4�� �E�0	����9W�<xQ<�	��t����I{���ߪ��~�vU��ݝ&���~�v�7�o�w�����w����C������Nސ�{��4�?���u��Vq2Ĕ�|6i�B@��^����`x�&.;��>y/jy>c|v�t8�s�i�u�F(�Lޙ�Z-�z��R��J�Z�>z9���8.u��aWX��b��vw�*��6\)�B��w4h����� ����;A��ױ�;󌶣��+l?PF��ڽ�a[)+,�x��ږ7��E[�X��$>�P�U��;N���p0�r8�AaP�;��fo�?�~%��ˤG��L��a�e��!�JNpƮ�jc��_q�[�V�;kl��OW4f�&wD�I�v��A��{��M#�+<�Dt����r�2��xm��GOS�WG��6e1�[�v���	n�;��C����QX�������̵��8ײ���SO�N;�����9�t�DHT#��6��T��z����2�;�t�q�{sv7IPt�YZ��M؝��
2�����בN���j�2��x~l_;{���t�lo��{rڹ׋$"��*��vsH�bt���k��*�����Η, ��6]�f��ދ���G�T�h�����L�jc�����O���\����0{̭���?]�i��ARw��lg�n�j��޿�`��X5gn1CЬT��Y�u1�/�h�Le��.��iԢ"�Q>¸K+լJ����^�J+ѐ��k���wΑ��y� [��,��St)�n&�<qW�����ò�Z�m�W���w��q��2��`�إV3�F��|��<��z���w��P�o׎V;�z�Z���c���!��\/���{Q>�8�]��22m)��=��k,�m�Q)��k^[6(��l��`�,��F#񐱎���^�l�2�Qqb>�a���MY�{�s*�r�HHr�V��r�V�]w�UW�jI�����;n�̺R���Ä+�RzԣN�L���l��/N�H�#h��ei�y!8V���e�s��;BEG�!�d�ܨх�]D���&�.2i��\)�1�G�^�@X#��x}^܁,v>�5���#덁�����An�K��ۭ�y!�]/v�R�ee8?��^b;R'�(Ld��@��<Z,�'QI���c��K��!���ǳ �<ܯA OY��m㦗`��b<��B��s�$>�ed���G�х��R/r�~�oJB��ȑ)K�|^��B@z�AY�s��&c7��"P���|�dL�RO���Au�wl;S,�f�v��M���tZ�Z����v�EK�O|�N*m����q���\5=�'-_�2��-K�{�/��ǬLS�>���rG�0��Ep�x*������������.�hV&�����'S�Qʘ�a!4j�S��m�N��`#;���\��+�� l|�7x�r���y8G�F!����������EcLf�r��B d��c,ovfoԜ�VK�@-���mJ�F�tZ�Vj�j���p)M�v�n�<Q��R��g��ZKs�-&�Ʋ��q��Z8�>�ff�a�A�}�iD�����Bo�kE��s��%
Μ���
��[�Bd��3�+�[��a�ڼ�5�=)r�������zQ^��Pzp�n�Ȁ��00�%c�a7q��wq��{S�uAuKH�	q�l��v�Z�^��˖���8���K��u�KW������M˦V�5����^v^Zw���h�S�Ioy�1��L����l��	����IK47��7�^a� �ph��Բ��z��YfJ���Iৡ�%�G`���q�?��@б�.��>sv$��q� &�|@'Sj�H�����{$\���`��9���2�����K=��d�m���s�Lw�;��� ��	˝Tj�ScvO�4gR�4�j�N�R
L�?��� �K�T�J��e��)�jm�9m���|���Ԛ=�;�8;��@؝ǩG���DFL�b#�=�.��Z8�>�od@Sk�ހ�KP���~a�7����=�D� �;!G�9'�+j�(qu�m�p���ƿ��N23�گ�Z|�%���ʖ�CdO#�}�g��.qv;4�&�-�)i���C�R/�P���duR(�,�[R���sL��ˎ�o��S�{V��I�Ӻek��g�����J�l�9�l��
uD�*�
#����/�A��R1��#}�@�zq*�J�0HbM�9ݱ���0�0�s](#�I!H�����8g�w �IƉ:F��4�ܫ40�IM��Y2���:-�b��#��?FFbor7ctb��Ip���:w ѭ��)�k_��\>@��_�j.����G?C���g���x�X{ww��>�y�/��?.�����4���T�{_�vfS���Cw�T�ו��y�;�SO�e+Ҋuǥ�D-�|`w��W����1u=將����B;#O0���P�7o�^ �F]GF��ɹ��ljp�%���A�w !�ƽ��9�k�17d�K��#�a����e�l���	�-����}�k�@�?�����v��v�n:� y�k�naͤ�$g��@���7�Ŀ��/���u�s6Q8��s���ɓz����IEo��@��D��z{^d�⊍K�;�W]s\���t�=w�]۽s�Բ�43=��_{lz�K_�V�_���_�����D`o��N���@T���i���A�L�l�� [#_(�4�����Ї>��R�1cr�4�>�bg�,��Ʀ�0�j�AS��h?��?�wQ?$����<�0eư1@� &�8�@y ;�b||ϳ��]�ʝ1�5��n�������
x�	s`0�3���9i��N>�Բ�bq���-w(�g���Z�6U:�Ԝە��ܞ�voK��L�4S��wC�dT�Bڪ�Ruٚ����R�0��d�g����O~*�y`W�*2�4Y��obx��{k��`C�Y�\u�U���漋/���+z��&��n5m�?ڿǩ�9~W��N�y��6b ���������}�O�ց^!yzق�~*a�8��>�M��A�z����&������ۋ.�(��+��r>G��ӟ�}0��乭�a�T$_`�7���_n�Z�J�z���.wē6}��t�Mo^��g�n��2�RJ��~��t��ek'�?��?�;��Uw7j���ac&>ӹeY���\v� �mDu%�*�
�qC�#{>9":s��rC��h������p�0W\qE�����2'TР.���h����y?L���2���svW�%�<���tf�x���)����n�|��~���;5�~9p.4P��戈Nw���=3�3�} �ukW�jj�NcWz`�m����4Q��r{&����F�of~�rjWji�]MS�O�ם�Z��4ۮ�=Ӎt��@15�-1?�K��s�zPF�3	�ِ�v�=ٰ�}9��/�D�p�����'�5��0a�Jr��y�X����c�3F!p,&�7  �����D�6��3S.�4�ͩ��:����U^�n�����DٰU��5�\��i-���og��>���c�9����{�2�mL���� "ЋqǲpH#������2����\�iӦ��l�r�;�5۷���]_�K���w��?��w�ȳ�j#�QL���]-K��ŀ޳[* ��>8����7\$a��ѝT�<�Q�A��pܓ�`��@�k;� �E�t��(����.L�Q���t[-#�lE�ar��<��S~�2[�Ȅ�;����� � �lي4���W{�9g��kV�j��R}O�ǖ�س#MTfS��Y�n��@�E�Ze"��Ժ����N�ʊT��Ү���k?��y�� <37}X��y�`�.v�� a��QA����:�������b�N�	���{���\_�� ��7lؐI�2����� �eP@���r?���9���F-�S׀0�� I�B���b�S��(G?�����_y��z����#���1�K��u���;���hh��w�<�v��n�Q/������a I��z�D	ڕ#d�����O{��r�Q��S\��q ���(r�$�����1�"x9����սa�L��U]�a�}d�N6Poh�	:. Lgְ���k�M��e���.�4N�c� a��{Lx:��Yg>��{���r=U�3��Zy�-�$=f�e�<�f��ij�Ҳ�'�fuEy���    IDATjt���F�����;YK��Ls���ʏ��Ud�9����l)�0��Z���u��g��Äq�e�Ev���XU\G&s� �er�~�oܸ1�=y  �F��"���[^���~�ٸN�]���ס��s�6H�ֻ�޹�[����/2a۪�^O*�%c�yb���/]�}�KW���(G��Z�利5I&��G��x*]ȇ�� !t�8�{��g&,
tL��^���Jd�g� qɘ����?������KV��԰�);F9"2�x\����p ��f�6�=1^��	+G �c(�x�;�^O/�[��%�޶�0�VN�yu\^��`��3^�"���J��g���Ք��� �J�SOӭZ�\��4�^��Jiz�����S���v���j�?�m��� a�� �@8�罅N'�,�r0a^xA��7Оq��Q�X�r����BL8�����R�0����~{lSc�x���{�gF�H�����C�0���w���c�0��@��@x �B�:����K������ߗ��q!j��FG�h�DG4��R��b����3�<8��m�*��|����W������?��yGe��ʥ����p�x�2]EA�@@��	;"jx���"ƀ1@ga�(����a��Z9B&� g�#�ZV�a��.1&@8�NV�#�h�y�E�1=���rskV�j��R}Oڵ}Kj��@�5�Քʬ��p^�����J��=:5*+�\�H{�&|mᩱZJ�V�m�Lx���G;*���d���+�� ��V,[�`� ��0a����=�����*`L��Ӡ_�=��<[��1��g w�8�#���b	���w�0�G���g/{�U�~����9"t����w�ؖ[ߴn�֗���3��!G81�z��Q�T��dD��3q|<n�F�h;�c-ch	L�0�^A��R�V!��� LF��C�T�`b� ����
�v��d"�	kP��Y��݄	�LN��	+-��9�L��}r��4��)�w@���v=�K	
L�e�Tji�UK����?�µ�go�����/�tA���$���~X�/��E9"�	c�Q���)DQ��Z�N���	s���Q�9By��F�҄#����
��Ș`c>��h��-�&x�2?䜋a��r&}����Z�HȜq>K�;D���> �D�r�R�0P\)W>�q��Y2&�o�r��mY>��	+G�	�<����y�Atw�Q�o*
ed�a�0a�)uc~G��	#�S��-��&���l�P1hX/S;��&L��LX��r� ,�	�	�|E�ӯ�<� l]'�# ��R� ̵��N�9p�/f����l��gow��61��# �j���s��m����&<�A�&	O���=}�SKӭj�:�4��ѩQ]���X�=3�>�'�H�wޗ&�*Y
�kD�]�y8�� ��'抚0Lx!�s�	S�h�21�u��"fg����BrD$&��RL̙��? �L ���!!�� �=�	�Y&�g ��N���	D ۧ�=��Ȅa�BB��	wCtK)]�eo���x�8�kA
�_6]��v獗��~��k:��r�!j�	3� �0#��ZL� &���}o>o� ��R����f�a�R�Q�U2�Sa$�\ef��n4A���@g6�� �L�Ɖ��QR�����K�;1�=r�W���R��+>w��$%���e���_si_�/�gz&�zr�Yg�t�Ks�i�@��4^n�rk�|��	ۃ7Y� J�SK��JZ���4���ԮN�F��=����O\�vݿ3M�Є�~�8���]>+�	AXa��1���A�w���0�	h�Z�����W�l����8A/�&l�@(�/@� P�/�cC}�����%��`BX�K ��=��RF��sW�ƍxi��s�� a	~���.��%�n�d��7�}�D��Fs.k�G�X�k����w�9/֨כ$���>��E�;l���S:-yT8�'0�όV�D�<u����9Y�a@
��B Lc����]Ӹ����;\��o�9���c�+j�>����\ <#*�3�%��;�񎮜#t,+��,̆�}��O��O������"7�w�m}h��c��@0~<
���Q��� ��^���k�涛k�s�=���H�֯J�V+��{S��>�:�T���$=dI놪�"�Zf��jj��Ӳ��R�6����|`W�����������R�3.�E���6�J4�Ձ�� �ع瞛m���f}��`�=�~�d9̫@����*^��+%$J}q��r��r��/��x��!MG��^q�_��aꎸ}"���g��7�pU&�|@�Uϕlp���:+�5}vA}��_�܉I�&�ўMF_a�"��[��Vf�JLeT�奍��L��/a�s�  ��+קs�9{�����F��P4����T��K�g*�����6�����??�Ӏ�Z��!`иѭx�k�PG�<*�5T�����p���x��v��m�c��ѹ��+���3�����q�����3p�7#��z�wup�� v:	uI�v"�r�,�@�R�B6F@0�7��l厲wzw*wHu�L%�O�	JC���vzrn;uJ�t��.�)͗�?$�I�����gg�\�,'�!qζF����开ðW%7�L��Ja�Gam���{�mhk��[��`�\��z\�T�s�|��U��|����+Qh��Sڟsjȁs<��(a�+'�B���;/ u����_�k�\�?$��B&���	��sR2aޕ4)'�f����	� ����m��ǰ�{�	�G߻�es{s�	�	Q�'W��swo�'��< F�ȃ�E�Ӈ���z��X5B>�|�+�7C���Dy�T@9�YN�`�#�tw E����BY�{;���n���\~^4�c��5*#8�g��c�%ǚ��e�<��kG�<���,Nf������ێ欲J��;���r$L5�X�2Bml,��͜f2wn7G�3(3���R�CFo��vE�[#3[9uJݝ���rg�Tx^K��l6�� ����9��;_!�[��ڹgjF}�,g؏	��I�eb(	H��r�e���1#Iq�s햿%�c��R
�k�>��@�}�Q��s,�IP���2ǵMٵ�9��dE�"y�
���s� �sAl�ޭ�'l�믧�a���.�b�'\��u�-7_�n��,�OS��e*9���5��;�� L��
$8ډ�ج�4L-�M������H�{�~��,��Ÿ�[2p�<�09�k��w��ϡF仃�#�����������Ռ�P4b�se@�!2x�`Y)�@�=ޭ;����*j}�2c�Q����dڳg:w�����]�_��J�(l�����xNi鋏� 2���r7��lf<�̴�e��i�T��;k�ژ:q�|�w޵m����i[��AS�4�^+�B��-pm�%@�o%��mS����$]}'�<���8a>,�K�����9DGy c0c�/����"������[W^.��PO��sb��˲�񪫮���SNY���·�t��w���>}4 ܨ�Ҫ��U�ze�#����Dt ����o�v�cX�#G@�u�u�96f���e��m�y���hn��Q@ΑLY��y���)�=���4���"��Y3�]�0��s�G��2;hɠbB"�*0+KP&Yב	��b�֭�
p��1��m�x�,GĐ�ٺl�,h������>l�=�z�}25�����fNٓY��a�|􈔥�;�M�eE�q��H$M=M�\���i/�BU��{��s�;��2_�U�e��-Cq@�?���j>�y�s�9'�>Z,Rk� n����\�} ��O��&L}�f����,��d���F�	��c{u��+����3�8c�bLr������fn6�9N��/H��N���{`>D�Q0����o�[��u���+�뢱2�����?�gBۘ���'?9?)%��9%��&	���$`iL\�g�E���02Y��׭�ÌP�Qɂ��80(?Ȗ�`�r>��f"�y�^2�AL*{�;�ZwϹf���c��ɚ-�h���p� A&��[���;ώϦ�e,ԩw�F3U�D�/�AD�0�M5��Ko� -KS?��M��ڢ����� !����%l��%)1.��t۲ľ�v'�U��k��/���,- E�s=�(̗�)&�ɦ��+�����,�L�9��6�tؗ$�(��L�{�b�6�1�ܰa����~�]��<�>��n��<@xl�����E9�<�����֣̄͢��i�bG��#3f�W��ys`\(��a� /�1Ǣ;�-S�0a C��VrԈ���s-�@wD�����Fg��*���!���6��;��\��VR(x���a��L����>+�*���@�� �����x^|��k���|4��֟ݎ��N��8���gV��:�%2�l���}麉���C�8�AX�l��HF���CQB�]e�\_�I[��;��l#�g4�'��{�����ne�[��]I\��,_L�ﵰ}u�P�c| &���|en��}�c h��|�#�޽��� w�'�-��IY�񊃟�籜��Ah�!��,j`���6m�t�i��v�};��B˄�m�㼩ٽG��*�	31��lot���y�幹�A�҅���ő#dt�?��2aN cbε߄��b�fA��1�&�*�@�gu�ڭap2z��	|�}d��!:�g�3�\�<JCq-�����!"���xΑ�����!$�l�=J9�݂z�ϝ'�z�1 �;�ZBjH=�!�,���Y~�)�~�VsS�a�u�N��+��h��}ɬd�F���H��.��&���Q��DgP��^Ji��z�����w�C��r`'j���g��{>��ًz���JH�>��d��k0Q�¨�<�9��!I�I��)r�zDB �Ω���[Ǒ�Y/Vγ�l��ԽK z}������Y�����^��_OG=j]�7�R9O�,�D��+��y����	��0q'��s����x�.�O�8�1�]�����OF�ae��N����j]�!�ݒ����Ч���9�#��=�%�3�D�����' J�	|�A��'+f���$	��`@l19�9�9���A�_mI,9��7H�׿���9�����7.=fb9��LL�q�?�*S���Lx��`�x�1b��{dc���Y9�	��^3�?�����+0tm�;�Ły�\��
��`���l�N����?�:���8�4��Xc"��D��`�C��8̤��_�vԉq�s>E�2HT��IO.��M�6]��r��w�ly}�(V5�	���W��g�˫�ƪ�AX�(6Ha'�tK��t�8b�����o��[���ԣ���[����} �V"�l�8���t������9�> ��~�<�w8���m8������E���?��qz�1p�	J�?"&8�����b=쨕+'z�b���w5��u���Qwo{٪��Q$[�	��hPմs��4>9�(&ܯAc��j�`�:	e$��ް�aF+yn���5�����}�0.����}�5Qx�R���y��r�����#��?N��	n�6�M��~���\'���W�XLTw1�I�-�V�W*���#�m7�q��-/[��G��g"��j���6wg>��n�[���̣>�䟫���1��� Ց|�{�a�H��s��j����`<�����|�����]]w�u�j`��������Z���A��z� ,�ᤠ��N"F�̶U���,q����	L~�zr�W6n���%�# ᱻn|��{�z9 L�V�� a��L{oγ2,Ns�0o���9���+��V�P7f�~?21w ��=7�n��*�v�;��v�wys���q�r������a��;�j�+#�\�m$��(��|̓B�x������L���x���	��[��֗?�)O!��ȯ��,���nٚN�hw��Y.�(�u3`��[�,�s<�ai>Le�����1C�z��O�3�ar�~����(�@W&�pO���y�AL���_Gd�Ca(��X������g���ԐP%�w����3���?��������֋9�@��SO�:�^��A���ׯ�~��W6�fb�ݖ����Sg��[�D'�%,6�ofTn�+��=��w���T������[̳<���P��@\�{~̝�x���=����l���{��#g>���R�[c��,=Vف>�*��t{@9���k�S�ʠ�)�r��7o���SN9��Ŵ�� l��r�ZjV��)�R݅X��������X���`�����KZMFjK(���[��:���P9b1��	ˈ��b�q��A���\l{ŕ'��+5e���D�$�i�{e��_tԁ�ㇳ5��`��A�\��W]u�yK�y�ܭ7�~��0��c� �q9ڒ��\��s�6� P+��$��A&2�f�{8�ȽnE � �� .�D�E���8Y�jN@��f��u�����)��7z�#	��M�9��;�a�Z���j�Ì��uy��/���F{;��v�#W?R�k@Y��t��#K!y�@Ў��
eCsK�7y]ȯ�>+�Ҍ�in�w��E�nQ4*W� �,q$c���0&���,.۞�(��>�F;r�!�m\F���6B�g$i(Iؗ`����0�o������谍>�p��(���9���(�H]=L��+f�1<�p�d(��G�ɑXd�Er/��! ,�XH��VJF&`��y!σL8I ~�0s�-Yt�#Ev��8�r��0� L���y����g�0,@�\d8r��8�5Pd��0L��~��v�1�v�>$�1��c�̎7l��VaE���U#$GT*��]y�/;�.VZ�ճř�@�`�	;��	�9+G�	��Ȥ���!�mGnv��� v��y�a�h����!Z�u�
�醝.�$� \.��f���K'��	o}q�?���F.�/c �����_�żݒ��ѥ��@8.m�G@xXm��P�@�s���� �0a��[��;�dA�/���~�����!?��s!D��k��D$���	Ah��u2�c�ڞ-�ɺ��6&H���5��r-�0'�L>�;������ƖE�^
͌k��刻����hd�<�Y����[���y7�
[���.�L`�bbr:>�Ƚ�ޛ�u��s}��VH���7�t��`�����{mٲ%��|��e[,⹑����q9�^�B�R�~u�,Wsq^\��O/-ڰ+DM@C�L�+������ص[w�)�p�B�MxII{p��?�Wd��X��.}��gQ�I�e۴;OOH�LܐN�ܾ0lb����b�PW�@������'��S��T�KʱI�a�&'|����`"2CGgwדN:)�b�c���W i\�]��b�<��>��d�@��k�f��ʕu�����Ή���!7�i�������H?��?���_�%�n�S����1���V7vV�Ϡ�f����|�K_ʠ��I��^���];{�3��@�\}��Y]�'��C0����֑�� ����]��^�i�������`��D�;�=Ԍ�e�
<ĸ�2[���g�gyt�W~�~!GY�C4��5�{�����ڇ�T1H.��}�W.]�G�!��H؋���җ�4���+ۨX�	&�C�@0�������{���
�H^�WdVH0�w��]9��k���N.����Q��,u�cZ'q���԰��ߣ���i�π�Fa���.|Da�,z�=��[-]t�E�q�{\�A��g?���c����3��_�u����s];����w `�^�'���9>�{P=Yp��r�D�@�h���҃���U����3�*��    IDAT�SG�`��8�/x���J��|����y�>s�"~�gӞ�lL)�q�^{mցy.�����y��;+��>�����g�4�m��詍b��# ��L��Hq?1ȗ��e�	c��: )c �aN��3t�p�]�I'g��a\�}�{_ޠ�� ���
p�U���5_d'�Q��X�����2b:��Yf�Y뉎{��f��D�'�k�젋����~^��^l�~��s��l����[7$m
�������K��F�SIF��͠�WN�j� 4H
�*���U�
S��?�4ݿ��X����yW���-�{CD(�r �F��`�\�m�b���p ����R~Ҧ��Mw~�����������?l�#��&�@���8&�KÌ�&Ʀ~��adweS��i��?~�{ߛ�p��T+���<kT�AF�q��s���b���xc��S�_�T����Ox�2����:0&�*r Mg��;���5�I�y�c���|�A�B�zի2���������|%��;U3�������������ۜ�Q���m��sd�QۥLN��[���ҫp�,z9���l��MR�h������1�K�,~.GVjRb�l����� �̄'óAF�j$:T�;<�6X�s���W����W,Y*�G
cl�L춊����g�O̩
*���B.Ԑ�_�,2C#G������<�Ą@� c9�X��ʢ� LP�e��b�D���c���]6���>��Ol�
{O�e�����ԑ�鬀��/ǲ�9r������=���;rė���<ؙ��zg��nY��A��p�a�T�:�5~�9��b���.�E;�����W�-j�Q��3��('0/������� ����dFy��(q��w�v������o���F���Q����Q䚥�Q�5�K��W6o�|��S���!a 0�3�8#��I��[tCuU�����	�2h'D���p���ja\SƸ�b���9�=a�L���fi��놌�  �����0B��VO�s:$�#�L��(��ZL�!Gp�TF��L��q����7�1�9��������	�V��9ka�D��AH��`xb.���Aח�r6C�Q.��N�ˉ��ROFQl�Y�zV���v��6�F`�w$5'���<��z��ȤeД��2�G��2 ��W��%H���C���ny� &ܚ>*�SN���m���߶|_J��S���f�y�]u{����-:�����Ё1:.���ݗJ4��A� �@t��&�@e!@LGD{�����g�� a;���� ��_��E����#��֕n/�&���d�H	</� +tL)�����6˶�4�7�	�3�r���|�#�,_9F@�ikt�8�[���A�?���@�!��O��Osx���0&l=�~�!� ���w�3�atݵ�"ip��	�c�a< �w���k�ʹi��	��|>%�v!��y�(g|^�A�;v�P�n�t���Q��K���)���5�[~��uw�q����zXkֺ�����[��jz`)8����{;D�7�4���"�(�p7vh(�ݩ�;uA�c������9��>��W�V�	W4N h�����8"G�(���^���năB'�0l�PX�F�1�Q�_����!3e���o�g��2�
�<Ϫ���������8_�w�I��z-��;� ~��^7�o�+�№�ɵ,'�����p���?�=�FZ���N&qO��>\��MozӼ�<�~����0��'�����alOm�:����7d eҒ��|��w�ˋr	�9O���-]�G9�6R�,��^�[�@x�h��)�w&��pq0u��aus ���#��q��N?���s��<���5�0���� c�} ���+��vw�u��.�r�}[�w��9ǿ)|�����mGJ�ꕢ;�q�c-�Xi�� �����=��j[��O�
>$�����'Ot�aA�^zi>%^/>���x'a��a�D�7M�h�S_�E���l�)��wd�B�:���Y��:���y�[ޒc�9��,�S��L�B�����s$e������M���>��g�3E�0���z�	##`oN�E��{���afۺ�і� � l���7�Xwڅ �'��ڶ�@�����r�K6l��p�{��VP3���/@ ���Z� 
������eR^�cʽk�����0ꅻ��2acL
E��,�����)<��Q"S64M0��ו���F�TQ��������i�2>�z��B��MXu�yv4o@�mܓ�Q�P�����������/Lqnd�z%��Y���M������e�.��V�ݍ��H����as���� ?���̓�� C癉� zV����� �/|���$��~�_�'e��X�\��e�FNP��x�esPs.���Z{� �ddL�2X�p�R���.��g�qƶQ�b~pZ���7�{��;o�d�џ	G~�]u7��~S��v�0 �<ủu�
���S���;��;~�Cc 0����ig�`�w�V.g�3��Cc��I��θ�u	5Z�(�sm�=d�~��p�m�96���&<��3&���=�L�byY��=#X<qp����g?;����E&\�rw]ڊI?�vA\p�-b��vRʲ�@�2�6���^a�0er���9F�	����G>2ow��R^�-�ﬣX>b�#s�1�q��5»�6M��Q(�EmZ��kDy",�	�t� &���/��U����2[���Z��=����v76���Zٓ%`������J�c�k�ޣȾ�u�N9B}K@�5��0&�M&�p��H�x�f@6�������91��5�(7X�β���Ŏ;��
 Qޠ��� *���Y��9X������ d���� ��>�R��(j�N��J �����tz·5��Q���D��v2l�&����4��=�}r<���BR�;��@
�E[�ي \�+m�6d�!��'a���g2Yf�*F%$�E�*���]>A�ϯ��W�r�)�c3:�y�5�&o���AL��Z��
�$� ܝ�|�+�<R�I�n���N�Eᢻ!$���H:s���81' cp.���u�00\%��_��_�bp�Ӊ0NB{X�E�b[dg�9�Y�As�E����ɒ�D����Ʊ#PF�Mt������B������H g�yf�>�Iy�s�o� A>@X W"Xhb.��I�a�`;�vއ�b�+�㱄�!GD-1u��X�GT���g�-���@m�m�M� �d��0�'�m%4A��9ʤm���o��v�hH�� ��D�8����H���t��������HbJ������]�� |��/Y�c��與��0�l�{��[W.�N���I\;�n�t�ob�{nT�=N���ӊѐ�y_�E?�\Ɋs��jT�\�E1��b���#�.X�����ר{~��pbN�j��a�]��D�b���=��
��6�hA8ztN&�.����y���vz�Z�' #�������b]3P,�JF�MqON@��cT��n��X�e `b��퇁���֊ \�,�w�S����@��)}d697`���zaĸ����q1n��1@�xk0�f�&e�]B]����!%�9Qk���H�r���͛7_tꩧ�X��f a�3k�����ﾜ���D����{g_�Cݳ�a��h���}:�����j��0&�TV'��*q�Y+�K��K�cdE=�:���lK0�1.������jpAR�s��Nx�%�<(b�덢SzO���
/�0,�C��xQ�Pg��4`���d)��k��_	��Y��z�����;@�v
+���+%Y*�Y14[!��� ��N��z(��я~t�	��j���I�0:�y�hJJq��0�@38Q��-���9�F;pMV$���DB[uP���,�%�L��Gς�2QI&�G�&������}ǅ+�{�2������y��4��[*wR�\�����I�V'�:�<�Vnw�q�$/�
��o&�*�@�\�{��{3{zI�&�D��d�2���'�.ty&���ҁY�u�)�dŽeb1!T���E�w�f�����	1x�i�e�:7�M��1�î��w�Ȳ�w��璙��YR�ַ�53,~0p��0a��v�#�EpU�pr���dH䃞�`�nɵ-�sB����wK��e�,�!Ә��� �P����l��	�"���a�{���/�\�R`�N@�� �0���^i��IV�Q�ʈ��<�fFك�x,��wu�hoJ�@XFo"F3��\2�'�]�s%�+����磤R��H�zR |��͛/>� ,3E�貔V�}�4��\�䀵
����I�v)e�&�H�q����ie���S���Z����P��*ai�(�`? D�Ȅ� l�f9)#?��w�x#t���5��X���k6(uS!g��$�J���X���~@c2t�g@��{B�`5�ıL�8b�j�Q��<h��6m���O���~��3�p�,���gC�ޑ{��@�7,�{�"Pdi�8�� ��g���F����8�F#����q�!�D�VV�#��aA��A�:�^��#|�E��BC�U6
%�%�� j=b�Lގ�fc��v�-��ǹ�؆��͹A7����=~	G��:� |���ޣ҄�j�0�vW�7�r%�sY95a�N�u��*��\��.�J�J	�픺l���J�fbq��u=v���iPf�k�u��s�9#t}�������P�<��2��������s�=FP�ɢ�s d�5���\���ʬ�	�� �`����������5�&y�8�Ir<	'�;N��=����H;7:��td<��;qT��Ǆ����e��´1e�A�|G2(��y�����[z�ߜ'���Ǆa�k�x�`D�(��ނ^	�h�
!��KY��r�D�$G�������A4z�=Iw��2^c�9`�|ꌗsD�� ��R�t�[��֋O;���E�}A����[9�m˥��c ��Ċf .������ۨTS�\jͤ��z���U�ͥ���j��R�6ݪ��ک�.��c�fsY��^S�7V�z}��j-�t�Sc)��J�TM�TB�贲�� > &L�ct���/كF?�yR�mW1a ��LP��bd�fň`j$����0��)���f�ê�P�� �b�ѠF?� <��t�g�m�E���a����ׅ��ѝ�Y�����,��5�r{?����[zP���_?�L���y'�9�Aa���rϵy������d�9�LX��!���_�F?��p�~؛Ǒ!�&���'�<ϼ�&H��p�$h3�.H9鷐&���N�T�ߍz�9��c�)��ฟvUl�C��o�d��;фd�M�z3W�X*�����J�Ԭ�{R�wn|�����MscS7�'&��T���6Y�ٮ�ʹS�\i�&J�63	�+�����ޣ�ssO*��=��nWm��U���j��J\�ԕ'F�$��\Q���?��Og��I�/��8AӑV���NZE:SV���w��Y �(p��>�:�VC�]B�Ыђ18����Q:���֋L�2z�/���(.�1M�ɐ"���m�l{�e�꿾`�C�*G ���w�Ű��ʄ�7��A��0<@�d&LPCꢎ����Ya�c�鉆pBU ���٣��,�~ �@v@�brv�&̱ڇz���ԍ���^��� ��7e�c`�����AYf=���r�|ݦM�^��L��0��#R/��*����oj��Vj����3c�2�l�w[+W�C{j��Y>v��욙�������l���}�n��YY�L?��灧����(��i���q����J�N3�6�r��A�A �+�8�!Q���vt��F�㊑ZQ�R��+NRq:h42��������t��R>@�c�"tQ��%�<;�2�RM���#��Rl]�y츑!Z����o����έ{�K�ee~�{�s�m��@AX��>�iX��,�\x> ��:wlìuF�D&��h�L&DT�$S/z%�����`)��S3p��})�3� 9"�Dz�1W2�0�)e��[.p�D�µ�b��X�QZ�m|؁pK+u2�e�-�j�����Z}nrrkk���[��k�+�];��� C���sL{����v�|Nm��?9>��G&���ƚ�R�MN��#h�0#�E������w &��$KQ��;V�
V���t�4ѫe5�R��</�	a'k�+�RcVC�%)�𷱿$>gԃcdIԝ�9v��,���<����@A�瓝Y/� �?�`��	�3�fT���E&,k\���sBNonX�h�1�@�a����)<��A �|��^{2���h6���Ɣj"Qq��;X9��0�&��M&�aÆ�O?��{c/5��a]W�8Ƌ>8�e3��TN��DjW&��Junz�����U_k�\���cn��导c1�*{��k�֤��k;����};�;���g-k6�[֛�sqGδ������R'�zr�Y�Z��7y�n�����1���*�#'��D���iH-����$,� �� �l�D�;����Aȴq�H���Ag�I6�:`��"���@eaN�EmW�Q[t'רC:��2�������v�(�Y���eT{>P��� L����'?9�6��N�pϨa� ��aϩg!;�͌���0�{�8^ ؊9����Fn�G����w�oQ��;�x�T����<��?�	�Q[R~�;�xE���eMxes����!�{��H�r+5R3U:ci��2ͦ�{VL�6�f�[��]��1kn��4�5䨿�D�����{w\���Ϙ��[1^n�N��J�VjW:�A^��,���8��	'��9�4^��R����j"|�۷��]�y>�0��D��J���غ�46Q0�h���,�`���t,�����Дy�A��=�fmٸ�Z,���ۿ=����]��g"K^�u�c��.�o�狃���<��|�8���\�B�a'ƬdQ�����`W䦀չ��kz��e<�4 L�.��zأm�u�V�G\5�g=��*:��qo~繹 <L�o8X���L�)C���}j1vd��k&t�&��67�sD��y��{D���.���Oz7�����p���So�;kd�4�\��j��i��>�N�vܳ~�����zm�?��/ݷ�وv�c/{׉+v=�S�������?eyj./��R�B��f.�xg"��Ĺ��t��Ǥ��>+���X.�fi,����H��ܔ+C�m�p ��  �Ah&=hPFm&���=o GM���T��I8��2�  ��"WL��F6�� t�I����l���΋�శ}8~�7x�g�,����3~����j.֐-F���ڪ� `eY7;�,� 4�5�19�Xr�m�\k!���>��e��c��q/z<�����(�T@�6����C���84D��I�e�<���LDr�����3�YP��>t��҄#I`��J�r�[���2nV�	�ҷKS��9�5=��o�?z��\��l�����4��������{�}I��/XU�?�֜��߲�I��zf�0��]&�0��t�G>�'$��Ս�8S<�9�L_7FL�.�/��Ĝ�ј�)���?��?�,���.ai�u��0�0����1�W����y�%�X�Łf1 ���C���!Vv�le>G����$.3e�! ,� 
�w�w�k��q�@X ��q�#�u���X^m,�v;�G�_�d� h��I{��/}i�&��	pрIlO�RJ�@�X&'m��<��B��2�,޹���t:��箾���<�IOZ�dµ[���vl}���C�0 �3�U�i�9���c���=�c;O\����E����Sˡ    IDATuO���g�����w���ܞ�k�Vfó��J-䈉�x�� �1I���K�v�ַ��uV;L�C��#s�7�1\:�
�$�"�������&��w�+殺�̘.���1�����}�p�ا��� v"ʮ����-/E���^*-ulb�&7Dͽ8��"G�Ar,2.�9)�"��f��d &�ꫯ��a�N8�	�_��_���ш����)��@��E�������ZFuv�.e/ًԦH��	�n�5��3�]2�'M��wd�`�Oo��Qn=������yQ��7(?��uѫ�F�\���͛_��'?y�bl�@\�L�����̊�U?�����w\���`�}Ҧ.�=p�oMn�����=O��'+�v֨����X*�K���Ǆ3�k¬�۽����.ơE�"�L��;'2��8�AV����a59�.$@�}��&���4��t�a,8@�$�u��`i� 1LV�N�*;n�$�����8�?G�T�81����O|"���Q��y��8]H@N&� s�pm[$��l��F�j!9�p#R<&b�4��T\%���s6��jχ'lzMm�� �a˖�3\���Nˀ�4!�'�F���d��U������?�R���96�E�V�}vÆ�}�S�z�blv�&|�^�~���1�Fy.'`o��Sg�q[��{�Gw�]s���z�m�)����+�����tѲ���c͙��R'5K�y&�E��?=99rX01���5BfE	�2{�����(�N�ڀ8��!�Æ��"󛱔�� 7 Lg�%"���Bg��$t@����7��ܗe� :PM�_��A�p�a�׏�.F������u5�{���|�DD `$��%�6_a+L�E��k-���Uc�vŤ��7֕2	�c[\C@D��w�7`��`�b��=J@�rp<�g>����lX��; �@F��,V�Nd�>�&#k
v�R���ƍ_w0@����c�s�p�6-k�֝��{�9q��z���nԇ_����ZsԶ��M�}׹��{l<�K�k����m��]��DG�Kt�**y�vޝ��|��&�F,S�9Y���@c������ʯ�J�<�){n?�:2\-:.�K�q��=0a�4sNx�X��v���\��\�t'6��	�vu9�b��R��b���������mʅ��>`	p�l�� `NbE��u�Ġa�F^l<&l���@*d5Rx��a#8�	'�'�&�]�;֏�� ��&�0���MS%�]=�kRâ#�?�  a����Rٖ��x>=Fۓ��n)R�0O�� ���/��u��~����Q��<uPm�+��Єg˕�_w����?;}�	��c�E���n1�{�M�NW�?�����w��̩V}Y�4����I���p��/��3���cn�@;;�Fvg09����d"֗s\ygG� l���ς�7,�侔A���PF:2�� V��z���5!G o8��/�����l����\������&lG��]����8]��O����*1ۈv��`��9`'��� ���Rmu���(��?+:�Sb$�ep���\ĳ�l�76�A�9S 4���3�F��`�7eP�Xj�� LY�YڌVN{��K6��L� ��\�n���l�0 ����]�nH����������2&x�
~�����۷^\�v�]�G�*�6S��]B]��4ӣN~T:��3�X���������ǚ�UG$؁U`$]ѭd('��e�'ٶ�`�%F���L��c�9	;����G�e�^G��xc7���J�e�Pf��06�}(�0H��8���a5�خ�\�Q�})�sr�:������N��8qE�Xǃ���; �$��cӡ�Wd
0�:� ��[̑A,9�n�),�KԌ��
���@Oe�����2p��;@��q��s�OAI��I�H�-A]����b�Z�qP�+��"gt��w��kq t,u��9�6p^E�W�s�R�37n|��1�Em���,�0�]�Zz`�q�O���n���_��Qz��9eӻ3q����ݵ�7�7gO�V�v��*�+�Jn�N:!��ſ��kci|l,5���j]]�����t؅Ҁ�vtB�	��N��g=+O�D�Mfg��}��N':�M]�T����ݡ�/���� 	�����$���;`QtD���#�-Ĳ�E���ܶ�2�DPv T�z?�C���	{ �� Y�20��F���E�=�A���u�Yy~ ;�z���xGdA�{l���2O��J̮I�)�ڪ��种aĬ�ע���I�r��B���Dw�(��+��Ю%/��mذ!/��_�lk��#y5�����O�9�x~�՚+�˟ްa�	�2L���X{��G�~n����o�C/�1������;Ϛ����V4�>�Rn�Z�.�M*�N'<��.��rs�T���z��#� ]���^0�=s�J��b3�Z��h)c��#G��e�E0.���_��.�!��+�`5,��ED��H�9l���ʈu�`HLb�"u��bp�]�]��n���^d\��@�+S�z!����ds�>�%�� f�2<!@�A�$P֫�>mړ6 �hK ���Cޠ]yw�Rcܱ=mM�<���x��F}p.�b����N,bC������g	��\��B
EG80�\�_~�<�>T2���y�	K�[�"��������=�3��=v�-��z�Rt��^�ɿ���[~k��[^����G�*�Z�=�J���d��M��	?rb:󬗤j��*$���f��r���KC���e��x���
`�A0J�2�	�+�As�	{� ���ɒ��눎�B�saU�J�ɽ`($����` �a��2E�Ƚ�Xb�/A��8�q�g�}��f�e8�m�Cu|�m H�h�<�̗�$܊�>�'[Vo'��m@���H7���w���Æ�x9�c[��@�bsM��͔���[@S2��|HD�@d��v�_<��7�$F9����IN��v��="�a�0w���;8�=�u.x+ō'��6dY%6�;�$�	\�1?�i��A�l�����+����@��91��y�c>=��Qn~��YhZ��'m�n����dٖ[/[37}R�2Smw�R���*>�7�H'������Zᩉ��nv'��v{>�A����LBi �u�d�z����,�
�-��he��	�z)�b�iuDϧ̰6�Z����T��6��(L�g��`��ι��cȖ�*?;�3�I��I��2���D�������$D� ~�^�=Wtw�`�\�kB,���"�]��U� );k ¬zd�מ�� °W��6x&�Źh�xI��sh�N'��=�kڦ*�I6԰9VJπ��EM�kEF���xuf�}��x�����xhw�8�����ڰa��L����}B��{����ǟt��xMw�C�z�5�Ԧo�q֪-��Κ�=?2V�)Ä�U�J*��S���ؓ�����Y�@�hu��;�C`��>2R*�	;Y�F+@�M\�'� G���9�s�F�� ���r��������\�9@�8Sadh��f�j{ ;��E|%�q}&��0�v�������E�+ھ��n`<�yœ�~aꌥ耰��;yw�F�$t��/�b �=�7���t�#���jK@��L�~͹N��,�/�2^刮u���|~���}D	�ߌv��&.�G�C�6�]{��0����b���mګ�Vh��W��a�]��kN�������M������~����7^ݲ����l�t���*ө1¥4Y���N>!�uΙ�����R��������D�B�U��#��QtⅲEw����7���_W>>׏�8~.��,�w9�spY��5�% LP?���� "�ᚬ,lqy�g&FW�]3"��@,��Eh�H*`����3��������, ��F$�����6n�-Ѿ�%>Äq�ѓiC�Y��xC�O.�0LM�g6O�A����,���n=em���>���q��'��O��T�2�~:L�L�v*��se����(Ca��1�uw�y����1�R3�aQkV�s����kl��c����~�c7������<���󸍟Z9���WOn���k�{���S�5��6Wf��&'��U�צg��ϤR��N:�Ĵlr*���lwC��H\��]��6�52B�#)�����t�x|�C�]+v��Y��;:'1���V�	���9�������6��� 9�DB����;�%>�%�ΚG�x8�0ug�u��8�s���۫V��N�2t�Q�G �� L�	_�"�ri�G�6�d�6�@�k��6��b�y��QF3�2������a���Mm�gs���c]x��z��uE�NC������hO��>�ܴS`��!����3����}n~��z	����ʭ7\�~��W�g�n���I����\J�j����c�g��������L%v};���n|��m[ߘ��e�S�z*7fR���J�R����������/����Dj�Y���E�*�a��
��#D�#��{a�t
2_ѱ�p�C/�r�O�C+Pv▉��;�0 Ё	Q�3"W�v��vG}��g�	����/oT�ڟ�^�sd[2E�ⲛ �v�	�c�|T�Q2�����I `r��	S ��O7��m3@��e���@ȵ����=��1��,,bGp�+��8pM�E��j�� '�%(�;.tr��fH@,>��y�������D!�C�0�h�K����
��6�'3E�"`�\�Z���_�t!jh�v\��	��@��Z�j�S�J�LuC��?:}Բ����,j��RT�3����*w�������dgv�T�����Tnv�7�6t���T�=�ݗ&''�o�Ư�����nTD���F�F��AX�(~�;'P����P���x̀����
H=D���Pnf�)�g���Â���0/_��R�C&���D��sd& <�	kqp;��;��j���y3���] 󐛁�u��~ G/	ǐw���c�##�g,�׊R��b�ݐ[�I��3���(_p'yv�KYB�r�w�Q;v~������}�h�E�1��z���Qtnq�2��ā��Bl���~Ll�T�@c�Z�N��Ax�ƍo\��7^�v��� <3τ��~�<��Ԗ��<��/׏>������~ ��s�����o��_��{ǅ�=;�9Ѯ�f=3aB�J�Z��ȧ\M��qg�Uӹ瞝�y�O�Nj�z�;����1�+���;��E ׵uFZ�HqcqAa����袟;� �Ɓ�c�0��U�ݠ'�iGaY���+��޸V8���; ���s�L��zǮ���A��G$t!2aT�`��?�Êڃ	S�)F�X�~�b�c9�,�XO��9�- ��}�ss��f��}��)�xM����jM��R� ��sb��A��#�0@�����e���}����"��������9�������3E���6����M�ް� <vˍ��ٶ��T�M�R+U��t�R%͕ʩ^kͭ\�O�cOx���1_��Mu����~��'/�}�'w�󋝙ݏK�4�棭z��]�N%�����t˖�R�\J/;���'��͹41�l> �  ��y��0�;@d�<"F�v�^d]	�h���^l'�W�2�8����K�,aP>�r�atb\�Q�4T���L���Cd�����!0���EX.@';Q��B˄s��b_���= as���xG ƞG�Y�����߂�e3l,��`ɮ/l �m�`	pAg��F�oT�+%6Wͩ�82Yȹ6�AqQ�����0��*):!�)N�.��/��{�֕OH4�8@��AC? ��c��{�ڻ�]�����N���V7�D�r'uj���Z��}ԉ�j�#�����q)*e�56m*�X{�s��|�-�����R�������ިݚaX0Ӫc���'�����87����f�����w�`x��4��|\DA��ȋ���p#iB�<���X`Gh Lg�?/u��ϻ��������bd�0�1�c��t5����3 �V8F�c�Ja�_�n��P��.�l@���o��
�r8����w�3��Q^�+�6��K|,@(�.L>��m�u5_�-F���W�qxs�.G(��<�9y��*�%�u�,�n/��A�Xy��+&�)3 N���R�0\l3 c�\����p@Y���i�Ub%�_�u��z��z?�L�+�n����۶]��5}T�<�zk�E���DoM�ԩ�ӞT�4W���1'�oj��?��i�൜�X�cN����s�+�����s{�����i�*��ޖ�r�������4��ؖ���ү��/�S~�������T��r�8p=�d#b"K�E�sa$�0l#f����0��lh��ha4*߹-����u�`	�8@P$J]�w���N�ŉ�~Unǖ���Z'/�R�	��9�C��d��T^B0���vڼy���/ �<Y�-��}�M�CzDX1vc��h�zbf5�q��=����a�������zl[%.]Xo��)#�xõ���ye����9 ��C<��;����q�xe�{��>Pd���6�&�LD䏃L|�Ŵ��F/�߽�D�����eC@��0�,�T� �ϲ;o�t����hͮ�g2��[ޭ���RJ�R'ͥj�WW�gc�1�8��{Ձmq?�2����o�8�z�֋V��E+ZӵJ��ʬSn��'���c���.u���8:�Fz�ǥ��n��f����Ra!�(3���� \ԋl@����߲#����1)��VL�=��8 j�"���� � �	#IP&�W4�Q@�q�Ƽ����c*up>L���fۑ������(�Q-h�HGqr�g��mڴ)�2���d¸� :� ��&�8��.S.z'�_��O�m�Uk~�{�.n��GD Ҵ#�y�l��[d�܇Հ���p��v��l`㑈p=nX���_"�������m�6('�}'!x,���(C�] s*�͛7�aɶ7z���;jj��oZ����Z՘>�S�)Gnj�rj |��4��33�������cW���\p�(F��c�������<�����wl��W5�{��TO9�|��:�	�%n/U���N'M��R�>�M��jtݤ6�]@Ɛ^��e����Fo'���0V/��wq�.v נ/��	�zq��� �!U�%h�<#:�0&A�c�dγ��I
�B��Aw�ו>��;���#�At.�lLP���>�腗���W�` ������h��!u�{n� ����Ł3���A5�Y�0n��,�d�X~���|t%\tã�CS�y��(\5ʻ�2�z0�D&\x�eH 1"����A62*Sv���>�<�F��\�h=t~��>pRe�7��s��Ww�M��Z�]�r�L��f��j*�}|���Tk;��]�͹G�'�=��;^��~^w]�7l��t�g�߽������_&K�&�i�!�d�x�>�l��Ff�,��Ɲ�q��1�9�>�H�+��ҹ�4�� �я�c�, �L�bXLܙ~���\����OC;�w�S�I�{�b�5v�CY���Z�r �&��:z4����;c�A�:�SP� laYx&HD֓��^H�_�3:VoF�6����w�!^#�Ɂ*��L�+tRz��XV �]H��9Q��F��
�Q��Y�{�6{�a���8���$[��/���x�ٜ��� N��%�����_���-7�κ�;^��5s<q©=;�0aA�=�J�r�-�Ӯ��={V��������>��k[�,����������2q����w�󧦧?ٜ��`���"W(;� ��w��<Jw�	�J7�%��l1�Wt��_�A0C��E�l)�1׈/��|3^��b����͡;6;	D�0 �s�j.�'���)2�����s2��[1Z�/����f��p2v�A���k�J�  �IDATtQ�!u����"��4�5f{��V�c�@l�5��kjkʆ 0�a둡GV�5�������`��s,:=K��đW /�d��=)c������%K����ౝ��^���m/\՜9�]�M�v=U�K��.WR�Y��N���s�D��k�jc����������f�66$�tC��M�R@v�"�&2J?ը��q*hq��GU�6?Z	!T�(M?�&�*�
��T�U�4���!�/0^���̽��9羳g��ݵw�����̽�|��9�y��u�4SH�^���]s���6�۾Y��\ɩ���_o럟8�.^xP�_��?����u��8���BKA �q�тf,;+��t�@|Ǫc$a�lȓDH�C1P� �������Z�� L�<���!#)��]k�׆.=�	�9b�G�y��#w ������Z�C��]�����[�TSDK��-��3��N	���#�7���I��[�:�A�.��~��F>(����o+�F~DŭF_�lJ ��?�j�C���<=|5�Cz�vp���P�����B	=8�SY��5�[3I��v���g���?�	�<cn��+[��=����:ώ6ϸ��P3Ƚ��6�`:����,��@��\ԛ�zN��ު���,����G�vKc�TV����f�>M\z�M|tW�^�� �c��u����C&)؂k
�v&o	[��XNF`R@��gu@�5�_��MGd���I�A���݈ &�x�� �6M� ���@���D-4R6�H4C�Ǯ~�^��	�A�a4B��$)�r4�$��E��o�k*�@G�^}�U����y�\k �A�W� �)@���I/�2�w�JI��m��,=P� o�7�s�<2r#�����>�.�G|	���0ʄ'���pA;F:=�oS��	!&�'���?ڷo��o�Z��Ov杧�?����3�^e�Yd����M�1%{�g�����3�gU�����~�7��w�wYe�_�rx6)�LM�p��or����1�llL�f���]��ӫ��z��LN�U����hvz4Lj�%�0$,��L'��T�I��'�� `��I���#�`R3I�؊��.�`�F�du�����#�L2�0|a����(Y��?���э�ɠh��&�FPG���b��cF9�� -� �>�`���/�0��� ��$y�-�݂W���n�s��'�A;��yi�`�A:a���6����3�`��Z�.�v�$�?��0<S���;T���qz9vA�3 c3�%�K�w-���������_�+��:K�0��d�G�qݹs��W����\$y�z`��;	$O�m�Hpɐ�A&��ix��sΦ�d�R)�a��
�t}���I9<���=�K1d����?���ĮQ��j�M�PZ�F�R�ګ5ZĪjU��Ԫ��R�����V5�ؔ�����γ�z�s�3]��p��i��L�0�zo�y)@TYfvf��LS"-zDm�0z�EJ�Ę�y0P^�3�����=s�C["	��sPD8#���ﾶ�|B�����o��'	w��
�	.�S�<r�qҟ!��&�Rf?i��	��\�Y�N�mO�	$v��ģ�bHj���qE�ʉX�T�($E~���8�kq��~��s��~��VǈQY0�<��wm�3n�*e(��!2Xp)W(^FYȏ�M���ڐ0z��(���1%��Zp�À&�N�[���U�rZ��1�Y-E����X�:�%����Aio��ޘc&��g�����w?Ek��8�-�6[����j�1����?6ٞjW+E��M��q�F�I�6���F2�����D�< ��D?��������+)��n8E�	*�������V�m*����2/��}���$Q�� �+!���6h�I�5?E,�qI�Ʊ�6�:e���� Ì䠀u.n(=�f.oZ�*��ڌ��tZ�O��.x�*uS�ʩdKҔx+��$��ðc����:�ԸK�,��M� \����5(��k����wh�l��h�m��"�Κ-�Sڱ/�G�,{}!����;�~���T]��q��\���o�X!rB�:A~AǮ�w�ґ~k�D�"%ᭉl�4Ց[�<����3�XGP���:��[<��|^�8;�0�&g�7�K��8��B�w�n���aEߝey>�o4��v��%��4D�e�~Ʊ��?Ӿ�CM�5y��w�k�3�����d��%�G�o�=d�;���I��<�G N���v��<������0n�S����'� j���"�C~�Ñϓ(�<�+m�z���{@I���pY��9�qʇ
�#��O|n!�}�T"[��*yy�Z3�g�f�
����<��>�!Y�CF�����&Gk�sX�yy-®����2vW?-�ʁ����g���,x/F0��H��"Ax�Qu�����?�R-��p[�<���1�\�Քۡn�G�f�d�%���{�𞙅aF i��qee��#7� ��3��׏7���;$��iX�z}:��`�����LuB��?���<��("���y_���[9��ED��\�P��Q_!H���I���B-���M�B3jf�={�F,�7j�I�6	)�8�_V����>[����wkZiͨ+D3#�0��0���o��?��y�Ʃ7����?�?�:�>_��~�����Wn�J$����-�y�w-�U�!7�=�K���62���U�f��7	���	��I|���*,-�\eF�I�G��Q��x�銃� ���}�tW�B�� я�<�.s�վԣZ0y;�pE1��±G]�x~�s��duF1�T7�N\P�����K*�d�5H5��{���៏�d'O>���͎���xr�&�{�կ�B�;]Iwȷ�*{���Nŭ? Ѧ�Y�6���5Ɩ���Z�g�n�M���d��������̈́�+���]�&Fܣ3��ȝ����\��m�����J%�7�N.V^���lOI�W`��Ԛ�;��rFM�hO��&kSkwK�F�d*�=���e�yU�2J�~��s�<�<�m$�ȁb��A����F�1$�JCzG�9�0�X��=@��L\j��nl�˓�7��d��4�̈́���=E@���Y�����Y_ވ�o��N?�vҖ#b	�
�{�� %�R�o�l��u�i3����7�( �0_#G����W:�z�F�I�Sh�_���Ĵ-k	y�E����uh|�wrn�I���K]���+ԥU)�~��J�M��h:��,���0XyO0a��W�m����m�	i[p��������b�w,wk�n�i���2���|Q�aӿcOd�����ޟܟaP[_�BV!�,��
���I��ʠ�5W� �>���O1*��T��C�".C��±�$��&�^�o,k���`>������b�=`"���r�ʼ�"���T����n��րj�����B�������!�������Ѧ���C����I�ǯ���>ZHc�K�V��
�;	�`"���X
���/�����$�Ďv,�[��5�8��f!�-F�[i^�G��b�#�ۣBb?B�/_ɋݭК�Gb��xI�ݩ+��@0Z0c��]X�)��"����lps�lU֩ʑV
�&,��焾��;�E��sx�g�k���=���qH��/z	B�=���@�!7l���������Y��K��WCNC]�����:�0�w��0����ɻ	�%�e�4��()��c��+iY��l!{8� �j���%�&�Z0��ә�<���Pf��36?�[�z0�M�?���x~[�੓I[*�" ���.�$z��Y��f!1����>�g���D��UgΔ��2%z_�ֹ�\
���82�~Mg�kTZo�%s1�ˑ������ݣNw-��)k1��o�Z�F&WК����D���i�5j��W���r�mEwm;�u�`��IP����P㕗~��Ka����B0�A�q&�>B.���0בTI4K�� �i�?�R��1u�03<ԏX�7�˂%'�mj�9h���^����ivJ��A�P�4R�m^���P�MݸY��� 	3�ܩ��^	���E1�5� ��$q��lJ�O_&64��%*�����b���G��O�w��;�����F8P��cfpBiN�-1R<0#-p"ϲ���R��,���a�F��IO�sd���e3����I�F�]&�N��74}$x{L��*۸9��ԃsNVق>����{6�k�9�2���[չ��y�0�H�e�UKGd�V�)��
�?�R�:���l���<XIZ����l�j����A�h���r�W��y�8�X�;��쎈~�)S�v�O!��ێ}. �B���t&�Y��)zG�A�2y�Ÿ�3y�`�
��PeuW��.�id�sĻ���r������!?j�6�#ي�V��}�;�v��#7� �eqe=��q-MgDbc�,����<�=��]79r˫2���x3�ȧP=���}���u#AQ+��|��CQ}�Qűq�E���Ȳ� V.Y`�F4���w��o��{@���x>��	t�@h��;KmO+K�ҷR+��6,.��+2c��A����-r	��Y�����WZ,c�����2�*���1ۤJp�����h�J�������Z@�8�/ILM�����W�#�'�����J�|����q��ٱtǀ���Ϸ9��wW�wB�B�lk?%���������Κ�ꨭ5 �_R�F��Ԯ}�3�"��'?�2�S�t���(>����Ν�O��\��p2Z����4h~{{��8Z>��#@�Πu�Π�S0�.���sF	Pԭ��d��H��=��PX��x�v��o9q���="�J��[P����{ǭ����;o���NՄ�6��.��mE�������Ҩ(���<�պ�?	~�W�-e-6.�$���ɋFaZZ���?Ǜ������cU���!r��鐵�����ʗ;^';0i9fI���i=XI��ɝ���:��^�\�n�{7��>Ԋk�����>�;��Z_���0�7(penHV�3�Sx:�Ҹo�<��{@A�4�t,r�A���hqb�&�au=��S��
��.��E!��;\�(l
R�Tݖ�V�^�h����Qt{J�~aulM1��Z�'�}��:��~ϝz���I��`�ϊ<O�.��GS�؜��i���{�k��	�;�j���\�Դڹ�,`��>}M�=;?֘����D�bZ��"��V�aH=��ov��,w�pn�ө�o�Q�+�/?$U䴐�^��g�:ںf�c�j��д^�w'2�_�&.F�m8�z=E�T��|�����^�*`���r��.H|):�F0�ޟ��_�2���2B;���P�D�	��3�'y̭]]CGmIR�����B�|v^�=�}	�߯��5��M}�XI���n���2�S��ToO����ޖ��_E����KPɸ����Im���ˊp���D�l�"G�,cC_���G���)��ui|ۯ�u4�Q@N��)j��3�7zœu
���hPۋ������|�q-#&�1E�vK��/j�ET
#���A멃�,*-^�!��GA��T*u�*��+�6�6PŁ���\e4�Ҕd���x益�������m��Bj"�7.��̗m71�!��U����;<��o�]�K˰�u������������񏯣�S��FB��tC�_WW/鳇Z_� Ps��k�Ѝ��x �����ö�nv@9��s.ƒ�d�������%��V�C"��Y��n�qX�6�G�?��n���$>�z�c��,� �WF�.��}1�{����
W�+g�VK�Kb��6����w:Z�%�Ko\(�[�s���������2��=��($T���.q��hB�@3%��]d��a~~GIɿ$�Y����������k�*�[?Ceg�3��rƔ2��v���ގTڵ`�M�oOl��PK   �X ���s� �� /   images/6c5cc51a-5517-43f0-84ba-83f8b91107c4.png��csfMۅ�ؚL�m��Ęضm'WlOl۶��m�zs?������zwUW��{�u�3\^N   HJ�(  �  h64����|Y�� c'��  ���$Q#�  __�"��n��0��j�d�9��ʁ�F��V�#u7�5�ƣn��50��n�?�cm$�?���.��=~����t��&a�̀����3x��e#d���I��H��+j��ʼ�W���\������U�|Y����1J���0j<K��=���&�9�7����<��K�QA��-B!�[d��p�+e�c�n����뀿��T��!?d�� *8�[����_q?��LPW��'���Yx�w`W��X��ꈴw~��E��m6�Q��V�ņ�Wߌ�m����x(≥��\�Q3����ʻ�ӌ��f�p	v�AU�rn���ŷ�%�1�)���'��%a�sO��U���rӶӹ�p��"��w�ʽױ�{xj�㋼4�(��4���n��c�7eu�P�K��p���hv��{�Z�����q'���20}�_gk�3�F'9_����.*[G�6��j)IH9�X|nR�:�?��0!�@��G���B��i��M�R '	3���Elh�X]	�qӢ�����+����&jqy(>��=���������Ų�1"�����1�~��%�]0���N5>,�Oǩ�K�\���`n �2���P����b��m��[8��X�3��f&8����4]���UH<��xa+������0Ӈ�5e�e�B��Is��>�����AT���W�mK\��}=C��ie�)�>��ee+aM|�i�K=`���OrƵ���O>*$:9ݭ8����)!l��g�S`�:U��j�,�균����o/<KNj܊�}����t��� x[�nɤ�Zr�[a�}{�b�q'(��W���O0z�n�0��� ����tᗵ�B��
4ɑx\�^9"��:}�_��IH:)��۽B�{o:sN��u��XZ:o<��4����׾��I�0�M0���B|�k�y���0��p�<����X?|�g��T����&��9k��}�lb�F����d�t��2�;T��v��C���`U�:�8w[-#O%>��N![��}5O)�e۪�-'f��4*=���ƺ�~O<���X�����(�1T 4p͏���2v�*�icd�x�S�����U���|��k��z���K,�Z�4����q���_�Jqk�������6=��c��{�
=\D�fƃ��p;�u���e<D�$���7��\E� U�6�ll��-l{Y���DG���ц���@�Q�%�o��z�hNOd OlVw\��W*��B��NF�A�~��qv��h�����ĺ�px��L}n^r�>��RC.�֏���l>|�!lZsI?J�rn2||s�jlo:?j|� ��g��2%_��v�|li$(�7�J�\�6���6��z��~�|��n�9��W{_X�J��9����;k����,�Y꼚i�;�؈����s�&5�O��=��L)2dx��ϑv�Kk��+�>!��d��W��?r+����
��L`gQa:a�� SYֵ����b&m�D�0L���V'\D� 7�T|T
����J/����%�'v�xڅQ�G�I��d�"]����}4��}�c�}��X�Ք��(��]�E^�D]��f�V�|a�충g�#��^��F��m�mg��1����Y�G�����}���ږ������˴�'�c7��c�9Ρ��H�����^ T�q�����
�h}�݄ł�j�ȅ�TiT`M�U��&Z��r�;e�1�*��{�^@j�#% �ψ'�$wcT�l�)9,߻��L�'�"i�K�D �Om��ǝ�j�l���r��`��[ru˰|���g����\�Q�y��cQ*
�3�_��V}u�Y������-"��4���������J�h4bb�r������f�-S��e��&�46hW<��u_g�����M!�E5�c)�T�t����NOx.��1�YL��������܂�� ��V(0�6F�
�K�n�Ov/�X�cPCP�rrb�u���[��l����1H;nE?#a��s��*��������q��ULQ-s'������y����rСsr>�B#�uUK��i�}~ֈ�?N�B��πgN�u?dd-"�%���̥��[A6%W	C�	�����Cm�	�/��Ⓨ�Z���5v��#��9�v�7_��&0�i�2b�bNP1��M<`�v%��>�!4~��9|�'�n�p?���T�$k�~�/�Q�L��v���G�� �VK�����e��*�c�S&ډf�Q�F���.��iZ	[������+#���Fn7���|����.��w�^7��ziM@-G�W=�'���D�?�& ,�uMu	�q�v��>}L�|���6\�>z�|��=�Z��݊�����n�?w������m���3�Uv��)3\	���t�՞��Ѥ���d��N$!#��TvO�9�JP����F��E�G��w��V >�!7����y&п똌Ҝ� 1u�v���EDm]qL2Z����揾���3|V�U�m�Ax�ɡZ�<�%�<�R��d۾�b�p���W����*[�4u�S@����Ll;!"H;/��.d���b m���ֽ-*؋��W|9<�cL���A����H�p�v��Qkc��[�t�����4a�n�_.�6k4Ń�6NZ�����w�Ӏ�j�I*��]YD�G ܓȗ�	LO3Z13i�oJA��-�����MX~?7b�aW�u��i:���.��<ls���U����y4���'���B�vy�n��������7�P�bP�3W�}�[�K�-
3G��z�Q���V=��|56-Ż5:�I%D����1�I��Oc;���4����!Մ��a��XBWW��(ˠ�I|�siq��gkcc\KK�R5avV�T����i1B�T�PЎ�Bs���z��ζ����Tp� ��J�|�PK��J�gX1��h'V͞A+	t�u���W�k�ழ~����I�,��%K5��ړ�F�+���U�+���\{٧Y��p�O�����	�F{5⎊sv�gG���э�&�~7���|5zle�k�g$M(�{J��YRu�	F0�d��`5�*n-�.��:]�dY�K�X�`�U�?�B�E�����<��yV�h�U���X���XM�e��dI��rz�����O<$�rjk!���Wi0�1@cu�]*+t�u�x�d8?���؁�Mõ�z�U��w��{1�t�]�؀vC�o���kʒޖY��ԓKOSk��[떸�ʴ�M��$�PH�B��SI��/�<?�޲��w�ƀ����6[�_U�]qk8	���P�wq��k�[��½�Sv7z�Ǟҍ��q��Qp��$���g�d����Y��3u��鱦�4�T��gDY�����nL��cy�Ƥi�C�U��]���2r���1TeeM���G�pz�^i�%o����3ꅣ
��@"�|L�W���E�Q'�f�N����81qpp�}�=u�Y�>�����gq��w]u�d�v�z~}~xs�O�0vi�S��vd�/��xv>mjv��|O[7�̪�!��wE1f�Ē����ڱ<�����*
��+�A�sA�յ����R��Q8��d3!���s?�21"FE,���1����H��FbV�+T�~5��(�^Ey���ў�33B�Js��Єܿ5lR����gw�;N�A�$M0<x���
��4-��Q����Kͦ�ߝ+U���&�m���&R� 3�Ӕ�2�-�.�����W��f���$�"Y������"��݁� =�;��I>�}(F ~�!+$$�c���ʴ�j���u��q��j�p(,//�,oM����oʖ����ߌK��lq�!��"U8��E�C�n�~�B�i,5�z�C��X��m�^��럣`LP���_�%�/��9|ԡ:�v�U�?8qp��BkW���\��e�����>n[Z��5'��S����Ҥ[����.���rqݴ��S��m�?�N�Z-V��:��5`ٓ/�,oA��4���wƨVW:U4����cFk�"ۏ�C1n��y��e�h��Y����t���hs��OEL�����ZRjA)��cӰ�����~�uf$}�[8�T�m��P��>9?g���I {؅F��dm�a�c�4�N[���+�%�|dB��L� �͑u�9f�֝�����Vtr��ӓϣ��4ԁ���o����i)�U��3��*�Z�z�3����U�dǴ	9>4d9֑?�o�L%�ڎ(Z���ɺ����W,�\��Έ�_L��g��/��4�&_�7��ӌ�܀�β�@�a7#+������5�9���7\]]�{���:��|�u���|?_�����^��d֢m�kvޖ�]7���{�|j��<Jx���Q�q�^&���XV�RљH'�)IOCԣm�GdQwE����4�Х`���l�5���s?��2�q��$��w~���5��Xż)~��m�!u8��/$�TFu�qx�o �3�U*D1�jPf�#��Q�"K�<u�߀�q�� �>̮�;�c�u���B�.�4-S�萍
'���ς�c�qvj�vm�aw=��Udnԓ�̈́3)c�D��ڛ�xa�Yq�ŷ��,��n�>u��2ʸ5;IL4�L4�j�9�(-�x^X�l�w�LFDMO���e��&d�6���,�����}J�G�>t�:0jy<���iW��^��pMN�}D�5��S��6r��s�;:�����3i���k#CˉM=��2j�����	��Efv�j�<鸍�O����wX�V/�z��X� �� ʹ��Ҟ�S;�l�.CG^~�m!J�O�V�^��!z���&���H �u�Oz��Z��o�����0�^$�#)�:A�;$����Y��0���8�r��<)���iM�r�S���Ӥ��2}��.x��������
��K�e?���'��Ξ}83^��xz�mga�vj?�F �i�m���o\li+�}�a��^?q�c�uы��>��c| زj��=a<c��T�[���e#1�O���V�X�75gP��b���� �8=;�T	C����f`��;E�S��.�����r.�2N_�6�_�C�_�
�`!}������xR��H�ӂL��gT�b��>.�h���{b�Z��&R1�t�|lso� �?��>��C7*Z�O�p�	.G����a���#L�F��Go˚�:�Y(s�kxXvx]���]����ܦ�!Y~|���{�Xk�YF<�V-�J�*ǉ%&6�i��������mN�'ot�?��5�т��Ƈ��,�^�^�����ٔcImQ�Ah���Qm��0'������Lo!����E����/E}��v�z52%��RS~���g���"G/�j<*<�L#.��䤓���䝴{mja��o�O�n�l5�,ЛB˰�@\i0O��I������h�c x��)��$��\����?���I�vqro�C8�Ä�c�Nf�\��TS�|e�UC��.7�|+|�5
���3E�5�H�I%�"9�N2�j6�zX�lZ}�<�j2m�S�F�����6��'����uT���I�ک�ge��(��1lC��M#C��JN���e�f�_�OJ&���{�韔�Ih���Vc�y��i�ꔀ����I��J=���n�]���ݮ��g�6�Qna}��k��<&����s�د�h�@�Ql���ʼj�9ʍ;I����z;�K�r��F'���;V��,�#�����2��ˎ� �CiA�6D)؟f��FZ���	��'�V����q��\\a�E�9�&T8�_j&�B�����6�^����Q%s�-����e�F�ލH�G���O}�9U3��c���-��չ��`2�<d^�F �L�j���*U>��Y9��� ;�l�8~p�-�^o����F>~3���|8%ι��WW��ҫX�t���%� M��!���J�AZ�(�����0�_sCݩ#��T.QȦ f?�OcUA���Hw+�ι�W����*M��Ad�K���jH~+�aQ�G9f���!��N����D�`���e�Y��|��%�Q�d��
n�>\Y
�J�AY|���]�п�U�_��G����m���kX,���!�{�����&_��@�$�Μ0l�њ��eSS�c�GN���.��!e�~���c�����:��{Q�"��G���V����w�M[���uk:������!�NV>O!k��O�4B)�?���߲?����%�@Jg�����fU�62��(QT�\;�r%���MЉ�P�28[(���-P��S�;����Ȩ��L}i�Y^S�	Ɔ�J$[I�V����+1`�^|� ���L�Lؤ󹬓ެ�	W�?c��g�Oy��Zm¶Nߪ;��wB�BР�����/�Q?΃�J14�5h�~sA���X�
��e��Ƭ{�VT���9����\ƫ#�v�r����_�h�a�7���i�J�ƎE���FU�-�L)�9�
k/�Ǫ�.>�U{�y�� �ޞ� �o>$�����d����P��5K�1g��2ef ��NjE=�
.�5�MIi��ۃ������)��{�CM$;d�}r�@�w���xi�ʂY3�A����@*�#E�"W�&�b5�y��D�f|R�>m��I*{�b\<�]U�*%�VR��bV�g��_x�]k�"�@���@5�� U�q6!+�%	ۧ/,=�D�|�%���z\!_'^4Q�j�>�c%\(����.=�ǡ10�n[ˁss�Oo+�X��f�$hƤ�������U��5��|��M�V7ý�	�p#R?�ߕ���t'!i���p
���u�?G��S���j��S�B�q�zd@�����f[��a�HQb���_C3��'2�����+X���ze�����'$XiK���ďf�a��z-��}&]��ύ��P���~Wb��̓�hT�q�J7#�?'ޒ�'U�x�4lپ�$ʁZ0���<{1Z�z�s~p/o�z���NL!��6��q�\����E�����2 �n|3\d��d��O&��]|�A��Iqο�b��^�u<���"��?f+�h�c0�=Z��]B������9��ٱɎͶ�h�\k�*��?��Kg]~<��w��-�p��~�郘�C���.mêyq'��� �矒~-��<7��#q0���I���*]�a2�����$����T�M��Ha�H}��Ր�WjvL���p15�Ux
���&M~G�칇��Q�(]Q��I(�˴�_y}�[.7�]�D��|�,'�� ��+�}? ���S��=��n��|�L������s4��)�**�����7����ͤvv�����8��f�.��gF�%Nh�,<뤠�%H�J�rH�$d�
�V}��M�+gn����ϣe�ӇW�C�� ��[c���	x'��)�˨\i�հ�=���!M$I.iI���qu��͢����:?B�ͫ�����nt� �ԟ<)��֓�	��(~��.ڿ�^���|ޒL�tmJ��xz�� ^E�� ����zez3!�Sgu�¦4J��Uc��y������cvF��/�_�o|O�kF����)���;��m+9R�I^�Y�Ύ�����~��Q勧�6m'EH����0ޗ���%ن gJ?����<��|���oN2�׭1���cSΥ>fAU�Ϝ��->K�Җ�l��s�~����4�zc�]����o����5������6�Nwqc��a����6�f.P o�E���v�K����{�f�`���*�ϣ7e����Dg��t�]Z�x����ChY�gc�ᶝg��	P+H��p�d�0_��f�ع�k-�H�oŗ_�_�:ʨ���]]��c
Ά���̭d�K�̂(����W�I�d	��*-���W�M¸�޳{�ۊ�3M4j�y
����y�.���\��l��k�i�W�����A��q�BAh芓���.�fq࠰�5�^���0>�F=��5��W���{���ش"s�$*�τ�"�����T�����d8��!������:kW���}��y����ޟ�2�� ,�Ap�[iu4��G`�h�pɨӮ1(!��ф���(�e[��Jx:�H9��Z�U�on����Q��u#O�Y5}���Y�������O|���\xi�2�V�/m�sFg��J��0�8�x(ݾ˶�O��Z�2�oD⽟y��~\Q�}[]�<ݸ�y�8��$���NH?$l���P|�7��U19p���=��)�R��O.��Æ���)��:U���:̨N�g���s��w��!P�o[&Z�Y	V6� �uT6�ϖ�/�p�h"�D�b�q�6t|0ZoG�)H���@�6M�x5eUM�q~X�IrC�J&^���D'w<#q�KZ���1_�ԚMV��{C�3hH��Zޞ�t�>�l�&�x]7ݏL+@@-ɸәt���o���>����O8��PI�B�'	�l~�[ƛ�;6��L�1�,�'y�A�?w)�"���I˟ڑ����f���+Ձރܷ֝}�Ib{u���?��2{��"��7�|�uӡ/B��7������j�z�0����t���9��-�q�}�������i�L��t^^�?���r��zA�7�����&�{����A�RU�nTU%�h����Ϻ�£�Y��̆x{��_R�:!�}\��^�m�ao���ČM��v��<:������i�"�p��	�a��}��`���o�E$�$�T�r=�@�T[Od�ݴ�p/z�����:�1�roMR;Hj8&*���>�/ѹ�`�>��s�X������l����r�@Z�fռ�w9��铮�E=ѥ=�d��}��@U�F���W:5����#���t[���FJ��KKz�/V��}�T�҉PO[��	�A����9B��ղϩ0x�_0Sr����K��!��4Q�jeN���7U4�o��Y��p�a{=��X�AH����"����?�c�4�>�]90Be�͉S �/�-�x����v�eG��wm�f�w�%J4�⟭��Q$��k΍�P�r�CZ���c���L�m3�1�x��9��t��z/�V� �<�/E�3ly�c�F.�?8	b�}P+�B��M��J+R�
�4��6�=(����@�!%e��+ߴ��s��J@���DwIK��Z��0{Ja��[�,��迷��J�'Q��w��g3c�E�1������I+��ϳ%�7�\P��6q�K�ͫo$�R���^Pdi�*kPQ��l>&�c�CB�*�=���c^�J��5��P�\�
E|	����I�L��<��C$ ��!#�qQ+I�&J�C��4;:��,@��[�7"p+?����!�w{�w��<YV����Q[�@��r�	�Co�W�<�*y�ls�M͢�M%Va��
�~}�q��Љ``�7_}?�8h����'�C)�=R���&O�SۊϞ�	?��������2��2~L/ńT�Y�WΌ{�ɸ���eЉ�E\%q�BA���
,�/��3������K�C��*�fv!̛5r�!��D�/�#�QM�2QX��*3�۹���.����;���dP}_ߴ�M���=���@��_���s��}.�u�$MRdH��>A��ndn6���Q�.���)oF9�o8+���K�H2�Mށ/ވ��tL���ť4��W��q~Lf�E��-8i,�0c����
�2�y}� ��$h�d�Wa�����A��7�!9��jW��ڴ �S�g�L�;���05�{�-��X��#��b��+������ ��
�ԂYv@�q>!�3^�@�U�q(K�a��=�e�1r�&yGr��@�5�c6���p�(�
�ll�u�A��8١�[�?�ZA/6�>�5��Ť���f:E/p��RZ�bGe7���0
r���=~C*�-�^�`EH.񼹴T<��#,�"�p�R foR��a7ty�(�*���+Il�¹o�b��S��f�����l���0jا5��\�J�s2t��H�N�(�/�6�h'~�M��x�u�X�j��W���i7\D	h(�+Z5^����Q�rRE��:�p>q+����E\q��0f,��gG��9� &RP����I���p���{�(}�c�H��ˮ�-� P��H���*ж\";�;�[�(wb�S9�F谽"ݷ�A?�hx4��Ҵ���J~,tM�S����$�K
`�F�X�A���B���m��$M&��,�X��sa9!Ǽn�j		QL�ٓ����w��C2��);;;��{&=���2�﵋`�l�F��U�]�pI�!�f.6L�r'��'��Pۃ �%��)z�|"h`j���B5�����h�-�@����6#hF�G��ʄh�5��q�KL΢S2��1�U�Z�.Z��b����X/�2��a�i�M��^��8`��}Uk��Wg��jU#��#�P5k���p�+1�����h�oy5d珕Q��=��*�/��ZOȍ�wr�+�nD_w��-^C���X����r�ٓ�F���a�U���[^�d�0�E���k�n
�p�j�C���Z�Ժ_a�Z�4t��h6�8��6Yl��>7p�S*�p���G���k$3P&DݦT���z��]���Pe8�Z4�xF7�P'�h�`Zͦ�%�|�����T7���:�V�ˁ"%!  ��UHV 9X~���.����MGP$� ���0���B�b�U����8�)3�-��T�^��5j^\�$ݤC��d�T�v�s
I��`?a0�L��:�f�]�*U�j^��̼ ��㞚f�� �#�[��XE����O8Z.�Z��������!p5��+�%3.�Y���gn�����)�q�n��k>�x����/I�
����e�?����+���C-*�������~p~c?Z���
����-|,�Eü����X��7�v�`�t��6]�/��9V��f��܉�l���t�<T+��Ƌ��&Dɂ����ۋb�G�u�
�؎�hNy�:-->�r��9����װ��N�ςZ��	mJ|ޓ��DA~nmy�M�Mre�S[�o�#+���>���W�I�Y�p<������BK�={�cܯ��(��p��v��%0��c�-Ww��C�A�K��X����́�H���X�5ݤ8�<Hѭ��?]{�t���-�p��v�Ł��9��t�V�� �7�(���FlNFC�2�v�QQm�-�f&��ơ��"vJ�=O=�,�9{gx1igJ ���zƠ�)A7H����d��6�R8�����2b�D�
-�?��Q�3�~��&��g;�XΚ8~�a����(�8�Oc�7h��P�p �ˏ�.D`t9mV���V�� ����A�������F˃o6QՃ���	��t��@b�:~�~�CO�_���:Gz����Ď��������郣O���z��c�m��;��z[ ��n�@�B���sܔc���Y���s���JH^�Yy��l��!t���A���jh�j���JQ��vo��ISTR��_7�}�'g\Bu�y��
�fz�!ڪ�2�l1Tg%��wx �'�T�:  �K��'!�^��֌L���H-V�V�_�F�H	(fFtF����8e1D����6��#�&���<�ޥ/��.����X�-���m�l=�e->^n���i�v������f�_ h�����oAr�=�n��|^xK�J	�?XX<�aL�#�5`�(Ƿk��_��Oo�$���6� ��(� �Jź��U�YU�k=��<~�6I!�kvh=���ӥ\eDx$v���]o*/t����ol���.2���@��U�jm�d�!�ϛgվ�mk}���g���<�у ���q�v{�^#���[���3A���u�_|P��U7� (�m&A\J��5��u`+�..�^̕��S�Ӧg�%;*�4܍�:ձ��� Ȕ�8Kђk*ۿ�wD�bF����¼⠀1G/f��Ŵu
�6uU��)�^��+�+τH�5C������� �_l�4"�㸃�6�Q��V�	wqq�i݆�?];��{ +:t�ږJOo�t�ژ֞��>n3�_2^�zF���N@�U+��8��bV�*�A����d=�@�1��;�.̜��f�9Xd�{�*�:��H�Qg�	Az��6��%h@�?�.VB�$���C����1/I�S$�gf�=
Jr�y���ƞZC�n�\}��1ܓ�
��V�*]��m|V��i�.N�nTT��v�W��&@�ƙ��H� �U�P��Ȥ~�褠6O��km�P �Qm��گ����[�� �����l=ʆ�G�ձZe����b�%36��
u��N��{f,ʍxg$Jc+���+u�
Z�2�b�Z����Gǹ���7�)^ ���)�UG�,�_#V̧�5�ȴ
:U�]%DB�v@��`T��n���ǩM�u~�E���ώ!��ǰ���wؾ�@��{�8I����"�Σn�h��G{��8�O#X�,��&J�t��W�����y1�p	�Q�#��ːF?�6�9Ӈ��"�#D����8�Z�Q����]`��n�
/#f}0N����rب�h���R&�fP�$ ��T7��7[7|�:~�dl���)��T��_"�P�sVL|H	K��ٳzX&�0^���M��0�S_�ް櫧�D*��,��1�E���wj��̈́�>�e)<�I�@��B�����L6����wؑ+�љq	�
�2��mQ}/�7$��G�[0��^��~�kW�#�}8�� :�m� =$�߀>-�k�J!_S�#�h,���wh fL���1αx�lXG3������ҹRֹ�>�����u7G�E�e::���o���u���W/�����	��x���ۅыu�(M�TN��3E��q�qϾ��p��6\р���1�}H��*O_Z ��L�5�ڢ�\��ُy}zL��u�1��b�0�I�8;3��D��n��]}��~�7;HΔf���7�*�=U�W�]
����.���錸�d������g~FK��céը2͂�_Ũ��P߸
 (�!����0���>z�|���=��!�XC�k��f0^�ҳ�I�,���`�5�����[��C]�Ab7�L��'x�jYh�����-7�ӛ%r3�9[�!b�N8M�̫�ؒ���r�������i�Mv�.�Sa@z�!�Q*.V"�N���O�Ѩ��} >�gS�H�r>v�����IR�ӎp��q[W�J�R������UYNO�A+� %��eڱ�3@�1���W�Κ�����VJ��(-�����xD���U������ڃ��l��"N�Fb�_MՌ%v�줄fp9=ĺ��;ed9�l��X��}?!�:�p��0�HQ�� v^�K(e���ᇏ�������Ǎ-���x�96������T0�6v��a�&���j��a${�<�4ן��XK��8��+ȴ�܉4� ]�:��ѻ]���}D�z	[iIۂ���sYhUyY�|;fT�@*�Јѣ�օP�]t�M�'��u.(/\�E���A�/���7p�!�����Y�Z#�CM���ue$�b�X�63up=�b�i4��AY�5��|�9�p��6ēsj}6��z��U�,���;F���0Ǹ��C�9�����ioX�휯��E
˳ML�ï_0.�|�/�M�~���@�	��s��Kpd��"B_pk�j�=8" p�:-�$R�@oG@$�ʚ��U�q9��P�  ��~��hlr4do��R����0V��Q�넯��<�85��wl��`����Ɣ��.���7���s��%EG�ȵ�j�G-�><8��ǂ��ˀE��f�}Mx�}�  Yvj���l�t�4�㠸��}P�U�yk���W�G���E� ��y���Hn�׈����BZ���C�`"*���ϝ)iv�D��v(,]Vt�l�)�n�JQDjBwx��_���<�	#H�nWMQ�=w�}$�� ;�,mR����������w�Y<����,��1�*0J�J��H8P�Ը�Bc!�X�#Q�z�@�>}\�%zǟ�'&q&�t:P��q�*�7�ԠS�lV/3��-�%��.P�����C`��t&/4��i�8Q�P�u.e���u�l��q*8S��z�GY��F1�M���$�&�{�����׊~]�!��|��ou�DF�6�eд�����v��R�3{P�:R�����M;��#H���WXKW����x�1Jԉ< ��=���dm��C�2��U-�+����h=:��N��
'�LQ�/	�'-�~� s�ѣ�k��.�N������C-�����4ʞG+!�5گ��1E.�c�:*�"B��#%�4��=jQ��%�A��n�³�c��/������Xm�MPT�CD?Ȁ����A�k��ʑ���.1�"Q#�
�Y��[�.Ɩ�Ո@	�R��2D���R@9�Zy����F2�DA~�,$�6�c3��촟Z�~��
���d��ㄻ�M՛"�?�~�:�w�b"�x(�$�	������K $���7Zϴ�ynP5�.d�����9�E�0O6i<�����GB{s��cqft���:oa�+B&&��>EJ�A��9���p�,p*�0|��?�ƺ��G��04ɝ�nHG��
�ϐ�[<���Ź�I
�U�5D�k��e���!�����#0���f!P��h�U��K�xTo{����_�m���>Y��v��݉��w;U���Aw�Q����@�{@�@��V�[i��=������q�:�Y(FNM +�مq{+7��_��Q�<���-5?Pa��k�hdv����Q��k���|I��6�� ��TƟ���ؠJ����򹊩�@�L�`�������V�G��]"$�	7-lQ�{q?
ZUβm������רu=�PS�%qs5�?BA�մ$f@�Z�Bq☘4)�:)�sK�0ȝx٘�BY����"T�5#��bDe<�f���]�N� _��1�Ed��=�Τme]��ńV7�	�h�z?d_��t�}r}�~�4@�<�i�t�R7u�
�\��]�F��������P�p�a�1y�'	?���W<��ş�qb�H�~Њ+�#��tf����!�+6��8K�����5vG��L��|S���T,�f=��I|L��u��j.��U	&��5ƛĄ���K�][�L��&���p7$o\�Sc��̸��c�o�P��uy��=��4$i��>z�����^��Itv�6�}�ҿ��/ֿ����d��J�Kq�"K���������F��ݪ��$����2�{�q��~�2Q�=~s�o������ r[�ڥ]�q�X�oG���{e�XNn8M��uJ�?�tcyi�v�oO��¹�z���}��ٔ��V���i��0��i����OhE�b2�9����q<wM�d*J��"W�6L������~��AH���V��7d!S��=\]AlO�|ތ��V�-C~������v1tI�g���m�4,�I_*��DЩ��J>�<����v^�x��k;�a�`m��q�~JQ{/��YX�3�����.�d�)�w�y�m�Y�����n{;ץP/[`*�j�e�[dͬ��n߃�P�I�[��J9ل�"4^�Δ�V1a$~�y:�!tل^�+�G}O�����VBઊ1D��6�<��_�rImjα��Z�6�2���s��d����08�� ������Ao3�xv�g�{���R떩��k�H��<���Uc�*�[��G����mF���T���V��HǮ���]���X�Iۧk��,�D,�����2ӫG���x�f' �{���phRF�纎�V�����4ܣ>�����y�e�%~�h�#J�B��w��dd�$0m/����Q�:~d
|I�ꯘ-%��E(r;{�vϼʹUA�����v2�j�%�tdεrVD}�w\�P��m�O̲9��������+l��4O4����).A�O�ʨ2�d�V�����%���)��͔�@�a��W����V���т������O��J���C@���H�GF�ʰ_����X9�����/� ��,�ݲ�28�yڗ���ř�?���������DEsg��N�9M�Y�l&�VD��Cv�K.�Jl��
�Oei���gK���tS웞�I;���a����Qc��M��ҩ���厛&�
�as?�d���	Nd�N�vi�Y�0��A��J
�?\A'��������;26����;���p�tW�f
o�B&��Dɮ���](����J�-7�)�,]&o��*�Vk�o~Ov��+a �o��Q����*I���W�v+��&9xK% l�L@ �c}�E������N�6���L�a?�P���lU�dǵ�52+�΂p��s���s���f�463�,TX�d��;JA�7��:�y��S˪�eJ:�%e�xf~T�s�/�.7��!_L�b��J�1W��P��o}P����NUdd�!]��$T�����ؾ���[Cz�zd�hU��?}K��/�NB��%-���e3��dGcE<�K]բ��Xq�����
�����6_FY戮Vcx���,>eW�PWؿ���/٫�Vה~�7&ܶ��Y�����~}���v=[4љ��Qe�I����x!��%QU$zaO_ᢉN}�;��2��o�����Gb+N�ͬj�����hM*]�$|�T4��l���X5
r����
ul[!�wr��G�e3��9JqI�&/�@Ǎ��U�Pp��7�3���n��O�Oy�;A�2yb�ؙȚ��� 2��P+/
�L��j���6-����g�QR�����9l=��v o&;�.6�I.�����8��%OB5$��̸ה����s��&�D��bK��$S���ׅI�|�$9��gZ��T#�MC�]�TV;�s��L�2��&j���3�*��%+�
��{�9
�$R� e�p��6�m����,V&9I
,����A�Uw�i��3��Ǚ<�,��C��eoۼ����&����7������c[?l���;�Y���5�-�2�d�'H�z�Y8a�j�)�ЧE��4���(Y�/`p��L�/ۿ߰���|�f�̉�o�ެ���h�8n������*+��`��F
���
��k�S��̪.���O<�-�j4��틚�Bݵ�Z����������D��1�݊��ZU�Vz�)���3}ie̵����Gu�,V�g��:�5s`fE�B$4�^�7� ���<W�9

����?�X*�nAd�W4��l(Qb���Slv�\�G&����D�'�a��d>Ɋ	@���q���X"}��$�π��]#]�i�ifK��zC�jQ�j����/�}��:f�(������Ѱ���4��Fi���n�đzb�H�GN]�fu���~6^�=*�dql`m�N!���ѾS鄓��y��!jՆ��Y�tg�Ս���0�y1�H-g�da<�j�ڵK�0�}CdόH�C6
��8��e���l[�[��%�x���k�a%�7�R*�4�(VaO�x	*y�S#��Jʄ����d'��V�{��} ��%��zRcp ��K��fN~�nҏ�4yPRU#)�4��+�X�ȉ��u���� �v��e�H�i@@�ߋR)�h�a�(���,�T�� h��2��?L"g����y�)8�������� �"2�ae���?Fr0�Mg��:���@K_c�-���x���1�+���>�Y��x���a��R�<��(��>�r!I�������R�m۶i*K 1];�S�z`�A�8�#-!��3�A�I .΅�"hp4"�q��=;|�ˎ��0������~c�|�JAǂ{��+��_E�S���0��c:b�V��1SN>��|rKs%Բ�'A��ۅ��Gsa���u��$S��Q,c��(�o{ �ɺ���������.d�kR�J�&�* <�W֬]�+I�T�Y�e:�N��6Lą����49� �7�t���J;���I�6H2��x�
���l٢yG ���q�NpEf5`�ܑ���p��\ԈfYKm�93�p��Y	��[��V� �0���A�i,�<l�
��C�j�bH���D;ܘ:�h�ΔL��4�������������c�DQ��	q�r�~s�a�<��%�Mo�\آ�7r�,\��;��cTǅ�1��;'�oN��%>�N�dOl6S����8]KN�SsS]-)���i��?����SH"�#X"�Ѩ�#F놲|����4�Zo2.JW�����SU�Q�*�
(/ѿO�e���Zo����X���C������?�����,�d����N�����Brx 0���&�s�� �6lP����5XU�"bsu�	��Hb��T�qR7)QT2�pT<8��Wi�`��������Y�eX,bڡ�x�k_����.���j쏥������yC��]� �u��cB��P�z�pH^�j��?�fy�:y�O}Ɯ�,����D��G�AlݺE6�y�a�k�I;&���-n��<$���+�V��ɌVӕqN�Ľ��%*��W�xq¼�H��O~_��H�
�C���[eϋ(1�0��eX�[��+��qҭ \m�һd���i�݋�a�~l�TO��o�,U���~�µW�8V�� �}�k�����`mJ/�㔪P|�����Pc �.��'f0�0���Pc�҈��l�����0G]
���|��s���8�%?�D�
���ZY"q�h�0ox���V۲ap 0J]#y�\����Z�!�g��i�J�u+��f�������xg,1�אѡR*�Jo���3f@�W�W`:o�T���?W����]2<tD
�b��j�>��P���XW�f0P3?����f9n�9�d�n	��9X��K����s�>��7� _� H�նo�A3���yC|y����Γf貔���19|��3�ʥ���A�b��.��K.Q�
5�����Z����K�@LLw�xu�ʀQPa��ΦƤ�b;�(�3�_y�zl\�#S�� �h�'�ö׋��nh|�%	�	�7Ζl8[gB�da>�.t=hVN@ðq�/����P��-oy��p�z��䤑M�n�lT��E���n�]�xܑ/<CN[{�T�jR�c�2&=�>	¢�A��w���$g8����^��hr9�%��#��NH�qQft��.��Z��J�]��ǂ�<Os^pS}p¾]g���s���]ق��Aw�]�Y��5	#�T��_��������37](=}+e���%�sE��Di��D����*���7�Q���p�
��&�^�O�N&f�>q k�@�Ŵ  vu���0��ׅ���،�f|��ya��R�to81�
����v^0g;���1�`���K����R��
2b�ep����s}���	�~pTc@lc�Y��KSy2:,���o�CG�w\w�|��~P���Uw�-[P��S0��]m�!�/j`�����5�r�I��(@�����c���5'����QvfLD��ᩤ	�%��6��d��~>��d��Ȁe;�f�
	WW���b�D(�Ұ�;�U�����|�w�I^}�:�$n���:2��1B�';T����'� ��xF��o|C3�x���cB�L��+-���4�j3^���s�9G���.�/񼸨n�q%3љW.xիe�V���͢��Au ��2�=�VFZ=q�`�X*@O�

�y�# �����1��� �=�EB�C��&�r�3v�z�/ˮÆ�#׾��r�Ƴ�H�\�=�R�%����*�&�M7��?�>�cϑ��X�~!��Z�Ɯ���L�)�SK�|��3��ɖ�4�C����$66PR��(�hE��|*��'�#C��� ��������o���$\Q���B�%m�F�9X�|�f��gT�|vK"F}0� ���C���j�ꆁ�Z dۥUki���QË��0 j+ �m�]gc����0�#D��GG�sww�,�]jf?T.}	����&�B#��J�̐K6&����� U4uv��^`� o4�u�E)(��`QEóL	�aG�Ql�j�բ�9G]�
�ɞ���W�R(��q�v�0`s^YC>���F(�rA�"��Ss��2�R3$���F��o�'ʼ�� ���V�?��@��/��� I��]� \N�1*���֌����<E=�4�����_)Fz��PS�����N8r�5o��V����~����2��GU`�����) _���f׈㱁'�_i�L��k�E�8p>X�~�NJ4��ڌ4�m������zG@�~\r<m$���u��S�݆	�c��ƺ񼯶���C���vyp��1C�AXN��6=�e�#H�9n���`��=�Z <���F��$U���h���իW�c��_UU\x��rҼÚ3*'��4��1���m��ҩ>�^I��7�Y��̘�4OE��(�N_+�����^Q���,�*�d���:>��
⌗%S�5�A'�|4��+��B��?���`��ַ�>���W�E��:^ ,Vʬ����	3���������ň�^���o�G�Ŏ�B�2Ci��P�HB�CC�T�uȆP��#�^�3o������6"�p\g^,;`�c��g��n���m�Ш,�d�-f�p�GI�RW�}Ǖr��uf�#f�n$���<z9�!mCL.���%�񔵬BC[OOY�v��r�]�I�5�4&�=��i�3#`�
�&|V*�R5P����w�m��,�l4H���"�5l�>�� p�+b�R�����a�TI���+gd��{�n�u;Y7�0xtl�f�p�+�&�rF����l���0�lR�,�	І \�6��a	�G����+2�z-��5E�Y��=��i�z�5[^�.Eؾo�R�a)[�H,訙�r}o./s�mFiƒV$B.�J�,�l�X>�W!�����w�������a�:�I�/pF{���p��+u ߫��Zə���L��u�8�]��.�i{Eثvb�]�3��ZT�;n��av��f�d�t�޽gwa&r��s��!60c����KVb��	t>X�}��j��1z�3�ZSt9a�8�l0�x���L��k�&kVwK�ё�ډF���U��w�j v��\rɅv��h]B��a��H&���W�z�&9p�jƴ!l^��ƀk�*X@�c�Ft�}Y-dpI�� �|���U�7���M]/�����`a%�&��z`K�P�.��L��8�N^!6�0c�ho���%/�̉�����C�>�3o�G6k3P���8#��f�t	ܴ��Q��.�@����/�J�;�S�>h�d�Ri�hJV7��Oh�=/Ԥ�1�kʂ0��D��U�ȴk�I.��,6���!���c0�oɀǲk�a�f|�1y(�+A\��K�Ы9�%�&Ԣ�H8dU�v?�3�~��o���b#F(1�0���hP&�5p�2���`/�ʳ�C�'T�����̰�l�A��۱=NB�"�v��.v��e���
ɰb�e8�<�����m	�m�C�d�� t�p��<%�����;��N?��׿��e$62�����3�f�.�8�!��;����Zal��e��r���xE�D����9�����$���1|ė={�����ʿ��0@\It�KVʅ��L6l�,�jA��T��	�1�`E�m�ZWo+�(`��#�ZU�(�*#�@����/�O�Se� k����A= �
B�0�wbڝ�{L�>�1��X�Cg����Q丵�/�Ӥ=H���i7|�Sdͩ����v�B������22[l�9TS4
|�q��)�/lU�*h�x@sV����W=0ddT�R�����k*g7;zNϡ�2�z���{�,)���dd�%ʽ[oאK�)�z�Itù��r��a�a�xH8f:8jخY����1g�UW��zVv�8"Q �.Þ_H��bdT��.��	CM� � 緼�M�w�K1��f`�ƍ��g�����4M.��{�,@*D�­1��< )	&���`b���1���]
ޭ�֧%S�@�q���5�46<�����Q�W���iz>���'b�`���@��D�!��@��Q n���xȀ��׽N�?�|M������w�yg�˂�Y>L>�l_G�(P��Ǝ�&~�	{w�'G[��I%Yg����r��bѩH���c#����#��`��}��zV��L`G�B�a��ˠ��/�\1*	�{�W0䫮z�zI ����؏!�XM�}�ٺ��k�y��3]Ѩ"a� �
j�B�rg$�Ŗ�����W���a&�)Kr��ae�o��W4�-"�1h0�0���m�f��@( �3�T���x���q,Ap|���~�#�aψ£��A6��j�v������M1�tH��}�谖zA� ��A��9 ~�J��\��j"����� "߬$R,��f�r�[����%W	Md ��{����1z��3�Q<A���J� �
 @�E�[F�# �XK��X���Z�� j�0#Ѓ j�'Ӌ�4�[�*�xܡ��ry��u�}����I�q�K��0U�/]>(��|��iш�1��64*��P�c{�xA�ш�1�ne���́m�5�|���Z��m�{��#���Tmd\JT'C��K_#KJ����J�����{�O?�9��iL�	�{G�KS�	M���e=����͐�-j�� h�#�[jcCK�s�Ӵ�fm>�I�'���'O�'*K0h؞zz���茡� ��ؙiob p� `#	��h̳�d��c�j,�+o�\R0��EѬ�x��	 CK�(A&qs7�x����4�%t/�@4
@I��x��2�)l6����l��m�+N���ַ�_��_u6�;�� �i����m<���MA�v�5]��W֟�/���R�nؿ����zc�lT���@��K./S�ll1jۙղ?"�#��ϕ��/5�-�Zݗ�%�dhDd�Hu����%Mx�[(��N�8�˞k@ژl�bF�Q��>�W��W�{���El!#F�3�[L� !�*$�O`â������r�2%������)���Z��n����Q�)4 �?�p�P5п��@���ҵ��I�[�:�K�3-S�Q���I�c��M�����5������w�*�x�2��WF��(��1;ʄ
��
"�\�B*�]�t9R�*pT<�R��0��g��R.��z�e��f�4��Be<	�e��Z��|�{���!���R�� G��2P��f5�[n�E-��#�T����nE"��(��W�?2d�A[S��xއD�Rr���& L�\�ׅՑمpcL���7�$P%@����K�.�m�&�=C������N�n�mG�	������n����\�����~�=I�;�&Œ+a�O?�t;izG���\���}�q��D����O��/ɑ��a���/�B)$KZ����a��1�RK���$�$\d��![�1o�!h� �Pi[X/��+j�t�������F���4@8����Փ��F��t�F��(�=�ܣ���p�`��t�t�̺q���g�Zb�b�v���
�\��������O�o�2y�������T^Օr���Q��� ���AF8�2�`¹�R��x��Ы:�P��ȑ1�η(O?�O�9o��
��QU�Y�J	p��G�3)����%I��	!���{�fDw�$�D�	�� -A�o&i��JX�]԰-s���m��(��t�����#L����F�����Ibv�#��IC'�r&�a�N�v @B�wG�@;����'& 3���3�����y[���;�1�Z=���4T���!����3��G���p��cN+�%�s���(��
�� %@HT߈Q�H��=���o�A�8��B�*w�X-�4��G�=�EŜ[�h����e&ۡ'�"@�`l7��x��A�q��-�o��D���t��'�5�ˊ��VR�l$	��P�	�	�V;C~z��4�����!�M'^����%S^��G�=�xiE�$e+�:Z�\���hM��ukd��^��	�F2+k�'4:��xE�"���\G��	-�M����)yAM���a)���c>{�OFd����_��F1��;�D��h�U�H�^I��m�I��u,��b�h<���`��,��[ u�+�x;���ΤF�i��m~�#�:,ms7�RLg���Sh=���Ͳ�6�O�lp���.�ț��Z9}�Js�5e�����ۼVPȓF��rѺt,����%cY�r���(w�����0���+H���t����a�Q�
ؖV�7������*�e���k8���m�4 ��m����i'������
Ϳy�������W_$�>_F���oH�kn�%%Y�AA]��¹��2]7K��g����Uv|�����V�%�Ε�����=�<%�m0+��`<�KO�Ig�
�)h�iE�:I�l�j�6���,�-��`ʻmwޅ`��9����Y���r�\w�I{���kd`�82:�G�{��F@Å�HZ��UU��Ē�ͽ$ryy�L�B��s�(��q�h.n��W�s��^s� w�X���a�}�[8����
3�b!d*�k�UO�U��pڗ�H@p�}@a���YҨ��&���hp4/tɮ���ޗ�S��}���+�'}��_;��b�X�#inkʼs���*���o�`�R���3$�>�TʮV$�`��nCnP��W�zz*j�����X,5UIƴ��I:n���$��L��|�$l��C���eɁ&U�hؤ/?���Q� ��G�J��%w��7f����J϶ *�\r9f��T��������/_�Ï"��z�R����.����H�>f��"�_xN0G�1\ՌN�Jq>e:㺵Js���)��Ubs�l!@��jvA>Ɔ#���5�����ȣ�J����+���74K�����D',	�p'�c8�8'¹��2�N؝��Xj���Q��P��[��CU9rpL#��9u�iV�������Q-�nV��Ɛ�m ��u[U���e��j'��Pf���L8.��G=��[�k�B��;�=�Tn.s]6W�G��U���=*cպ��`44ܐr�Wg�(4������)��șq./_It��JQr�a�%�u�ZS��4�;�P� v����n� �u;�-��خ��v�9[��h�ߵ��>w�I��LY�PD��$�,l$��+4��&J�-�I��pa���Q&L�l�윞�R��J����2:��˨��<�s2u��C��X�A����eI��3�_�¥c�Xv��oZ�dfq��S��d�K�z	Cfs.����
^B�ό���O�r14���{��J�Ud����s�շ��a�F�s&c�d)C�u�L�Ê��b�[&�aUb k�� ˀ.������z킟�1�EG�d��$���a��1{zz�Z}̀n =�.xhHZϭ�՜�ņFBR�(~G�
�Ff8�^D
��l��j�T;п��!8/R�m۶��}�X͆-� �cr�%�ȩ+��/c�vH
^Yv??,���#AL�k'�aU�\���[�	���<(x���m���_s����(�����JWπ����@���$w�nB����Gi����d���$��l Z�s3�Ta�c��8����-xEl���W���6�+�0�u��o1��3a���&��PNA�4\���(�(�2�#�rc�b�ID�����d(�<�c,�^���L��kց�I}���=��v�{v��Y�j�,]f�����e���X�W�è���!륯p���2�U\�9Qn�w͊�e��+e��k��2#��,�{�"8�l� �w<I�kV���s�	��I�ƒ��E6��DJ\֤c}8V� p�եy�H��w(���cH��c��"��� =/����$?�b'���E;˄����:�:�r����~
h�,�����9���N�c�[�7��;��s�g����Td3_;��L�3����s;>,6 ��m��dQ1�����|�;?�姊\y�y�Uꑣ���<ui�m�M������Aƽ%�s��\���
�7 ����i��C>b��3r�+6��ҵZ�hp`�2������Wj��昧j�Ł��^�n���oЂ�x������T�A�3���F�!���r�RG^x���e�&� �ׯ_/7n�ԙO<��w�}
�L��4���0���.��eH?WR����ޛ[z����Y�K�}E��,�UHB�Y�&���ej��$q2���d<N��$�q9�	�+�8,�)��n��lV�f�EK��u���Ϲ����{���,��=}�{��Y����w�+��x1�����ԧ>�0av:���ݽ�,(=̗]��{�2�=I�u�<��:9��9dÂ2�d�����`�u	|F��]�I������ҭ�}N�շ�b�W�SZ �����56PE-�k<L�n?ŭ����LZ<:H�ƽ����|��7��[���q3����t�g���n:vl13�L�23^�2��U�y[�l��:�x�С��]Ď
̴w����Jԃ	�b��|!��`1��Lވ=���ݟ��g�b�A���1�y��:��p�ȌwRQC�; ���W_�����%5��vJ�U/� Tt `L�|�/{���������Ed�2Z�������M8�ߙ�]q�tF�s�F��4�ޕn�w)���>�^�ꗦ=yw�͢�5҄�6ƻ^1F��~������=>6���o���{aW�0:rd9}�K��y4��}n:�A��Uu���@�Y�0�5��0w�za ���//�-�+l5�ھ��o-Y}-��|�W8R8C\��XU�n8U�w�W b�
��`Zވ��q��B�TuG��d�3���b�W\�b�B'���Zn�����+��F��1�bԀ#�]�a�9�
�dԏ�D��3ϝ�nF�#��i���Ӓ��V�6G����#���=�Kg��V���r5t�u�J��ԛۮ���%������u�f6"��jf��↶��F����%(������{~nO"���)������!zW�L)���^��������Zv�.Y�^ı�_�����fS�hZ]j�=צ
�R��O}j�'~_�3��ߜ&�\cm�
 .���.�����P`[r^ r��{��ǘ/�݉�s�}hV�P���k�413:">�q��Lci�%[�	O�y`�=x`!�����w�tɥ�(;�m?��T�^�P]5��_i���"��On���V���[�A:ppoY(`��$���bj�T�r����`�a,�{�����׿>�����9sPi~��/�(��z`p@�<N�9F�� �O�g �#<ª��ک�� �:a�Ӛ,hְ�o~�bE���������Y ZU�_��إxO)w/��ӹ7�x�D�s�e��7��嚟��g� V'lֵ뷊� ��j��28�<7;H��ޖ�>��~�^�'P?�:�i�5̬??�p!��$�ο͢S�-K.��1���[�Sth\��}����y4@F?m��ڧz��rQ���vjYԪԹ�"vI��F��4�8��L7-�׿���;��a������j���4�5J����Mb h�8�=I�UJ�ˆ��R�N�Yi��S�?%D���h3��*N~��wx_�)p��7��#��qb�y�0����T�h'l9 �w} :���x4�-�-�8�-��~����78DQ�?�y�+�Cf�!�}�����ɶ�K��H���_������M/y�3�����_�UE��'C�U#�;���m.ޗ^"�lKL��;n�N�h���X�Dd�n������T��g����\��Y?�T5~B��������矕�ߟ��|� EY�̆���I>p�#�-O�w���~����{�-	�N9C�DL?ap�ȹ�Pe�u T�j'�JǞ]�I |�q�� VQ��j�Ӣ��6[#
����J�{��Ep����=g � K�U��P������b{�7�]��r]�Q�����¹0���������ƸX�^�i*��p9��k^�Ͻ7ʹ3+~�<8{R#��=��H�J"�VI�<U���$b��[d��h=K44r���T�	&��]<z�ȸ������v�"������n�yN6Rg���؎��/��@3-.U���>Et�ra����*��!w�|�+�}�J	 }��^W�v�3k�H���Z*�b<� ��wU1�.�<&�%�h���[ �ƹ  �����������[�R���� ޣ> ���}���RA���*2�XE���y���<�$��KGsM ��y��P:��a7b `ٺ�hԏ/zD�VTX�,��XZ^z ���I���X������{�M�Z�8o ���/"ب(&��bM��m�yy.&o6'�);�`����[�IVϹ�eO�ux�=�N�� &��4���L����a/}�ۇ
�Y\^���@"�e�f�\�>V�N��M|u-Q���i<#����+��+��ha� 3��,�b�DW�6d�u�yX�ϫ�W4*y�5br0>7�x%�Vq���ye�~{�l��t�ܗ!|�H�´���d\��bu=�N����C��DM!0�.���v$�Gv籜���ă����u_��O�E:�A��]�b�L>W�@{�(r$��%Q� %jy��K�V��ʸ����E]�j�0T5�*��=M5����I����C��Oг�Qi��Y�}���p��jYXN]j�5g�����@��}��<�������ԧ��g��IOf���	�B��B� ��x	s� >��a����// Ѹ��_��_M��dòZ�$K�i���un�cP��u�߰^ū`��5��'-�@�a#:%G�ca����]E}���g�C���9�������i����.�@�f�
��`��ǃ�q�tǝG������ئR@+���#�	��E��䩨� ����ϝ%��z������"Fa�EdZ���u�ұa��i�}��Q��jUE�#n�ކ��M���`���@:� �Ġ����N_���Ro8�v��W���Z�J��5�m٩�8!�vQ?j8CB�s��$aF�I81V!��=���ʈ�bU�-%�9SU��t�[2a���1��;�t�X��JS��aEݬ��q���*������s?�sE����u����I7L��9 !�z���q�U�5h��ǎ.�ߙ�T(�D,/̏4d�͉��N5U'�!�
�'篛�����T9�хq� 6�kâ�@A����n��i���zl5W�ˣ�l:�o���}�53�f��i��+u{��U%s0 ���s}����%����__t�	� ^��/�B���K_��d=�*+s�|1߃8��*=u2�zL�w����T	�����fba~��0&x��߰LK ���/ܴ"1/:��A;Oe9a�Oy�Sʵ�h�r8\�{BC�=G����c�V���y9;w_a���ZNS��}[IeY�n35ơ��;�!a߸Kc������x={_3<�Z���?��	�vr!��>��p;�&s��0�ۿ�_��0��]��G{i���+���t�y&\������'�u-�p�*6a�Q?|�_,ċ(]���[��������19�	Ŕ4M,溚V�^���o�h͆���j��R�#3wX����������V�\X�5�!��%�_��&��:��"2��`��À�d�X75��XIaȷ�r�:�4�2p:�n�����b��G�s�:����k�]�9������/�M:t?.xc_�̊[�,�dq�2�<=����L�i����y��18�tD#��_c��Q� QU$kv����Ltth�5.zi�&��w��=�L��6S���XF�@���a�xhu���UWѥ��t���$}������w6��ką��&k"\7�֫�G����R[�w�1|ٙ��xo��g��y��c
� �|��a<�V~W��.~���RZ��I׿�����D������kj_:t�r���嵚�d!���R&;�ɜ0��}��������da�>D�џ����xЪ���b�c."	j�S"�?d̮9��\�:΃m��a��i��= �k�
h?��9�Fg�ܕO(:��sh����u��Iv��`���>|���$�G'� �)�n�p��x��_]������c_����{
�}֞�g�{ݖ��]�Ϧ�G�������q�S&:��V)-]�p|��8X�N& �7T��G����*0���,��~LT�i��B�A}����P�'i�L�{=>TU�QF�`��p�İ�hP@���gU/���	N����9�*MP�|���Q�V/��-���;�s��ϣ���B6E���e���ܳ)5����s�-H��<����@#�qv�H��;3Y�휛n�클w��|?���᠚�s��
��b_��hyȚ}e�-9�����8��:"��+[UltWaɟ����٫S�
��0r�1���c��K�诺�:b0(;(*�Fw5��3������Lam_��m���{'l��N+�M�/
 �VIgG�'�k��==' ��Qrq���:�I�Ȼ���=�%�N/}�uU&���|�_|�+�
�K�V�\���aqY��|���	�eE���=�š�Ɂ|�^���|�P�[6����~ٲ#:c�����S�]�)�9�ދL32Q�aLQ�u����q�J��#�T�yd�V_�Y�z�D�d?:�K.<w��7,A<J~e�5ת��kՃ�di� ��IdA?�d�3Οh�	� �5�'��1�W��x�H��習���;��u^c��kj!�3c��0����qǹޜ�(j4�o<�)
xUn.���д��է}�[[,%%�$��F����cc�N��a\H��^͋��΢��b�˼�E�/��n�_��0��.�@B�I�p.�n�ݜs�M硎` `����?��q�9�~��	 ��3�w��?������w|/���ki�����x�̍˸���p�*�{@�G�υ(D?�@�L��������6�}d�ѵOp��h��Ah�4Y�b~+7(��5Cb���	�Q�$0{?.n��D�n����5Q̶��'?���JUo�%���M�׍ȹ%<�����_�ӯ.��q������� nbq#s�� 7A��im�0[4r���Gy�U�����O}6����p��x�cӹ�<�����d����_�&m>_�SЇ��<�����@U'@�o�1@���ߙ�V���{^�_ԅ`��h�h�9U�bK��r��
��Ro�Q����93]����	(?���"�
]���O �u��7�u�v�s�5��l&9�'���an�=�9E���6l�Gü Wf�L�t�Э�ܜ^��Wd����n��(�bW-3qq���l4� �lP�0h2w�v�;��0�3گ�GH�=/}���t#�n8NP�;>cK�^9�qa�Ff�y��
�W��2�"G�vL;% �G��q�,�MH��8u�)����5"��ܜ<FՖ��(mE�瀯h0�*/��>c�37P����p^���OfU$l���Yn�;����,U�;��̀��S��?���L���� �H�3{��oHވ̀��Zq�g&ܠI"�wr6��C�;�L i.�p��Z�7S�!�W�}�1�Ҝ(�ɑFh4�K�Q���Ǆ�����ԙ�&ʰ�ȳ�FH�������9(�n4��X����R����\�1H�΄��Q���
 �~���0,7B��$N�i�w�f�4�.��QZY��zG��G�^���Q	Ψ�q%jn���ˮ����7�'�('��G?g�&��)�9�A
pH �}��|0�H�'Rt��.:���rl�L6&㤟�`6���`4�����S}�s�0>��0|��F7�� �|�����I�B��'HMH��ؐd�qSQ�%{�) C@���Z.���/�'j07�>ᚑ�sN�ec^k�+�����=��}�	r��n��e%�Fȋg�3���X���^��X��T��d���֓m�R�;@������R�mi~�=Q!��.�t����VW�\�j7��h�q#a���H+lB?#�b��ߌɾ�O$k )�1`��r3�|�K�.k�����i���=��	�pY��qb��Z$7��}�U?_��xy��ޛӏ��C'`���V^���O��ѿ��22u�V\U��.�-�.5���#�o��]�1?��47ߩvw\�y@�����]|K��Z�Zd�47��X#��%�3��cq�|8�`��=��b���5�y=@�	���sr=�'��1n&61�}��pO^܇@��`� ��K��T�6�,����*�(F��l�8�RB,�8��3D��碿8 ���>�*��d!r� Td��C�ٍ����FgF=;cʼ�xv��k�q�A�����Z��@|]��+7����^釾aL7�i����y���u�hlr|��V\c�H�ֵh�%�0������-_�tZ^9��W�TV�Ro��O%-�Š2�>��������L�N���$b�c�}�ܠ����\��܏���S棛�7��������4���Ä�P{ǖ]v,B��8=3��;@�A1؉�Z���� 8<��� L�2��������X��L�]�RGk�ĐBrZL�ѱt���k_���o?U<�٬�y�\|���xK����c��+�s��Y 0A<;;����d�y�(3��Ȩ��::`�o�0��bԡ�W'Ɏ�(e�dt�������E��Z�z ��4��� � '9�x�\�  	�`��Y����8��XO�7��H�ȸ7�ɴ� ��/�ʋq�1�[�+�2^�J�^\����Fk�Uf)���z�2q>4�,�v���M�f�,}�Z�J����l&|��������D���jc�(���u���^���7�Iǎ�*n��3.4Y�_cCl��h�`�C�����9��l|�w���*PؠKQ�<2n�ĺ��2/�|�Ӏ���uPI4OGe|�h\�����a��Cgk}&�{x ��i@Y���q~ݓ\�.VZd/��5�e�F �<��n�X�巼8]x������4���.�;+7"sX��D#���a��g�0� ��A �=@�Ŀyo Qt�t�@�
:��d<����u�q�0q����@�_���7@������)++��α�ȸ��m��c��
��: 'ǨnBtw�	�	�@̧Ap]�	аy���>�=�T��{�ч,n���o,Z��A
r�`�m�9�
�G�c��&2�ڜ�{��$����w6#E�`4P�M��J-�M���dW��#1���m��7��1F7S	W��O�Of��
4�:�t��OM���_������ݗ�^N�),���3�ɿM�յD8�$9Gy�����$��x�zt���s�����%��8�W�	c�ԤD�9"f�~��eW9�v���'��ڤ1�&�L��Jv��]}��.R��04���N� �N�\����H��ufK3��dYJGg �<#�kp0�1u�<��[�d��hX1����So̱.>����j� ñ���KF��FR-� � E�n:>���cf�WU-<L1\�~���Y ���L AF
�D77�Q��T8��D��F]8��Y@�X� �̒��&�Qm{���g�"�2H��	�P��Fù ^���D#z谈�
��G>�w>3/�~���s��K編 G�����������@�7� :�W��Fǎg	e����=��I��{Rz�eOI��q8�%(� ���u3��z�5{�@jڏ<���{�n*V��Q�F��-~�M�괂���r�Y_E�����;���71Z���X��7ͤ�c�<yVґ{o/,xi�P�`wםKiϮ����V��-�T|�["�.�BTsL��04&��� ��,� Xu���H��Tt�R'U^[�'���ٟq�k��ا �WG���ʱ��\�c`|����s��Z�Z�#(��k��Gi�DyY$ �U34[=�Ϡ�@����ʽ�QﮇC]�eC%�􍢪9@3�2 $�����k���`7�=)��F�8+��-�:D7P6DI���0�w��\^s3�3qٗ�{9}�����9���RI����!=���46SoP�0X�������h�٪m���X����<Y�:U���	��E��J���^w�W���xF7��4�I􈀙�K���.>�.��|��t�m��UG�u��ؗ~x0FB5*�Y�k�=K]Ɩ����+�5	\,,,�	���{f� \FE7����䥩/s#�ݱ��q�����
U�?�������q������ת\x&�	��S]��e�����P�%����iaG��Ёj(� #�� r#]Ԝ���mi����2���ߨO���@�uݬ K%#��|����W\1�ce�@�õ5������_�}���;679U{���k�ԯ3sԞ��J?����P�;�+���l6ͥ��=�Oyj:�����-�O�Ae������Q�3��~��\��8Y�\��hC�<R���g#p>m�9��6��Uҝֺ]*�������؅, ;�X��3Gv��r�{���ߕ��⢴�'k���8�5>n̂U��kTV��+�0W�A+J+*��M[ɱ,,U�|����vk���;�"��C���T�D��!@ �y�� 2T��H�� J�h��J0�����Q�j?*N�o��c`��b� �1�9�}��9@��M��{�e�</��Xm����,un���x��Ϸ�0��o�v�zэ���=R��� ��g>c��yO�rO܃���+����mie�xu3��ՙKwޅ��0�u�iiq%s�,��D��_M_��;���O��*�Oou9u�k�ݴUD����<��u+6IQ}�D�9n�_�P����V�Ś_��q*t�悎�Q[�f��j�	�R�ޏ��Z9���n�ñ��ư��2���x���ΕdR2��;�LD����H���}I��E	u��'lN ���Ɇ]��O5@�0Ѓ{U���q�����p��waEi)�J�� ��|n�7i�.�2{p֪���N���e���Pk �|&+���>��g}J�����oA�<ԧs�z�"�s���_�{g1���G~ �㬑Q��:�is�TZYi�@�k2��H��k�lg>=p�p�x�ymeIs�f����q뭩H�7S�P��dY��{^/�;&1�cں;�6<�>�j���CٱQ�w�����hQt�܈��)z��]���w�?�>��v���ۊM���͋t�'}����ˮT��UڞQ�r��\@,���F��K�]��_�{ݗ�C������{�u��g��M��GР}m#�	���c�e�@�H��]XV� �Ȟ�q�Y�C�X]4��n�V���F���7���]m6*���ٜ 4@��ͣ
�ee��*[�?���+vC�9�q�T��=��<�c�}Y�����97� �q����g��8�\�f��'�u��%B�7���AZ�k璟ɛ,��a�V&��iqeX<%�>;o��"�s
��5Ɖ��/nt�s�"^�}�@=��u����I�N��Vmk�Q�7�r6��Q_Y7Z�p�e�N��q���Rv\�?J�P��ꫯH�w5��0ͤo�ݽ����+--c��)���l1QRe�{���X,�7%I&&��hp�K�j�c�O �jl
?�:���M�P�F+�6Lӭ�H"��d�|�ƌV�D�@8q,L̠��	ȹ��Y�d���� 2���Or��{�J�O�HI��
2Ґ��q�:�ܜCC����;�99��bf�������a����>�zƠ�յN��^.1/�sϡ��q/2f����y��o����d2��F�w͑�}%�⫟�^�����\� ����F8+�uj��ހM4K���q�8#Q�g��W���؅A��&���}��(���	��)u� <�'Yv�F{,���+���޴U֣�L�"���Ț�nRu?��8��1�W]�_WV�r4O�t�y{Sp$�u���{:s�U�fv��"Q����Y�k��i��gq#�i��j
<7� zpO�v}!c�W�u��b�w@s��Ⓟ�j&Q�xt��h����LQ>NJ~g�f܀��70<�w��ƨ�t��i�y(�4�Ѧ��c���{NXolO�1X$����iج�5��|��i�IT�9��3�a�ul�;��^ �^ݸ.���q�D��g��v �����!Qo���XIg�1����J����=���'�o#ϫQZ<�(�`��crS��~�n�]�~oJy��<�u��@c�*?U��,�����.�{��%Ap�E}��w�G3�^�1 �{����w;��0���F���#��ZlG���zb�]`u�v���2>]��M�ڠ����{��(�w�Bz��.K�����Ky?�J�'��+k F���*߽U
Q@@0S��ϲ�Q<e�I-�ɈQ�b�f�p���Km����n@5`�-�u"�J}��o�i�z�&���N�E°�wu�����7cqu2�9N��bۮ�9��4:�ˢ�k}�5��G�l�C�ޓ��M�����Q�yZ��G��j*��T���&��������:P�p�W�e��m�=��m'&x���.^Y��6�����:��e n5�A�hI=�və��	�Չg&"y�v��w�F~;�,��h�(6hx�^W?΍�]Ռ�O�G�VW�Lo��^�~��^��ҽk�;R��0��󰪶<����/���K.�l4�ϚU�{dN���k����0����������2�4���߭�[\ [o���������A���e�ݴ�nv���u�'�L��5�	�H���l��¥�L#��|�ӟO��ޑ��I���/K�?[ x~>��X&@�����	�/�wd���h<��� �$��c����mc�e/��ؤ�9�!"��6a�m�j��G��(�ɮG���&vH��d���F����n����=��\tx2>E�1�ц�H��L��ٕ�{)}�c�~��ǧ'�����xHL���y. b���,�Z*�4����]��x��x�C쿸����"����xYr<W��~Rډ��F`u� 6��nv���Zu�����F`_�~��6z��4��U�l���0?��>����wI��L�=�?;�R�#HPe%]7Қ7Ud���X���J�UPۊFN�EI3�����|����͙m��{)�C;:�̄��l��`[c ��y��C?5�;{�7 �X�aS�?�u�և�
02߭�u=My�0a/�N���O1�x�:`AM��s�Y��W�����7�M�K�4�!�CO?Uي�ͱKZ0Ѝ6WG��U��F�G���
S毕�}���$�ƈ��KM}q���!=���=��6E��g������`i[�ش{8Q�?۩0�킿�4ͮm#��4��ζaq�Dm7$��Q��������3/�n�B'Kγ��[J=Ԙ���iϢ���\�+�*��Y�u�F��f�+mp����_�fTc��*��k�������;�AC�`X�,�kT)�V�Ki�W�^v٣J�E:�/���N�E��� UQ�&G1�.j�26_�-:����Ź0��c��q�������/3%z����G������´ɜ?����Y�ze�h�Imb�
�e�5XV�R��s�S�z��'��rpC�Z����^@W���&�h��3��a\��Qo�O�O�}n����|�����j����`l#��Fg;s�e�o�JDe��(DXE��BԯJ���8�1C�����׾�����>������+��h�ǥi��P�{R�^y啅0�1u�\��� 1 O�KL�Ͷ�)��v�QF�E��2��	a#�ݳ7=�Q�MO�3&��`������N��YB�2�X�Ɇ�\w׏�����p�&U6�bt E�?��?.�jb��Xbm��ĿF�'$�����^���s�={h�~�2̥����ƨh�[�[���L9W���`�L��4�Q|�( ��	}<�~�
���a�s�2���I�Eo�6���7hlv���Է��&��9��t�����O���uY**J2�eN���ۓ^�/H_���gr��slD�Ƽ�g;%0jee)���KC�;���\M!��iQ�F<��,�ɍsL�)��X$h� `�qx�@H��v}qM�#�]?�9�)XCRx�m�JH�`?�ߝa�@�/���xEz�S���@y���9���� X-���z�K^���O�tRa"zV��Dڋ����u�1���Ό���>s��6�K_��t�����yr,��ե�UP�F�P��p\�5�b��DSfu�F����/����
���e�B�-�4�<�����RLS�._�z����'Y'|*m+�jlu={�|#�矦���s3�]7����a�Zy�o�
O)~���	 �ٵ��qՕ�w~���S��t�E�j�H���
��t�+(e�x�i�z^�a��3�� � f�j�pǊ�G`��W_]��
�`m��|J����{)X��1�馛
��}�Cw�v<bn4LFX�O�9�I���?���%q�s#hS`f{� D ��l=���� =P9�ܮ����{�yt ��}(}���ۍ���"U\�z[o�\�B+U���׾"���t����y�V˥�܈���A���H��	Z�6
;��U-T��GU�F#�9$��琨_/�b&�k`�zf8���g|��i-�F��'�m�з���TJh�����ot��x7A�I����rNKKi����[�>��\� �c��ֆ�N&����Go־m�b�#�Sy��J�:�=�;_gO:Vr��t��/J^zA����b�[]=���K3}���� $����Ӌ_��w�[5@H{�;�1I�dȼM&R3�������;L�B���"zd���/6�I����a¨#���w�V������Q��С��y9D=�D���H90����t�;m I����e/+�!₺S���O˥���;jW:���F���oݖ�;wEs9�J��]�����g�9i���q��x��/c��z��������\��j��J`�d�%�ƅVw@����~ְQ��,t��ͲNG;ϣD�{��xZT��bܘ�<Z������77b�"@G�����M����F�q�|��p7������~��<W���=i���]EW<U��� mU������ �?��?+��@L�Ԙ�Ԡ$��T �%8
�dyf ؠ���գ��z��������Q�vm��M��N�Ǔd�ߪr��t����
Ӣ�0�J���������≘��c�w$���~��������=�yew2��:��ӛ�[Â��i3��a7����O~$?ǝ%yLw8 Bno:t7eY�dqk0f�c�`������B/��Xj��b���gdr�䜗�nu�1Z��_f ����l+]������~�3ݝ�h�L��T<�@�b���h���+螥Ǐ�o:��^O�Y�:k�N�
M+�d ޕ�����#�#7|*�������ƹ��O�:�y�i8GC��6�A�^%g�)"�+�>��t�7��X<;����s^I� /�����D�Dc��zt����<��#���O~r���k�{O�O:�7;��Ǐ-�7LG`y��7h�.ߣ��0�$�7�	�����s��a� UX3����ԸP�b��Dy@x�A׻2�=^,��A��[�,�lwW2J�;��z�H}���Dp��P`����cSP����CYYd\����v�m3C�N<{=�JF�/:���M4_O:�]��Cg�9�c��=��!�y����������yMt2���Ez�kϧ#�g"p��^�x����Sk�R����Өt��3aUeJܣ{Я�گ��O�_�ksx󖷼� ����rN}�G�R���g�:��F���H�@`�C�Q�BBQÊ5����L8��Q<�IfЏ8�s���&�Ao�>���6���` ��P(>��3���ท���e��X:�����{�{Kgt�����N���
�u�U&%9�3C�Q�O�!��!ї�ۣ[3�g�|Ƥ=��~q��|�I�j\b����g����1��� ���!?
��V����P��7^s'�7b�H���S������77�9,Xi�;+�u�Y��$N�y]G���:uuDQ���Y:�f�^�ղ4��n����i���k���-@�_���&x�j'�cLpϽ��o,j�c��g?��x~>ӥR�˹�_�
�f�i���4�D۔BL���&�W��6�U`o��`�F�?Z�,�,����������l�UԈ�~3���b����`h��\Oy�Sҫ^��I'�[���N��z���]��a�:"N���]>�Z��,n�K/���ӘOݕ=yw�?�g��#�
�� <J�zz��|��؜@$]��ͤ#�� �A�z�gN����t��$�}:��MR	.����3]'Y3,~2���5ZCD��l�w�D��Ѩ|�����M�fb�����Yo�Uo+uB�Ľu����8s�T��hB��L������g_���\,7�T��1�s� \E��<��5�����t�5�U ����T��?Xm�g׌^��4�=&��:JVR�n|f�cQ\pW��Q�qj	�OHQn�^1�IRv�V��Wr�iD���b�[��s�P�3hQ�Q �'bɯ�ꯦ����(:|����g�z���4�M��bzы�Lg�����-�fs>�����?�'�:��j��W���/� �Q�$�9�>���V#�d'Ϧ��	�,�v\h�?��Û�u�T�
�N��9��֯����1���T�*Rm��Ҁ C�a����H�G������P��������4��/`��be�8���h�jN��ʀ`����tn^Co���^��g��YI�n�v�����l����h��Kq��\�'�nhu�6���/#���3D�����e���7}�zrܢ�>������Q���4�
�muO�7�n�5���kV7�5��wח{l5��x�~Y�zN�ĺsˢ-?��w���\LX6L�-�V��!�b[£R%�9���ܩ��E�Jn�NZZλgcWIFR"{FvY;m���m����lOQQߡ��1�}�p�~����QT���
F�i���ТԶ]��@�o:����o@�o��
�3E�����ck &��1��s��� l�k���y�?�Ò
��ꗴ���R^G)�;�.�i��N^_�y"W�(�����̩0�q�Z��(<Pi�ˢ+�U]1�`8��e�GOu��F�K����@�3:H�� {su��5[�Q���7^̣�I�JG�@FQY@�n$��Id�E�b8���Aa��/�忤�����x���S�{&y�@�p�}?梒�w��]��G�N����R��Z,�s�3%�)Y�ƽQ�xF̬yKl�Ec@l��R��4&N�i��?��(��F ���F��,+&������i�#��?kL[7)�)���[�g�f-���5%	2$��9��"o�����N�� ;�y]3���X�Ъ�Gp�B4�q[��sh��(#&��
 f�*"r�~i43�����8�7�?��R1p3�G�/�/��/n�b���/K�ܝJ5���KH�s���&8a��qݲ����o-�qG�x/j�4��{��__6�?��?�����T��E�UF����Q�i~��I
c����j;�;ɶ�N��7��(�����e��1��y[/*���w��99�w�R6|f�Z	�X�%��������b7gpaLl|S p;_fASE�:f�i��n��_�n�t����%O&&��4d�..h�qhGs��;�����@�Im��;����X0GНi0�`L޽��آH����4 ���z���UND'�[V7o�7~�� s���Q���4bT�_nhQ�S/���@$g=p�qtKs���G�ܕj��J$�)�����.[\<�n��O���7~/����ї]����/���5���R�s��� �e�;�=�)��ozӛ���jbw�"}�Ā4ab*�[G�n-� �Smj$�����)u���	�����/Y�mt����,���=�:���ݭ���CE�a8L���U��������d춵�����L���|�L����7_K��c�׿4�y�A:T�s�@����}I<2S�Χ��f�+Y�e�yY�GЍ%�l���nH��F]�|i,D3ũ��1(�D[�}Ǘ�C_ɜ��1Y
I7Js@ˤ�}�g� ��Cp�XT�1�Y�}1�Y�OՄ*9ƈ�8/�G?�u׵���GԵI�3���CZ�d"���f5}�7�C���y��M�3Ӡ�7�h&1�RH����Z��d������Dʰ"9}������whх�y	Vq<R�D�9+fG��͚��`�5�8�n���΃0MŽ�ą���yl��{�7?H5QxX�G��N.2` �cd,�6>�*���]�c���g��GL$�	��\�>TvI]�bL��ހR~7K���G��_ �LY��~j���=UG�\�1~h�QO�99�������E ��u׶�g����bFOU�=����dT�O�G�����kxV}���KSt�~������y�K�[�$bb�� �R�����ѕ������
*B4���'Ԋg�Lj6f��Z���������轻:�\�2��ۈ����^��i�Ա�y�$ B����}��.}�Z�_�7X1�d�a���9�:s3f���/Y���4c^���q����Ou[;��F�q
���L���z��x�v����M�f��e�WUh�-�����>P���y!�DL�/|�El��8���7��t�'?����L X1zb<30�=:\g��:��,���`�i���iq)�`��=�@z�c&�gH�s�ʢ�f�Ԩ^��S��2���/�7�c
O�l1'(!��[��\� @K�����o3��6ꍚ��µ`�0.�1� �p�_4�>M���`��nP��Ju�lWM�l�����cY�(�l��Ak@��Nj7��L;R��	/��#.97}盇��b8"'L��Ȼ��>�id���ɧ\�Vz��_����� ,� ��9zaT�GT���i�/ǰ�+��`!T��4�G��	hƏ1��p!؅���0��lХ|��0��۱�^�w��~���(a�;��$#�����N!β禠��1�����fq��Pο��o.�9���hX7���-�F�6;�L�\z0��%�N]�_� ��f�z���{q*蘆zrv������C�YZ�1a�VRIo]�L�aEU�V�a"�D}��1M*c���<��s�n����-O��'���p\�HP��{�~ ^��^�xCf`�J��LMu�L�>�m��舭��� ��֔���r"�=��g=�n)Rz��l+�3��O/~�u��dl�I�|�h�
o��TI�k�Kq�:F��G��!�}��^{m��AU�O}j�p]]:}��Ma$�%�C�s^/��'�8@��%�N.���oi��#(�93����ц<��?���{�t�ŗ,�?�V�Šk8q"3	���X;����Iq�1�,nM6��mq�G>�ѓΨ&{�zhL�ed�X�|����W����ͦ��}LZ\>�fڳi�t�T%ܝ<�*#\�3��2�*6�g�[�%��1b�A
&2��&d�ɞNT'�zz<������T"����d��O�C ��������@4VG/S G�!�Vw�aql6�}�dqN��kV��5�� vӆ�T�ek��Z���'y��3�`�V��g\�Ĵ�ey}��3�<���#ŧ�����������I}���-0��V�@y���EE2��&�s���֞����#5���������;�#�ӯ~�u�6�p�����Ύ��^&�jeG����z��/|I�ǗIȎc�"��.8DU����ތ���G>RحF#�TY���/:����4YX��D���v�)-�.����%鬳�(�t[���N+˽<A��Օ�0����үQ��l?���80F2��W�i��f-�" �;��/-���)���ۉ�~�w ��5�(��<�����/��,Y/�!kG]vd�����l ��p�
�	�d�l��j<g-r �=�����:hʹR�C����l/��XI{����v��鑏if�r55;Y:Y��n���k��j��ꪸi�o#j�L����!pT��y��5���y�hxv�XHϸ�2.�	}��a�V�Q�~F�ÆŹq��5�Z�C#�X=��L�֘DUU~�3c�gb�`w�ywȆ���*�� �b#���_�bQn�� ���7t3�~���L8���Q�Ϣ6魎E�n-�����ay.e��a��׿����oڃ<1��مt��y@gw�!���n���+nzD�u�U���PoV���{��aA0A�ie�Q|*�������7��9�\�C"�N7�	�>��O;���w��2F���	b/�k�˭���K��3�p`�Jr���Ƴ���1�[/^f��.9�˔�fb��X��E������' X&AA�eʅ�f�`6[���0K����3�%U�#�����|��Ԟٗ��=P�� -�ߝV{˕zb�Ve<��^!46|�� I�6!0�������4�K�����
!Τ�%�i)CCntd\�_^0p���w�l�������k���qI�CU��7*��X����0꾜:��a�kW�zе���"��q����%ȸ���E����X7���a$ ��濺1���Ci~���*��O���Jlj�˱�i��Rߣ�����Eo@Ft=�FٝhηXbD㿑��N]�y"��^Ի�7���=�O�`gp���@���FBc-���%`	%����u��ArU�l�w�u�T��F:�z;�t�x���D��{����Ꙇ�� �p0�ڙ�\���ff| ��MeW� �������6`�N��7���FĜ���&��aM:��T�5�$�[p ��CUi��O��ԙ��E��������9O8d�\�v!>�3���[&��&�| Ev�<t��%�D��u���ۛ�PT�3 �;��z��q��p4�}�����O��9��Q��=�A9��ü�������
�x�\ԑ]2	g���Dܮ��j$���cܙsQ�|:Z]']7ј�z�0�!"V��l��74�&4#�8�u�� ����%��M窚EI����>��-�G�>��^cl:Yg��]ψ��TUmW{���3��Ŵrt��9X���_��-��/s�V�L$'$���� ����-�;�o6s@���(�<1(E�� �IA)Ƅ<��qyŠ��n�Q�9��G'L�j⍳菂�����swpM�nn��6�T����h�h�����u:��	�P��j\D��������i%���l��#�9��V�$q�lU��A�\1�������4`����i1
�D|��jaEN�4�o4���K��<�Ws1_�����orQ}�C�S�+�3ݫT���<��=�C��=!y��6##�p5�O����I&4�yu���J��ʌuZy]f������R�]��vJ�!g����J#��-���'�U��>T�#TI��FP�n�5͋F_�hߊs=[O�m�;���h��n��\��ϢU���-.$���4�n�.78�fLL;�D��5T�pK�/��u��,B��H���^�5O�cu�-�5n���n�R�c)���?=�nէ���P���;�
�űӛ�;�ft���m��H4�,Vw2��vԅ��Z�Z���)��1��(�,��*{N^��#���6d���F��:��sˈ���gh�����k�K�]rNڳ{��Cbڝ=xg�Ӯ�*�{�y�T�k��g.�������ّ��b���t;�y%�?ٱ��J�FqN���ʃ��{�T6���|�M1MuSh��	��`T�6֘Ҵ���\����J,�W�u}�h��u���&������G���E=\��h)=��'��g��r�;��sF��H���?�n�-R@��xs��19�9#d�Nds}hMvb���vYpl^C� ��wJ�q"��!���4ؔ4~q_|f�\��F�ׄ��t�ENc� . -���2Gn[ �ngQ]ǵP��ր	��@aY�(��&6��uy%��e���=���k�s�{u�(ޞٓV��t<3�]{2;���\���SXtņGE_K~�z0�FW�W��r�(J]p���TM���)��,�.�Ӣ�'��t�@����Iw�N�G}��wu�R���Y@]����ˤ�R���kO���0H� &���Iˋ���=,�<)�ͦ��F:|��#��w��f���VTaT��R�A���ޢ+�(7MdU��i��3T4�L;��]���玢*M 0o�^9,t�$��F��u�ܵx'`��ݤ?S�ZA�y��#�ٺ!a��/�fߨ������G�5�]��/�^�)kp�Vj��_����)�0����J:��FqUC3�j�O�+�t������L�=���cX���5�)��Q�ZR�8���������M�c��c%xu�1�6�Y���{-7��MAx��M��z�3�)n_щ^qJ�(]�Q�'{|/��3���Ȥ�P;�	��J�k�K��>��򦏦K/۟���G���۝Ť����®�<��lK������i�I�PWO�uc���i��Ӫ	�Of(�>O�q�~u���z2p|�ȯޅp����`�F��o����� �!�%�3_>l�	U!���u��X�����6"�h��k����:Y*kfiq)}��_I����ӓ���t��Jǎf��ٕ�-��(����-^��Z}�~ҝ/�O�F�C�_�?�Ҳ�$V�u7ʺ5F;�T����n�:����RS��-��Y�hQ�R���5�s�~~~�e�^;2��ǧ���Z�TϏ�i������t���7қ���~�.�g�yR�������Faヰ	�~$���|V7C�� ��d4ҝ����`@k��D���TtC�'{O�5"��m�2��$ǉ���A��n"��`%�B\;4Y6�|��*�~�<�$̣!��;TlH0������'kl2y�`�:��bجW���g��+�7������}��ON睷7u��|;����'�Z�*׮䫞s$�����9�;��ű��N�w���:j�5rwJ�~S���(ߘ\b|�k�_q�h���q�(Fx�'��,������_��1�zu�s)�=�O�<I�����&=�W��>��%���2�Gg|���Q��x4���N8Z��i��t�<W��  f���������<��w���Qw͹�zy-�g�C��Z�ܒD���Moð���)F� �sN��P�{�X�ي��:eذ�]"Q����Xj�Y9���Ψ$jG�<r�h���8�Z��v/��V�3ж��LN�G��z)j'��>C�=U<��umu�`���D����'8�q<tџ4�Tf|0;!VM��1�Zd�3{��^p��:u��|b�M�RUy��,�u[閿�3-/Qv&�R�S�=Wr#�$��I��Q��Pn����H����.q'T�m;�[�,شE��N�s�r�df7u��j9ݩ`�օ�� f���� ��c����9A��djzr�⼀7��]Y-/Z]=8MT��o�RN=zdt2;˼��b��Iw�u_&7�t�E�|+�ػoWQS�
��-k��N�7Zw�mbE�k�q�k�uf<V7��)��MA��sv�dQ�ڼM��`"�	±	�u����ؚ�q�E����w�-�r����R��f暙)�"��ԙ���"���3,Lx<l�ᜰ��u?tq4�E��rӌ��p;-2���9��4�Lk�C-�պ�wBg��׼�ll]r�����a���	C����bXSg�a�k�� �a�a�oX��Du��wDɡ�`�@%�kZ�����Un�Ʒ�$ٮ�g��m G@���5O��y-�:?(�H�Cz�fk��+�̠1>�f4u��ApZ��>#�����ql$�Q]�mLQ��e4K���l�gQ��-�.*�xg����c���n}���3�����T�k��,#���3��52��}/�ڛ!x���K�����t���ґ��y�P�1�q�[o���w{�b��v� W�nd�Vգ�h\U]��X�!l�EU�j2ϭ�D\n(�\#�ȑ`a[+`����9 W�lh.�h����P{L�8+��p�>�&��I�F?�Ra�|+��g�s�>�wϥ�_��t�p73�R�����JZ��`<[�ёw�0��cp��r3 ���g7��X#1���љQ��wx*lxsn������	�t�2Y�����|ŉT_Q\����Z�U�#G����]�RG��ܮaz�k_�.�p&]��+������r�s#ZM�/�r�4O�S,)��������� �e�i5Ĵ{��	6�	ڨqO���QԮ���4���zO�> K�Q}Q�����OY����wo�(Po�$K�?�b �k�G���f���Ͽ�{_I�����������lvP���ٚ�l�\��4���>����>'}�w����URY���-��J.��z����]�˳ҷ�	�9��a�
�p=.^�q���MAx8h�0��0�:�x1)�Ư��x���6M�+�C�k���D.ӌtu ���E�;�^��̦��ܚ�7�^8�Ծ�$*q2ڗ�7TK�>��|�l������C��h]7L�	]d�&Y����4釶���ʄy�f���}�<��l�uт.�#ޏs��PQIX)C�<���Vu�=�#�9�I/%}���h�,}1�2&6[5���n����O��s��tB>_|zgJƲ�\�����ݕ����Һ���:�J��]y�<��oN���E���$��.}�O2��\�`x�x��޴K�an&�(�`7�N��5"EG��O���/�[��t�f�0���AT"��٠l����h^O|��5�\S�g�'�(͝�&��*<͐T����~�+_O���L�+���);�K�~����6*�\)�R�yTÛ�M&,�g��o������IFK���͌s�xND�y"M/1�Ĭ��ɫb"��PĔ�Y������`�(���d7&׻�K�{%F��K�ϴ�i3���6�^&+�O��̂WZyø'}�K�ʠ|����p.�ʹ�{��t��invO��-���8^��h;����������I�Y���s2���<�a�)�S��-t�Pr�.+!���j�<��^z��W��{Τ�9�2LE+�3������:M7�tS9>:��>c�����/y�����t�UW����-��9d����o/;M�B��}|�����A���[I����Z��Z,9���y"��Nǎ؄��@�DZ�Vs.�0e��P���x�p�er4� A��^�<�����9����Lr��i3�>��O;6��Ģ�3�+ L_@4��i�\� g�,��E�K��G03�}��v��Jȵ�t����B��R�'
Õ��c�(j�Z	�ڿ!`��"ޗ�8�_��{���tÇ>��A��I�wq��OJ��|)������)��:I�d���70���^���� %%�ԛ;M�M	��4�~��+��#8w�7g k0��G�Z�CI$��<-�Q{�h5[�����)�1��,�'�ܓӳ�y]ڳg_��ٱa�N&��x �EN:�T��V�K��V]�j��ԔBd�?���.ߛX<V��X�1od���|�]��d�{h�Ҿ����f�f`����nx46$4�9XmuD�iup3�D�&��n'\��O�\UCXN����t�M�T�V@��  ,N6ve��*ki{uۀ  ���+nz�����Zt�����PE=�6K�����Ozz0��O�ռn��u�Z�MGC��s��u[fó��S�Y�UW�K�Kl-�{�/fD�oc�SQ9V��&�8S\�����7JV�x�3������k�9&����=8l�l����+�O5 ƚ��5��d�A�6>���yIf�ץ����j�h;1L@����`�щTL%3�ᛑ-��#�9���`>N\��h� �3�peۃt�H��bR^L��2��8��9�x$�#L�1�-7�J�<`�n����n�r�	
�7bB%��E)�%�j�ZQL��+{�0����^��Έ�6a���(�\�����8ǔ���0������?��-",�Ρ8m��lR�W=��'���[�HEs��H�����3N��B'��%��WRZ.��о�v�=#8X�a/-����[�y���+éj'��-�K���������x�;J?�[���CC�M�o�q�4jL@L"�9�U�P�tp~3F`�VQ8�͕�v��d���i �����~#?��t�W���~=���3�;Zyo��I�P��s��-�Z!��>�/y�K�w��Ǽ�u�+���b'�X��0�z�	�$�LN�����GfJ�~��-<����S+l���TJ�4LH
>�A8�t���I�	u�y�K�9D{栬PF㦿�0M�\��y^�E����cX��0�EC4��ҏ��wu�y�GI��晽v�H�k�Ɏ$��௚�r_���V�r$]x����F�T����.ܥ��<&u����/�{������ )�fc�!K;}�ӟ.����P3��1�>�&��� 5�;*��1:ڊ"��g�������1c���}n2��N���h0��/�,t�W����)`�t*`�e��{'+��Э��2QM�����:)asF�=�O}�:Jv�v�Xz��H���I���4�����ݝ���/�Gjj�	��!J�V���|����{؉T3>��殺���et��Ǩ�nX�fF���h�Z 0aĬ�]�ۚW���7K�RSVE7W��Ut�C��)1'�a��sG76��Dl��Z	�5�܉��s��RF�f�iv�\z�/�<����N��^1|�;s��qX�\j7����uG+�_���n�ES�B5�A�1}�я~��R� ��RmK�q��� ��
��>�s�^�(fx���3
 �G�h���X%qzK����R��L������!|��a1 vI� 8�BG;���� ��yk��s�k�oD������_ˠ����[�^L�������<@�i+���{�&��K���RvTJ��Gm ����H �0�y� �9����3�h,66]Æc����s�噙��!��t�YG�M��:\�M~���]�Q"�𞱁]z,��F!H�w��r�2��N����]��^<v��/9��~B�������L:v,K2�nI�ngf��R��y��ݔ&�rm��7 Q�#ρ�FX�)��4�0�h3�����
=�/��➼4�2���ê�X��;τ�VAv��^p�y�#��~XtK�nR<�)�5�#D�B=1��,s>����ꜛE�e���zX)_��W���J�]�1@#����X1��=������\zFz�k^�f��<p�8_��I�L�s��@nϰ���EO��&[cc>���U%�x3���0K�u?�m���h�tB�l��>�����@+; s�z��u#d�3���"F®)��ҪM�T��y�7��Bj5��K��0�/9��I��,5馛>�>�gQ��ЏN�3����?���l�uE!b��}G��׿��E%A?��.�U</�y�w��]�>%%<�x�3 �/�P�Mi���Ҷ��8��q�]C(��
Z��q�y�s�����bqgh��}��W�� ��Ibuc��T��xH�-����B���qC{�k_[vA���t��t�;���"��qq���2�.��#�/��>������;����oo-�r���L�1�e���"��DܿO��Qׇ���ԍ�X��X����I�J�,�t=&;�`�Sl�ޢ��{B�C2�'��em1��x����~�1�&M���;�K�X�a��fܞ��z��L��+����=���_~�3����ҡ�{�7��t��{K��fs6���R�3>-����y0ȿ�e/+��.��oxCynt�|nE��!�XHb�b1(��(�sn�EyN�Gm�=�G������ڈ���UG4Z�ҵ�[%x����$���ۀ�$oc-��;��+�1������"�y�~����������芟��g��e�q������¤�sh����ӝ?�7}�O�:��U�K�>��H�b�+j�F����Uʲ�Fy�7i�Ֆ�"��XMs�[��m*)���&���b�N���&�Ci�~ΓY�^G�k�s�qm� '�I£
�{9���K��;2��
�3�%�Xa���`�,q}��XŢ=Eo	����õ$@T�"�a�;��owf�sdm��U�������t�������aw�u�T�f��3c�W�,�	(�̪��G�e��������˛���"��;�,+��������x	YS��O�~�����S��k�2H4�L���8����'=��PG�G�V���ʺ]6]���k�ݍ��S��dwٲ�_d
ՀV:a:#�C��ab���\^ӿ�ɕ돆ie9�C?�/��<IF��[�H�_p^>���� =��\�u�-���+�? � �Rg�?���.̦?�fA�U��L��۽׺��k1_�/�L#�� ���h��4�kØ�7���r�fk~Ƞ�E�,��^�}��Q�,[Vա�� A��D�M�!l��WW��J�b���]E���݇Ұ?���ޔe�|��������\e������7� �w�H�آ�J@����'��5�)nk "�D��^�)�|3zOhP��^��	)1���UQJ�4Wv���R�hT��/4\cavRw�f-��."ѰJv삈I5h�υb�c_�җ�����I7�pC�\X0j
\G���?���"]�y�oa~&���H�>��tɥ���fz��}�J���+m�����yo�F�>�g�����:ӭn� .8�n@�ewd0��E&b��9�ew;´�[��
���Pώ�z�-��c�y�v�q|�<,�A��xǄT�SC��W~�p���O�_r@iD_�6Qݻ�s��\u��<R�k�Է'23l�Rg��.zę閯ݟ�C��WJD*�#7e�Z�̂���~��9�x�$���7��<�9�?���T�A�~���wxWi�:q7>]cـb��8~q����X�X���W̭���l�s;��h��y��r*f�|��z����;o�ܰ��sx�)ylԁY"����������$5y5l�I��|�3�)��23Fm	LS��ưL�QZI������_|Af�g�W�+CIU�QXq����vU�S@$~�ӞA&<���T��fM���YwK�Qb�m̱���T�a���*�#�ى��F�I ]�̀  �� @��)1���[�.�c��!��ڊ��kK�aT�`��QEp?H�lJ��j����!�W���if���ϥW����;ߺ?9�/u纽ci�ފU.-/�
+V9\��+V;���'�X՗����o�v�P�oHƀ��싸�}x=n4���x*�4�����}�mu�E�b�*�&/v��@͙�+
Ɇe���Z����g1�E�gXA�F��D�<�'�����u�G}w���)�Y<������t�#���_qQ&�t�b�U���**��J/�~�f��6��D�u�0�L�M�)����n\��N�im��4����U�O��{���(��J��!q|��z�H}.�D�DI�s�o�g���Q��X-id��2�<n�[��/�a�f�XmF�6F���C� ) 0��	k*��}�������e�|.�������͡�OOzʣҿ������Ng�ufa�Ԥ�u�a�_ȼ��p�IG�z^?~�����/�R�PF5>plԑ��Dn��TS���Iċ��Qu�����d�����}#3��p0� ��A����shb�b�1�4�ޱS�!�L�Cǘ�'2X�75�:6un����uT�E��;*�|~�0]}���}�.���X��Υ���i��?-�3#u����q���6N�=c��:˵�.�N����f�Fu��'{�h�ޮ:��D�`��+�v����國sW�<@�8�0b�)`k�M��vp���ͺ@#ܭ`aVW�	���_e���fL�!�s��@o[�_T����iFs��������˳s�t�Ż�Y�^�n���L�qSg&ϙ6*�n��y-���R��0�=��O��C�����Pb��sLc���8�Ք�ԙ�;��6��&��W���y�Z��E�q@����m���F�v���0��i/z����+�t���ID7�>Fk����/f�ѱ��7����Y��q7�9\��E� ��� δ���}���T�$:gG�����A������-}�;�����M3s��޻���eί���/����ԊZ��@�iQ���+����K{�n4.x\`������������4p����:�Ό��.m���ν�U_��A2�Q��	��L�f#�dmH� ����Ju����m.c��8,�kFC]TM߀6b���y��3��D��k^߼��t�_|=�gKY�Ngwcj8��Rf/--Ri��:YR����fSM�S�+=����ځ8��~d�yғ�Tp�M�d`�Ȍ���Ȳ������r�ʪR��$��Ҋ�B 	#$�	!�1k;lf�D���3቙��n�{"�1�&�=xŋڣ��2b�X�&�RH�U�de���߹����n��r�L$���Ro��9��?��1�DԲ�1A��zL��Jrw-�asc��T��v4�[et��)1,�D`�+�ޢ�۽`�{��Ŏ�������Wy����L@���F�dI(�tg��}��Q�#����
�ӟ�L{��L��¿�@�8��}���h����/3w�Y;rx�*���E�;��7��Zb�]���s��(5����yc�6!��� ��Vmh���ă�V�B�K o.���}��7v]S�y,iF��3G�$(.��LR��浤DU�`�(E*�6��������w��W���wJ����pkAj\�}���K����LP���-��_ ����	ϡ���ȋI��趕3Yx@pUL�����?�~#��/�R��ؐ��y�5�p#E���g�
0��_G�)���ø"���F�cUdֻ&�u�N��N�2<�Z��؅0������;Pc��i�3qxϮ)[�De�(�D&U��N�k!�q=�0�J��@�
��#��2����[>��:'¦�C�?��V �r��ӧ���O�f�`�Y�\	s\����K��f�5�d�^?�@=HϹ�+��_�^��u�RE��T��4��ȧ�	ӭy�C��km(\
D=��m��@�����,��Ԥ����"� #n?��|�"���"�6�÷��.���3sԢ�N;�jVo��|���frpWm���|�*�}aN�D{K7���+�^��\W�\��j#a�������g��0b66��J��ؾ�D<�P������g��+:��W�͠7���8���ګ#"��$fg���ِ�'�z)B��'í�!�K���L�Ag��@���X�M^I/X��r7RzLO���&� �$@��85�OڲU�jV_���#ǭ:1c�V�z��v��@�2�IA��D��p�C�\�QQ���8J<��_K��:��ꈥ����leD�����d�S��S��B��Q�{��ET/���6�ݻ0-#� ��}bڎ?a����rXS��%o�	��'S(�j��i�c���*:��a�b~��T?ZK��BlvHҤ��qc�C��y\�{�H��s �T���O�6�|<W=��
�ЩY60�sQ��N��k,��(ّ�XE~u�
t�F3�`���X�Y]�^�Ʌ���|gO�-'v"j���:�!��e/pK�u�7K�L��'���UJa'���!ڝ��}�f6��Õ�9;���?��#�:\m>E �6��>J_��+�����J��L�Z3^�/0՟���|//-��x� ��Bja�.�>�l�Y8%��|���eo?�n��%v���5�#z� �Y�I�)
@'P� v#��<Y�|`�����/��{�Tr�
9 U(2�-!0|�Y
���RܗvQU��<P�XC����W֨v�$�^���I{:�r���ZqY1B"Z��>�������_�'q��\�zΐ��@�K���޲\B޻ m��@����]��a�hu欓�;x�����_{o��ɤƦ0�[Mc}�,:h5$jM$����������a����К�R	m ���rΫ�._�����z��h��>�e܉�O[��`�j�6o�loy�+�U��>��k3��T�@��Y��rS~r�z+%�2f��e��sA���u��l��7�
����=@����x�8"��:Nc��2/D�����*�ʟ�&F(��,�m�\o�s�O �Nf��Z�bZN�t�dgR�W����A��%��x�(�׏ϸ��`�Y����Oy�=�'Æ7|��1	b�FY�];��J�c�d�S[�f3�n���[��軒Յ.{#�!Gq1�!|���a!?^�"����(�96h<�~	x�3�j5��rA���m�<k5�X�����42����~K�[l߾zn �t��@_c�&�����20{젚��^T��� �0	���SQ	�U=t�✹&@�Ď�^AJ�i]�������~
�N'�\��70�-��kWzX�ۄd`P#�������yp�� RM����T%x���lI�A��B�n������l�[n�:습���v���WZ��l�&vx5���݇��Q�<?��w��Q4�h��9y��=s�{�]��=AF%��ǺQJ��0�[aݶ�6Q��q�ngE�x����W��]q�Kl�maΕ�L� uv[�Z.j>�G��(�P̛����9W�DEo�(F[ ���q�W�e,S�>����6Y�`/�&]7l���p����jt����A��~/ZD�����-��	<|��>�Ĉa�P�E�����}Z���[��'�x���w�զ'7[�r4�6�<l9��WJE� M4���\�0���?�/��V<�sL�gi�Ӧx*�ޜ�?�Mb9 X��d{3"�z��A��Bs{�d�)��v5��i�����J��r����ޯ��/�gs���_�2H��1�p30s��Mo��n����&)�3!^U�DEb"���H/=��5ߕU���1�:����=��/�^�#!�ƒ�-2�Ҟx���GK��r>�8A�*�����Jr����b`� �{
�}���&s<�[�m[w�S=i��������ο��p�J�̇�N���CE.�G�y#���'�7��P1<�/B����s��h��o�ɴ�EYW�zf�(�X ���"������e2es-�]T��̘� `��>��v`���n='���/b��S]R6�����^۽߭�Z�&5�"D闯�&WL�_ᑷ5q�2���^Hܸ���=�y�s7�k�.U�>މ7��jJ$�7�sG~��8�;�{=�����Hw�c*��E]�o�~ǿ�ı�yX2e�����_&I5`������ӵ~ވ�j��J���@9��I��z�i�������$�C1��O�q��j�<W/	�or�7�&��U��B/���@�Y�7h�o��"�� .h�X�_t_������'҂�����W�)�iX��\fv�ZSv]�*Q�011�3X��^hԛ��Oe* �YX��ʞ�d��_�
@��4wG1"а�?����������=��Q9Y�U1��I~2�z�Bq-���������/��}8퉙8�ʕ�.��۹k{xo��t��V�~}9��"�<�]�[�=��O~qkg����{ ��{Bxg-t/�d��-N�a�i?a�!Ë�:��j)��_ۻ�s�ħ�/�G?���`T�t���W1^��g染�,λ#zfE��v����E���Q7�'a��}�;��Fy��/8���^��:1��j�
�����[�;�EXj�+���Qs�8��ڄ<���or�I����,pdE.�����Z�IEU������{&�ũ=}�i;}�6{�O���\p���(���u%�ig�o���2�[��" V[��P��s�꓀ƃ��"�i<}ٖa��Un�=��Kaq��f��C�ߨ��B��p����"��9�9�^>�gy��1}���W�U{�$��o vo��QHs�?{?��}nkKX�[1,���6��6��j?��[��~hG�խ�:fI�a�f%��$�eU����W��=ޟ7L�YOZ�\�߰�S��r�=jw�R�k��5�c�up�����;��sv�%[�y/8;L��(&MLe��-���p�J��(2���U\�9��yqT���X/���_��׵�3�F3��},r��V5>BI�F��g
�;/m	��o��R'���6z�H/�K��P ��`��I��W�����"�΢$�LR��jiZ�� '� 5�L���y��߿~������y{Ίf�y�! �i� ���)�Zq�x�f�r�.5Ǉm��1�QHcA��rF2��-�P�IQ��5���S�m�z?Q�����v�i��~��sΌ9�X�[���U�����Y;v4tvi,	�X����٢�������@�"Ǩ1й�ĮS�D�g���^>ۛ^���{q3� z^-N�Q.I�|tm���;���{�aݛ�DG������˟�!xc�f��]	g��� u�R�)SB��n\/�2��Пٖ ƍ�V�{ٕvڶ���ө9J�g#�q�,J��d�5���Z\�K6���AK�?�v���%#�hʸc��R��*Z�}���P���z}�?����そ-�,J��a�}�DԋA�*ۉO�7��7�f�UȎ��r|M��e'�fƾ=ŅU����1g4+��8*n
zv��w��O��^* q��+��7ho����?k]S����(��{5Ű>�;Iҵ�;IR#�;^}��QR��&�$!���VQa~�VL_����[�,��=��>�����֌I�[��"�N��ju�QNia!l�]���������_��r�Z���.ُt0��r�=��T<]!��NfolO$~�{����b'�J��|������|��B\U�J$C9f��sv`5��Rn�"�S���}<�P�,+��Pa��E����K_����}���A��V䊼�<g\��.W�T_4��,j�{�N.WV*ZI�>
|�a�f�5���>A")r�(ɍ�L�GD��z8��TT�����&�K��J���I4(�����s?r��ү� Ҫ���)t�k���A��aR]�y?Ӫ�����X���i�gp��⮏؇>�ak��Z�bڦ�7�UW���\p�5[��)�5�>�w�D�a�����U��8�Y1LE��4�+�%G +�b�_2y��{Y��QT}�W/����@�pjo���!����ჶ0Oٓ�0qjv����z��l��C��o^I �e�n��D��$�E}��d���s���< �L��b�J�_��m����< �"� P ��r����W���=�^ �$D� ��|~��⺤?����??r�@�������ƈ���8s�~ ��e�+�\� K}�Ky����RO �ܟc g�!<�M�~��D���򒍣����D���&lQ�09U�Ns��	\/Z̪5IY�mZ����=}��0U*fn<ƭ�s�Ԧ�S3n�8R���o� �MP�N��J(]%j��	N8)����pd]O��"�V%d/�	KnT��0�8e���l� Z�<���x�x p#*�B�#�|)}�>H�H�I�3�Q(Iw�1 �<����v�B�bY� �!���$} �'�61�C�u�^K� �~��u���.5цqEu�(Ւ6C�K^���o�̓��92'8_9 ������w�7%�`���"�2/�@"���k"��]f��}+�������L0�h#��h#���+���6����?ǒ��{r,� �	k�{2wi3k��Tƞ́$2 k�q�����_�r{
������w|j4~����uJ��a�F7ϰ�5լ�ZxtSd��j��kA
	��MQ�#KE���'�c"��j�y5�E����E~���}}���>� �+U$�}�+l���)V��><#ի��t��X�u;��p,;==K�3Q�<I�(&��_n�^zi��|k��`�3AI/�����n׿�;"xS��s�+��"r=>�`�Dz@��E/z�IA�J�mǎ�0��m��CN�(�M�O����7��3�ѵ~*˥��W��O�FLyOx=����|_�qC�TE@/�CWCE���g
�3��c����U�u�ߜ�Q�X�w1��1?�r`�q?�x����[����7P����CF=y+(_,m%/�R�z��P�[ 5�q]@S��5�Us���b� �!�2����e�P��,�	��)R�E����l�36���X�h"�&lێ-��+/����\km�=�0��Jo̕��3	��gI��T�����͑�����G�#�LT���K6=*� }�I{���:TL��Vj3~�G��E��讽N�RIڝ�M���'����n��^xQ �kbZ80�k�d�<&���&zB�DDB&c��B�g�g#�������}Q�p�7F �a ��\�EḰ�� <Q��^����D%�Ī��Q%��������3����
���Im��~�?���N�YXԅ�[�i�86J�Q<�$=x��]!�S�aj&�=�L���	�c�Ј�,0/��V��H t�|f����8�9(�8�y�F�25�#��1��X��E*#�a��\-t����VF/Iq�Q���y�C<�r�;�t��}���Q��aé�r���2��܉#�%aOڵ];�����F��/��Z���0��Mx�V�Z�6=#�2�[����I��V�4&��+^�
���ۣ�8�ӗ���1/0e��z��C������|��:,���4���x���Y�<�����v��),a��M�,�Ns�n>�l^t��t��ag:�W�
΀�!�p`�Ʌ�]���j�}�����ʎ��"c����Q��w�i?��?o�''+��u��H�-��h�����ݴ�w�<,���/>m�f��E�jŹ�>�F=p�)���֫5�u�^U�d4!5h����NznΨ�5�����,nE���s�3��� ̢�w�ׇ"�|q&޸��<wDI�f��X�,�é>`�����.d^�^|Fg�x����u��F_�I��SqJ�bh �J��A�h?��E����0�6m� �\�)��?sԵٙ �NV���F�c�[&�3�Zu"H*iۦj����M+U��Z��e`�ݾ;$�P�UkC���������+_���9�o|�#C���I�>��&ȳG�T��넥�{�,��!�0�G ��Z)�px�k�	��(6��M�͛���l�� ؝��yf���	�>ɧ�I�?X{:���.�"���R u�kq>0"����ܱv1_tO�$��7t9G�Өpן��sׄ���l��M��Hy�p�q�y�r"�[=��N��0#����H-�QRzMMl�V�<�Oj�0���a@�O�(�PŰk��7@���b��es�).�k�P9��ec���9ǵ8���5�
��\����yϢ��zp���,\��p�p�������%��}�o='����0�5N~��S�	j4�1Z7m���
���4�ԷT����߶˞s��>繡�%�Q�+�$�����_�U�!�C����s�p�s��%%�o��Jq<c+@FR�馛�3a��5�^�%FI�<�c޾�/������/�g(}�����%��������&���9�X�ͯ?d���ý^�`Lnu��G�k��6.�,nC��{<�������|�#��?��?�7����Ap�StA�`�]����:e��_~�����oٿ��_�߷r���|4ט(���4L� @�B,�|�m�5�G��a<�4P7�:r	[�3�rh�J��\@J�x� ��yϕ�����g�J���E`�$��F��@��a� �Ap�0��o�}��ĸs���}U�$�F	�̱0J 8�7��b��pq\��dh�I�+ΐ�2��8�L*>֟�����$L"�N�n�#�Gn�F����������{���j�˿��&'�m���"��������$�Vyn��u��W��mx����'���}�8Tm�b�Ĥ��c�d^������u��'H�K�bs��{����VXop�k�����Q��������"b�1�i�2�h��XJ�"]��3vFO��f��Q���ɋ�C�̄G��7��w<����"��t�ϖ��M�y�t���#v�'ﵟ|�+���P9n*����fä�M�Vޏ뽎S�n-4�>7,���=�z�azY��E ^Kf8ԟ$�le�l�SD<t��@%zz�"�1�Ƙ,��A�����\��z衞�!b��ay!��l	�7��g�T 9��& * G���Gnm*���K��fA������c��J�����s���稛�Ƶ��n+z�;ٸ;ڱO}�s�������4+'�Y���l�1�5b����?��`l��/��^��WG	��t�a�P�s�=��s57 l �b~@|���֐rxh��yހ�7�7U��P����a�	H�ؑy2LT'�.�{�!��3���#��YF&;��/t�I̎�N�D�a` �{����4zd:����_��x.��E��̊�;>�x�ĂQ(v�DÞzr�]tɥF��VNx2���Rf�[f�r��񐨥�#ø�a���)�P�/��$2�3�@~���R�9 ��� Wɜ�h"j	���3��׼xj�h5�2h�!	�4�>_5s�{���7�q�=��I�r���K�"-|��w|���*�#��!{�|���q��~��:>P�$�>E2�J�)1?6����$fJK����
���u�)�I�կ��??/�O�������8Ό��-�_lzR�ȷXz[ ��Fg�f���o0~y5�X�3|V�E�2w��
a�k�	'�r�M��	�X�t+t�"�GG�k�B)�(�Cް^'H(����u������-�qD8�l�z
0���s�uH���=�)����6�NY)�����n{.:7�T��V�\�ʢ��tn.�D=��* ����`H��wYS;�G��-F���������~�^�Q�;�"�2X�T= �`?�R%� MZ�s�������@T�u����	�5�l�"����B  u��@�W��j-x ѫ���ŤDޯU�О��5�s뙣0��N��ȅ0|[� �i&�����OX'��|c. ��L[XC�6y��ܐ��m���*�:yI<I�P�T$�1��JqTr��v#y��j����ل����J���	C�i���k��хl��YR��N�T4��Kc�2h�J8!������G���:�� j�c��B k�ypF�R+�F��sv؏���p�r����=�U�������D7j{1�b�������yė@g�ܚ���3+�L�mY)yN��?f��kMî9N
�������N�F�v�bëE`�����^y�=���F�4;|�`�/��.���S���0��,��#�/���XI8Tc�(�$oFa��d�+[æ�C}�6�  ��IDAT�{�jS�����ݼ_N8 �8t9���[e�G2����h�XVj-h݂�ᢆn��[o��	_��1�NZ�F,�.�M�Atmj�do����=n�+_p�M̴�Qϸ�Nhnti�p�#R��'��9*m�E�ٝ%���!�sJ�@U . �$V���=j\�3��Î�z����\�z�0�|Q
7�0����n�C"��+i�!\J�����_�cs�;v��^h_r�=��&gg�n"��U��\�U?��i���} �ԋ0(��N~�#�$8�G��! �^]���$n��:FҔ�^��Ͷ·N��ˣ%�m�5�Һ��G�����@ ��7s����� P@����G��N�k�1�<<)=4�HK��\���E�{l.j��]��l�.6�#v����n��a�L����yu��&�KDU�5�"?Y�ּ�B",˫d��s5 ���Z�"�֥���~����b؞
��u�Q��b��:ܵ%|�����a=LN����a������mێ�;�[ϳ�~�` ް��Sf�w�.y��֩�\�ۆХÄ��o��0���>�v�0e��B>�M82�z�(5�����z�a����n�[.-.�xB��&β�A]�:#�_�ThpQ����������K��p��{�[�b����i��{���g��6�t;�|?���|�R;�[��������a��)|��N�D��FgI#l�$@+���Pz?/�+��(�k\��B���*ǩ��Ѩ�4��1~W���{H��c~��+w��p���@�dڴ90@Uk.�b����}���Y����?�J�6���ێ�B��wZRg���|��	k��s< X��{���{��8E4�ە@@�A.i�� o�	�e��Ƒ��K�Nw��5J�v*=G\i���v��¾3ޥH@Z�pQ��nG�uL�k����aN�~Ǻ�կ~5�������Q�|�3���ǃpֿn����_�;v䐕*d|j9|�m9�:s����Ls�\��H(��,�Ч��n\㢉(5�al���Y>�D���E��ն� <
�W�E�jQ�����b.~�/�� U��%e[�_�|�c������8d��MdJ�b7��j��Tmr*��0g۪��/V�2^r3U�� F\$����ߏyq��-�H�X�!�&x�Q_�ˋiz�K�R22ڥ,o���I��n�V��XQy#�h"��:�E����x7o$�3.':ݢ1�Dˑ�G�O�/L�b���3(ɱ�J}PKc�σ�f�-V�$a"a<(��<��Ӯ�a���9g\BU����ë �,�q��ǥ/�q� %#�Oj����J��aTԉS?�>+1>���j�.v9���j��6�g'�B� NNLe��e�I\A��R5��n�gm����|�N�~��̐U�eR^bY�BI�a���d��F+\�X����C���M .�_p��3C�Ǎ���KF���q������{��R��5�Nڕ�#�����p�sϏb�	�%=O��_��1*@C9\��A�NGu�)K��irD̡�G�Agg$���g�:I���V^?]�K�-P�_��j�H�X��Z����J �ސF���ؤ�ܘ�Ae�řӉj�h��o~�+��-�������)�J�s�Ji�Jf�x����(z���&�Fcr`���F e�%Ҙ����T��~������%i7�7�W��>�ASSS�Q#X�w±pɄ����������~�5a�̎���XT��{W@��9C� �|0Hђ��y��-�(�BZ�M<n<55w"�.����H�� ��=ј�n��%�����̎�O1���:��D�d�#a@��1�	���5n+<��ﾻ��ɷ�{pm�����p�u�f�b��J9��ɔ�����M��C�	�K��W�f%��C"���;��+TG��{*r�Ec�8�wW�T[ƵkԹ�8�����h�x=A�_"�&��e��d�sRH�KO�6��8�G�ݳ1�?W+p��#>}�v�/��?�Z�;�
��l�MK���=�	n��{���Ђ?��?s�p�hH�G�-; �8��+�/8�ڒ�?
��:St�sA"������6���^�F�N��ֆ�$�s��2cO�����^���Fu�SO����>���a���� H �`��JN�Ί~"<��?��?�����ꝏ[�|#dD<�8!];&�ڊUx5�r+�؇��]ĕ� �͘O�r-���������~4�C1N~`t���a���n�=[���V �e�6{�Ͻ�~��o��Z �:�Y�&�a}&��%������E����N�5��;�w3�E-b XA�ɢF�@����%&��j'�va��سgO�d�/� |P�����R���3DFGp��Db�i��^-�	�I�XF��$��:���c�Չ^M7���h,�T�'�T�$r�:y�]��^٬C���[b;%NhW�@��A�c٦&7��][�J;2�ɠ�8�<� .��Vb��aI)��6h�����T�42@m۾c��s޶�VH_9���w����o�s�6Mo�)/QS�N�*62N˾��pq� . ���uWK�T�J�$��WG��^�
��ʵ�����w��3�( ��b�b�Pn�bދ��r"�25��dL�sքƱ���_���z��#Gˀ�FB����B
��X�6�T.��蠀����t�ܓ�Jގ�T��+]��q醉�==k؁��ؾ�����fw���љЯ���m�����a�V�Ֆ���O��A�σ��4�ymCkY�q�&����ڷ��d`��
�q]S�sj����/ ��>S� ��T�p�bʊ�%U�����6@ޣ�p/WO��&Q ��6�?���PR�3,�'V	K����Vo.D�����"G���N�)3(
�``v+v!�F�w�*�Ă��ك���׼�78��2@�Oj�z>�ם��Ժ�m�|�}꣟��O�#?x�����ض�;�`i���M�;��,����l���$��X�� �Z���\îҲ�����7��v�������v���ע��4�b�����Ի�*��u�]9R���J��J����� ļ�������B�;`^!��Yد����Ғ �@�)2��-���H�tsp��P\�"�a��v���9%�� H^9�F��
�O�B ���Q^ �{����6��'�x��򃟴׽�v��=-�GIE8�wx���E� ޠ���D�i*�&ʹ���0>��O��s69qF��b�2x��,�� �:�0惫�//@���4�0�!�D;>�I*	�����&�
?1�ΐ�׆��5�R).��h<�Ԋ�^�8.��U;�>3�Ocu �Vɪ���3�C���2(��b�xQl+����������@. UjA�, JVI��g�*z@���R���V���{roVl�����ٌ	���;Q��A���r���ј��Z��o��������c�nٹ�LS�=�q��R|��ԕ+�{H�VjD�2�B��T`�7��W^	~$|.j>s=��Sp�H��ʹ�
�����.��}n�4��>.u@�\NN,�̦�x��b'f���є�V:9�= [t�@� aY�"qB�t\�xK�C�1��AɿP)� �W�|�'�*�z���|Ĭ6�Yi؅�m;N�l�S��ޯ���)��ōN;����ڠ]DE\cYǋM@2 �T%��-v����_�o�*�^�lW��B��^�1[=&/̏-���*F�J���>�X�J �+^�n�a�|ДWcB*X!X�}r��֞NZ�4�#r�t�U�([ϐ7�@�H�G�x7�������XY6�ex|>
��j������O4��w��t������ُ��z��2ʦ���9�T�F�{��h�c��Sk�:t�<�6��r�>����҉k��X*}^4Lx������#�8����+�Sc���}���?�$-?��w\π?6sIMJE꟭o��->E���[|��L_�NJsHY�._��V{�<�k�0��}r%1!�̫V����*�ʡ 	Q^GR���)l]��x`Z��گs��y�c��� ���o���ਕ���ݑ��LD״ޜL��R�+��杘6�&�<��Q�����1�L ��>�s��Џ�;>Y�`�Rߓ���G9����,��8�-�[@��V� ��xw�!4�p�/;a�N���[�KΰK/=�&�Kv���3S5�cXr߻�%����DrX��F�o-7I��W@L�ߚl���&���姩��r��Z#_j��=�H|���r q���ʷ[�ڐ6I?*䟵 �K>Z��_R�(O�����;��RV�%SH�.}cqS���}qU��6IH̊6X�]I�z>>$]�D�/%5��R����7�{����͛lbj2���\w����
{������3b�#\:kթ�����w�����*Z�&T����
q?��m_iE�C�'�(MWǍ�>�����/山��a	b��<�����	9�m��l��Y|�v��������9�7��2CC�'�.�W[.YV[��J��>���X���.U����xx�b��B�X!��6Gq�R'	�]+$T\�mD ��8�︎rp=y���(N�K;j���|�ө��F_�Sz?-lq��bf.�y�bD�U�C��,����$�{��Ӹ*����K�.���a��E��j�/4cy���b��n�풋ϳ�]fss-k�� Y�H���kw���h�h�9��43��+!yRx�P��J��an�9�F��	�;&{�Cn�}����K����&�v2-�QC�������M��i�Z���>:g[gϲ��<1��sP�#N�W� �}�-V��L�,�Sq�J$.S��D@ ��X�ճD��-p����%���(#վw�����H�Tj3��i��y�R�S-7�kN���j���ࢴ8���(Jn}�(4����^��D�}���o�z�r���m0^#�Z�**È��#���FO�jeҞ�7g_{��<�0�l��B7[703��1��Z����3�Tb<����o��Wh� �dFp�˹�l[?�[A��Q;��Z���RWxqP �wT$5�|�.ngs'�W��v�:h� Tu���g�D�F�'7e�"ba�NLa�Df8/���*	)����������1Y<�Q
Pe'�q��	I|g!(���ŕK� (��W�G "}1�䪦"qO�*ݭ6��A{U ק����p=�)�c�VMqഏkpm~�]��~�-\[ܳ'�M`��Xc+���zR�����1��6L���b(�����p�R6�N��@Kܼ�U̢�^�g�ev�;z���߹�����4�Sj�I;|���}���u7��]gY�4��b<Ƣ�/�8�� ��y߼$뙸�H:����\n�9�xUߊ��'��������M���vs�Њ"?f����>wb��'�:Ĩ01�h���	 ^�n���s������	[?��~� 	���cq�X &�^��^�X�8� *�-w 
�)~�J~����$�^zit�Q�@��K!^/������x~���8�w��{"�����M���{|�rJ۩���'ek�$��]ʅ�爣�t�RPEW�� �#��O��v��2(������n�#��$ƕ��MQ�p1�2���H��u�;!���>JGK�i�*�r�+��N�6	t"��"�h3�*T�gGpנ���2^�햔óճ���I�6�FN��X��^I�U��'m ���{yھ��w�G�.xS�Y�ͨ#�:�#q�^�(R�.?�8�w�%^�9�	\�{�����5��sZn��%�T������u\6�S�5�-kwI��-��0��NసVu*��rFT�]�I�"���ʑJ%j���ű�	�Q��N
P�  ����>�� G\v�����ߜOi�����+��"�/`��v���  ~�>�`�� m!3ɺ �.� Ĺ��`M`��T��K{9�� � �r_Tuc�����f��崝1�ܛό# ��*}.?S� ���r-��f��f$� �6����@9�񑏻���w υsy�<��&b�1�;�:���z�$��� @�b�3�����G����9�TX.%�N��2F-�AR�&Y��tлD�J�3ʯz��焇q�ˡnw��	Ot:�ҞRO��*�x�b����E�U{u�#Y�ДA�u�]�n#N���;t`�@����dح��a�΍p�ˢ�?�<�_�D���Ćdܒ�	�L�Z�3�� �D�X�$,\@���x�c��NΉ�R% . ��� h�� `D;��-�K,.�������m��s.`�m�x��q-H�5zv�E�JWʸ�+���u�I;��6p]ڦ�d�4 j���6 `l!�9%cýd�U\3@�̹\������fD{�� ��OWc���<S�XQ(�TO�������`֓�;b�S5k�p�u�<S��;�0*ktӆ�_��g�c�\}����9���uV�R��D_;�	R�TORE%�Ai��ԁ^R�h�@��ƌ�n�B�wB�b*���muc"5���kAIg'qKzE�(�1�<�(~ �u�� H`��`��y\������9'��J%�햛�cS��z��&j%k5J��ɖ���;��G�Y+��="�Mn���W@�� ��{,�0u�҆�Dn?�;:�K�'�����쾺3�	��BC!�ø3�(s@���9�c/�<+�hh�D%��$��Y�� ����/s�Ϝ�=�N� J��xp> H[�tʊ����q�@��sƐ�܇y�J�|T2���U���O�c�#��VF;qb|��*1���޵�����C� 6>�'����G�.���).	s�����ǣv���so�I{�-W��dhC�n��R�[lrb�-,�y&���	c���G%F�A�#	W�S����|�Oگ�. �������9j�C",��]�*�{ch�9�n))U˕�g9 �lpR,�t���*E�%݊&��E���a�8Y����t�,UP�N��]�;`{�O�=I���~�v۱}6֜�v�V�۬�[���1��s�>aϏ&�����A��Ȋ�o�	q�qg�XIO�o�	 �ɨx{�ѽ!D28�y ��3D)U�P2����K[�r�&��ui��^����W�'O�B�űÙ�8SUX��T9^_�O�6-T&������㽌\���r	 �pќ#��r�p>=���4��kr,��o~����I{�'����b#�06����H9O�gq�P!�v]�)��UJ�5�l��	��bpu�[8f�v��O�N�ԯ�����a���\���V�6D��v�|e���@ء�^̋���xx?t�����P�Yv	��}�Oi�������N�'��.��J��KY�Z�U�?��N��w�]�	�B�=��.���jb�kP09`Y�e ����鑊�vSQ����!;��vÍ�И�a�[�Ul~�p���p�eu�'�·*�_�\�
�3�f�͸*��W�B� ~��+_g<�^g��H���4�p,|~c�s�V��3���(��Z�<x�'�����N\���k�����f�zCB\�<+Tq�X��Q &�����9G�>��NT0R�p�Bh[��8��~P�	`�g�ϱ�j,�K����5.�˜��8*�>�y�kȅϯ�����c��-�a�զ�9n�G�m��?f���vɥׄ��u��Zb�z7��"�$ϙ��|7�օ�Ah���}��T\�gc��O�m�k2y6��4/�!K��p%�N�ֺ�r�SI��ݥ��%I2	M��o?=r  �V�5$�*�c�9�ゃ�k����K,�$�L��0&?�0]��2�(Z�����q-���B���"7�o�-a��ڑ�lfS)<�N�QˀXE=#wrP^? �����&���r�J�˱��G8+���� ��=L*��x&;�	�p<�l���\ �de|y��$�ȆH)��\�x�<s 
�gŽ8O�)8y%a�E{T6_ �v�0����617��ע��ƫjJ���C�i�Wp���h<���W�1��1�<��8T�)�8c+uc�x�,�+m�m|��d�L��T%��gB��ӆ!O�u���~��b�l�X�1�O��b�>����w���֨W�~����v��o����R�<���`�~�T@�� ~�y�KV�"���j<4��K��ld|׫M��y��F��#�e�+r��Zµn'�R�s	�!p����v�,����.�k����)�� ��o�ǔ�c�P���cLbb2�$���K�����U��7p����8pЧ?��\^"�(gu�	�,%��v+�;����vϧ?o�yͭ1�O�Ӵ�MC���:�����[��0F,x9������?�X�Ð�X��])�����(%�:��s#LD&(�v ,�ǳи�:
�г���t˼�N�$��㸮T
����C�^q����7��g@�k�l ���o��y1�|/� s��.��`^z��IZ�pO�Oq��2�%�}%Y�_��I��gmb���U�z�}qf��/~�0s�fd/(��u��U�am���S�Q��ԩ/�����=�������T�t+'ӱ��f�oe%�� K�qw�qG�����!)in���{�9I�+{�|đ� o0HA/�S� �1e�W�B���=7I�2@��T�+�%]�*�0���Xc.�i�p�<Q�s��+k\p�E�E���!
�O�!:&�@
7C� 
�]D�4�p��	1F�ǽH�|�7Dq�kHL�V̆��g��'�\�&O- FXDO<f\tVh5�8eN[_�����~�H��s&()��p�^���s�3�OARoh2KO�݅(p�2�
|� 4һ�;���>�d\��(	��) 7��k'5��?�%N^��?�M�`�'����"����K���2
�~�W�\����MB���`L7qc
~Иs��q�0���$$�D!��j=�:O�M�x"�#+��j�yZ�	�0s;AWO4�-# �Fla�y�k_�����7���_��h$��<|$����{���o����iH0���#�y��`n�����ճ�z�W����{G��J���R�8���-���XE�`�����tǄ��Q���&5�V�X<tL�*E�l &�o��oG���^�:���?��k���o�Piw*& )�L��τ�|�.��t�𢳣:��l���"��,�{&9ur��J?��:�/����o4Y']�<Ε�����k  �X%��\�+xC�S�%�{�I4=�-�M%��.�N�~s����w��T	>���@��~kj��W�s}��tw��i�)��kjQ���8E ���&�!�u-�Qu�I94��q�&�st��W�K�K�ubn>����NEIy��;m��h[1x�"�����Q6�'�O�^ �+�XA�"� E��Cf|��К�3���*<�Z�瞽!�k=��Q�^������C�k���@���ђ�p���X�ʅL�ո��K���1=��
~�|�m��tϋ_��o��A;:�����>f��[��.��!#�w+iaxn��p��mb*v����{���Mw�y�i�a�3�r�R��rN*���YC���3����E��G��G�����=�h�c�}"�aM�H=����x�s�
�+�&?�ݑ��Z�i��%�(oȟ�=n�ʵ����@)/���,JUޖ��R�/N,��J�����a�z���^���I�T>�k=�����,X��h�R5��nD�6���U��;��}v�ȂMLZ��C{�S�c�Uצ^���h�;��^��F�����_��CG�J��ɥ�'�B� ���1>��&�ׄ{����o�b����jkN0!�ݩ5vQ�&jUk/�^�'C7s�aW`p����bO��B�iBH��$B�HG�%�R�����ϸ�� ;��� � 2���}�}�*��g`b&kv�ۛ��v�%����1`��Y��8���'^p��][���o�I�*���Ӱ�x�����N�c��ŰW��W��ڤW�J�H,�P`Qz�ܠw��QM��}_�F�߆����v�����1)��u=��k��|��~�-������^m�c��J�i+��9��*���I���DVmrz��Aj��*�5/��~��������q��m�\���P����f>c�Fs`^+i�ThzN��jozӛ"|��}��2.�%T��n$)�5��M	]�ʪ�,TZ��X��<`�6g�Q�̑)�I�_�.jI���S��4b�2A�β#��t
�I<7��g+w��,ƀ1��Yq�pw�}w�0����-G��܀��D�����Rb[wL�� }��۱#�6�y{x0-�7�<��-�Z醋f}*�AkA���5^I�R
LWg��������T'��vع{���?�Ή��'�mj:K�Z)�֤��b�@�D
�6*OT� ����ƜB�yEj�0:+镘6y�h��+�א���_hp�{t|&��C�F6�iH��j/� ��l�F�L�ð�J=Ile�؉����DW��Y�pź�@��)b���$���x8Oj����%DN;6ޡ��쑇�N��Ѱv�Px�m����ID]���Jv��nu܆���~��l�=[��z	�p���ѣ���=�����*�n��F:�险 IS����K���"y�H�º7b=���+jL_�G��C�k�pˀ/x!5��aĠ'�D��M�eWP�*�,��̛&�%�n
Lv�P���N��ɸ��������4K3X�(S��qH�|Fe��d�fgH�++�z�w��Q1���g�$B`��J���Ur<�B����lM�7�}��k�a�MTÎ����I3�N���eJ�c��X�z�σlэN�A�l�L�6�@{z��������]�G�o��]`�]���%_>���zLeI>a��T#RN�fP
(Y|/?ie��3�AZ��Y��>��0�'=��G��s��K������S�k��hRD�7���+� ��EQ;R_x_\����^~� ��IB�) �?��?���>�яFu�9�3p�8��.���Mo��`f�q��ܿhS;-��lf�|�zb�3a� �M��i+(m4H=\<�67h����nVA���ٰ~�n��Ԍu��ӭL�x��>N��f��J����XC�h���Ry����3:]�{Yìk�<X>��OE��t�rS�a�����e8�1+H���}B~�5ہq��ڃp��q��[7�F1B�R|\6����Y\ ���y�\A��c{�SH�p+y����z�1�@[ ��N+� {p�|��d �f �2b�Bh�p�.�ռ�\��a�;bm�����\?���ؠg7��\�
k(H�ݬ���d��S���歜�����vn�f�o�7��pl�q��rC������;�c��^��UKF}T������䋷A�;�D�3�	�꣇-�R)|^���J�Y���_�L��Q;Yp��w'����+������z�������=��w�;�K_�R{���B�ey�h��So�;�D���$:jIe��{�b,@��'73��#ùS6�诺�q��қ�Rܰo����mг��:���4�`Ǐ��v�F-s��t�T �ik^�%7<�v��8�i���j�u�}�=k��W��r;`��B
�Cc>^Q>�V���E�D�*I[�
k�y���}��T�]-W�n�j����	�y]�#��V;A�6�w��."���h�"����9�o�v-�E���+�J~����?��N��R�U��ꂼ�dR
��> ��ІFhx��l�&'6�wz����-;xpq]�����'��z�S�ݍz� ���Ӧ�mo{���c���I���Z,��l�lz�Lkf�Ըa%�'��T�eyT�
C�o�u"����3�>�$jSHҲ�	�A���w�ԧ�QT:S��@���D�:I��D�Aة#�IT��J�ȳ�y6�GwIE�� �+6���?�{|������y���}�I��
����$����f�mE�h�j2�w6�9۶���0/)����I�C��½&��J2��RF9=<��
1��J�$�J��g�����S�7�'6h�i��N�Bnz�@$��V'���k���g��/<C�1ĵZU{|�U&f������z�b�F�T�6vDӱ���Cs ����f����������/^c�S�#q��-˭<#8߫E�6�^ .�֟v�̱.qW��y���'�H�Ġ��^�je��8"Kv�
�KΉ:٣O�%��Q����X}�+���s W>+K�t5R���!:#`�w��X��F/��"��8�Z�G�_.��L��#����]x��v�M/�͛C��cG�
�KF�0q�R�3�� ��<n��9o��mp�]��'.bra&�c�R�@6 x��i*��;�T�3�1�J˶l��c'��?�����+��Ѷ���`��-�N[y*����n�lO;mG\D�¬��y���ڽ���ɵM���`��d�)Xs>�]�
��L*<���'�e��e0�Y�$O�ߍZ�Ռ�xN�UNcxa�"�~��N�Z�}AVS��а'�Tt�D����1��j�XDՀ:]��#�b�0a������薆h0)q����.�Ї>sI�d<\��[����8�سx\7|�e�t��G?�����7����s�ґX#�رV>Lr�
��˃����76�c�q`d�/�`�qL �q$��mг�2Õſjd��������~�ؓ���W�������R
@�Uo��a�#7�l��������7�9d�(�>p_#�Ǒ���D�:�%%Q���8c�8�R�zݰ�Q�(>�s� �rM/�gx��:�j�Z�]�3@(ƥ� 湏�m^|Af ܇���H���dm��ݞ�:;~~������H�z��*�΀������_�r�.�|�!���@Qe^��-ڎ��؁}���){�˯��\zA��ь��F�����
g���p�
���:�Z�X*�����J��#@�C�E�|�7h�~���`�K�G��0�N��'���}�{�lv���P<���Z��zc>O�s6x��|H��k��62kw����R�]|�����-�t 1O1�Д'VH�7�+Me1�;8'M� ^Z*i�h���#hI�tC���F�ވ�����Ύ�,��*�*��C���w ��?��_(���J� �<j���/�F9v>���^�̫2�y�4�_��6w��Ϻ:؈���'��l��4��G�%y}�n:�М�!���f�9}�}�} 6}#��6�ڠg%�[J�i��k������m��>�P�yr&`C3p���pV)i���a}0�J��}��G׶V+� w�_%��^SPG���I�4��aV�I��UN���7��0�!�s���+>�Ւ����r�i��t�h-�U+U�(n��&{�UW�J��2���]�݄���p���۫���>��A ��j�](�������$�����I��]aמ��tI)j�;�o�2l�ਢ�s���K=1���sx.��=+�u���Xk.�/ʕĦ��A�<߾�бhWR� �S!X'F�Yw�+�ֲ�Z��r1�E�)g�`>�L�I0j��)Ҁ:�"��{P���8��a�9B��lujvr
�%9a.i�N��I;>�E�5��c��j����HUdP�T7L��n�q
C���|�)= �M���n�\Vy�RL�A�Ӌ����z��J���ѧ�~��]�v�o�˟^l��#sV%�`���k<&��{��MP1�|�
��J��A�l$8�t��r5����t�xo��F{��O��G��l���c�@��ԗi2���jL��QM���y�Y+W]uU/�?��)��d��mF�W1�
�� X�u�W��b`� b�}�.��Ҫ�Q�t���Z�10�1@|���X���5���)��p� 0�p��Q���������NBf�.��}�ԓRT��D�Und��>9U������9gO�UW�g'�"�[�N�����@�j���?ʋ�9~���S2δ_~����.j�LS&�����Z���m�4k�]w�]�ޫ���+��18��LF>}��k\0 
SsG�%�W�<��4�~R���p��L��t��ž��RQp-�
�J	g���>�ǹ���#��+������f1���Pi,�b���Wg ~���j��-�������㚨-H�9SUd՗�o�_��/��m"�`A����j׽�;����N�s'�����7�3 p��FE�� �H�{"��HH.6���£���T+�x��a�7虢��f��5���Vg�R�f��b���>g�ݶy�:Lj�,9)Jq�v"x+D�x}H���d� ���+12
ʐ���WN5��H��6����\e�P����7����S=MW����c�[�� (�c���L��>��z�Ii�=��tU�ŗR	3ދ��<���&�7�#�Xd7Mc1�>�&�K�i�Ҥݲ��ħ��� *��ih��{U�b�!|�ѡo�=[)�}�lwb�j@\��}��
�;1����f��)]�l�rukTE���h̋�[�ը>T)4�-~A�]T�Hă.��u,�[��:xCls�F��0;0���	�� �F�p>�y��=�*m�g�(S�F�(�OI}xG�r2����a�ޱ���y�,�U�6՘=���h�����vp�!�P�
�]�|ʞz�m���I�:c�&
�JqStPlT>e�j�A<x�	�VLH�td�6�YEi)���*�Arl��C���|���g��VZ���g�i�]w��>�b���	�\�ienm�{婴n�qz��Tд�-�I�trV��NO� f�X�A��?����TWk�[Z'��Ϝ��I��48P}�-6\��AyAh�9:��~�Q{�����.�����'�SOcF�Vc1�HFϵu�i�,%�zE={nj�Oe	��>���#�A��*����X,!�A�l���mƥ�5��۠�C�
�����}�o��O��B��n+��ö{����Q�s��:�vO.J��@q��cJR���{H���[#�9�^'�(��D�LAn�(���@�Z��G�)��8`�
����O8���1	��� mҶ�R��� ��N\��.�#���&��q"�X@[U2'>�
ߠz6SVA���$-���CZX���� [f*<�p,?\Ӓdb �Đu:�k[�ֽ�0je^�w^Z�I-*�$���b=�y�X��U��tu��OY'�5��)�2Р����uvyNЋ��|uoo������rG��V_<'����hյZ�w��B�~�Ⱦp,���#Mb�����$��?�+©�'j�zUF��;@z�6�YI��j\X�额q�Vۺ�b��ޚ�s��]v�U����p�R?�"	��Մ������5���$�� AN1j��O���H6]���Tii?a�DH��Zn~ ����V�(h�!XMt��z��v�^�<���޳c6�W_n��-�Ś�j���?|������ر� {)��HO���"�̠rV�5� ڢ����}�7h���T�%��`�mˌ����[n}~`[�a=um��67_�a�Ie&�#N��)=%�����n7�}J\�d�Mѷ����ٽ*B@*ψ�qN *�Yb�|�Ȩ5_���	���#E��:?D�{Pw��� �kt�?z ����s��f�!�e�v������	�N,�Ƈ&M���U��N�/<��\$�`%����ʡ�ngbX���Ǫ�N����x��2ܩ���U�^?��\��jh9��Y��^�u�l�F&�X�`��;��3�w�Xu#m����v�pÚ��=�$>�oV_��,P�aD�K�A��t˒֚����^Y�y5�O
�ϕ﫶g���ѫcAx���C��s�A�+���*�E]Bw�XuZ�Zu�lG9B�+� ����3�]&�U��a�p�jK�d�)�C���m�����+���w�����|�}�O�(�@���rf�����%t2B��B�op�0¦^-�:��I��l�\��˗_�o�*��Q��4��R��R�Y)h��~Jr%��,�۵!�o]�x�R�O${MT�q �g�}N����=ީ�NY���$���nB3˨ۺa�����R;���?����z�.��j۱����5�;rׯ�t��Y�~>a��A�+I���F�x_d����g�<�mO�XOb*{�D��I��ז���XPH�ة~��Y�/�?9xP�}U��X03�Ȫ�N�����rq���\�R7x_[��	臹wr��}�l�鿱���y���+���6=���漕p*��=�W)�}�y%( "@ݿݍ.p��K(�fc��}�y��(�m�O�4�7��Jm��/��;�����c~���,^��k�_c�-�1Cޤ�ڻ�~�ܯ˓�4�O},~�w�G6������W��N�ju"���G��fX�����o���g�]��b;��K��8����X��{���4�Q{b��=0|<��yU�O/�lW�>@��N�my#�h6�F��=7�XHe��j����@����6-�Vd�S�s�
x�,H���ي�-�O�V��(��|�-Λ�����|�^�����ZDZ-�]^��r5F�� ����Z������-�]�{F�|𵨓��pN��o)�Q *p%�����n���9C�4NF'��QB� ��Ԭ��KI|��+�&Jm�s��j�� ���u�sk��F�@x-�%L1=��LZ��i����'?g�~h���E��isI#\)e�M�D������ƶ��n�����o._�] -����yK6�`+�� ܩ�}l,�`)�����ʸP*���`�����a�^Oʥ��2p)�Z��T�c��I��`��*�D-�5�f��܍��\Wk-8�n���y{��OU�uߗ�|Ggx�2��D%0\ts��ߋ�e����w��'����ˌ��7�4�t�t����`��`F����n������Y#%]��t��z� ����D�2y���*�Ν�2����TT$�U+i]��˕ؿ$5K�6Ab�̅/�%����e17Mx���>�J;f���K�r�C�j�+&	ދ���jSM��_���H ��D���-u�z(��6��v��/�ZKlb�j;��bg��۪�vb�8��.8i�9cX�DuD7^�T=JK`��h�\o�r~��p%�㊟ך�{ݜcNY����a�e�Q�l��C��1�x�t	�xO7<��a :f܊�LO��rX#1�	�-*U"`x#w�_�gG���{��X�e�ڭ�u�i���b�F�Ϭ&Ղ|��LNs��KI#�r� g`!�TCT��ҝ���V���?ߊxLǈ������^W\qE�
#O��z�.D������ܞt�Өݍ�a�������'�r{r-�Y����2����Qi��C{������7��]x���X��C��7��K���:Ҥ�c&ʎ��wm� O�!��:��2����NR���.�kb�������� 5I����r��uXZ�b��ü$L�C�_��?�jfړ�FQ��=���_m��/9��^�Z�
�Нw�Ҿ��'챽Ǭޘ�fk޺j����Qc��h��<�Iֶa�z�O0XA`��H��0��
�k�'���A����7]�.�0Z���Du��k�F�J�lg�}v ��ǜ��*�' F%J��).�)L�)�C��Т�1��n��6�����x�w��gϞ���/y�/G�6�j�	��㜤� )Oe�~�m���.;�^��Kl��h�Fh��l��1=/a�|cґ�G����M���G�~Q�Nu��2����+����'+�(/n��A*3$�z�68鰓X���9ߓAx3Nt�3���#(�,
mPK,�6����a�fw����Z��d��"�i�����(id�ն=�ϱ_������7	��lۼ�fǏ�#��k+V�Xb�����P$�*�DMb��.�,F�RH��ɚ+}�c�@���7p
�����$ot��"���0�SS�5VGt:\� ��v�M7�ƞ�Gkr"(!��o*�;�������P5��ߒ�g��뮻b"旼�%��W�"ޗ�R�q��b��~�R��,�O����-��^�[��T���F�h|}9\r���,�c)Z���~�䋤c�b�l���A�������-����v*���>��������Wx]�w���뢟n�����̆y��,� i��(z_�( 0^bj�wۻ�h�O�$'��1�O�Լ��� 9���P¨T�F�w��ٳ9zE|��='���/'�ru��@Y	x�/8B�0$v��/}�KG��e[�� ����_p˔bS Z�ت��涬`��q�0����m�{�����}�=��S���J�̐��ΰ�$աc�(�Q?N:��P���J"�s�=�^���/�rs��2���>�у<!�d{����)�ͻ�~9�V��f�R�ӴV˔�?|�)+_W��Zf��"~�x<0D���6�1/E7mǪ%���K�r_�Iu~�si�K���dƻ~�`�+�8�����t`��~��n��Г$���uJ��-ñ<��#�L���g�G�17�s�OJH����~T�W9��4b��Rq�T׷�h��G��"}2��)�I�[���Cf׬�J�����w�"�|�gon$݁y���3,1l?��'��R`&Y&#��V'�jWVs���;��*a,��G����0�m'����l�D˶��;������<RD+���^�M��z�z�9\)�õ�R79��L���J]�q�6)@ə��ԗ#:�{�qn��U�P�8f՞��X�����ʓW���fl���:��`ɔ[���a{�5W�A ��x��hx��I@'}.`�\��܋_��8����IKW��?�S?��cء0 ���cy0��a�<��|�3C�/�wa�,����w�=����c&����2���aB#� ���{�>a����G~z|�R���Y��1��8�(P��n4��� �Q�
��`���{@8U��r�23���/��[� u��Ja2�ݜ�qaR3�}�n��e�}!��ϯ:�=h�ő�d����'$��t�'���Y�U	�>�po��N}���ə��ONTs	�q�����Tع$*�$jb���[:�|�[��{�id��)�r��$΅X��m}?��	�pȾ���>���h8����;ڶ�:�\{�tû/)=+ 2�06���	�.��(�mw�����k��Q5F�+��2�� 0�l���1Q���Nػ�o���3��y�e[o�˽��^���[qΈ����ΞC�Mn��WLȭ����~$}�~�;*�����q�u���9�~~:�Evm�nZ���ޭ��׉zǩ��x�7�Y��?�A/���׽n�v�����K�
?�^�8�Z`ﭷ�:탹9o`��cp>�{ؐ���
7�|s��*8�O,{�XjG���� ��r3Pzn�|�}~CJ����w\|�nL,�������7�G�%��q�q���"`�2ep���g�Y3��!�9��J��o���1	=����~f��M2WT���J��q6<p�C鯾�t���:�6v�����P��l.�n�A7�[k)[�[7QF���8�=]�p����h����r��zʠUp߭\���y�G��zg��b
S{l:�L��섃�g&���ի��,�O�1}��ۋ�@����u�r��9��m����"5�0;n�`�m��n��c���aTY�)}���D��kw�-����&[l� ����T��׋ 9�4�7��w��&���5��0 �[o��m�\��6�ݥtp�ĵ(ӃS���F7=`����ݕ�3wB���X�N�d�J��Zݏ�M�� 7`����������;�i�F�"�Hl���z9,���T.	��>���旁p �9&����Q�;�nq������4����@t�w��/D�$�(�iYII}f��er^���"]e��`~PU1���y����|B�LRC�h���kl�	'�
d�,�
0�c�-�&���Ғ;HKt����u����v������ݻ���t�=/^9�m�	g�h2]ty�����t�iAZL"o������̛�*W `��g^��l�) w7gyj�/�NR�*�<��@��P��T��!3D~�F�ϚBv`j�޺�1Q1P5P%>�&Xiky��"==VǚŊ�?��פ)2���e.�.=
gBh��X�2UҔkPڽ�NS�?�$?+�^DƵ�z�����u]Ϝ���@|� �VZ��=�I��2�k{i�����d�ʢ��]ߠEX�]#:�׌���*��\r��bV�̒`Ɵ�ɟx9X
����o�?��OA���� ��� 6�͑Z���'hͩ�3�������F{��Z�n+��S�+ƝZ��ˢ1�㼳�q���4D�q���(�VC����x�)�iB�c���(�x�����L�W\�R��ot�,���<Nn�Ml͠����F�&Mz.n��0�|v:�HJ����:�w�r1�k:"D���@7;���C���ܸ����x4q�Y6_g~e�L-:)�a�c�Y��ô�������eS��T�t��j�8�ndǇ��d�� �=��)𬨦P�h�v0��ݛ��o��t���7�������0�qݜ�6\E����X5N����6�������^mV���TL�S�M@�aX�g��J����4��4[+#��Cs)R�eb�k�ήk�B�6�� �:�u���O�{��g�p��X�Re�0F�$��5�\N6kM�r!{ՅM�?���1C�5���x�);��x;e�h�9.���bn�k��֣�!O{2r5~R��f�T�Kf�h놌�C"�����%X�i�$7�$e���&`��,��g0�^{�4u	6~C�����+L�`��` �t��m�:��al��Z�r2��Fo��G�������j5L@�$���ÃE��]�yԱ)p�=��WC�ѝO']Q�0�����`g`�"?`�f�[wh�_۠��R�/��Yh��d7�7��)��� �ڌW�U�&<aM7%(ޘl�&-���U����	�%�w��`Ǌ/f*W�'��@a@�!��+;(�
�^#cR��D`'�\���y��I�Z��ʺI~�2���r!����*���SG�y(_1��?�����o��-�T����y�SGdfХg+r�9('��9󩗳#�	sϵ,-7�l�����^�� �XTה�C��`q� l�L8_C��,�&�ՙe�u%h`e��05��Ɠ\�&����q����&���Ν�Ƭ7�wҀb�_z�F���(�!�Yk���E��/�y ��d:�S��׌�,�M߃�|/U1�ħB��^��ċ�T�Mv1���������X@@��x�K_�{���Nf�	��Wjة{��>jU�~�4 ����f]�E$\�i aDv3d&��sB�$�`�Y1/GuB7���L�z��1-�E6>�'��I��?���/��/�Q�����漊���G���ƄMjV�M��M=F�0v�YXX�L96X���&u�Ė��s�i�S���ߑ	ov�0��]��ls�曞좲�Q��zn�Rf���-:�ڰ�ONIU"���F��0j;��Rׁӯ�0iR�9�7V�:C7�R�Ә�w�^70�pV�{9��N�(;�r��4�����{���^���:�(�iH�s�� U�
�E��`�M� �|Î����V��ͅ�7i"�f4�;�j`�,�,g���,��<S��l[,-�=@��ݘ�h��g7v���|e��'��j��>&����h�NV4�ko��38�βobc.��q���zӨrF\����`ves_u����m�ct��p�MZ�K�A,?E���ϵ%4�����k���{DǍf�F���w���h��3s�����?O�*C�t< �m�N�U}+c1���fl\NS��q�{] \�#��S�z���*[Tl2r���r!Q:�dZPؚ�KD�����U���~�{�s	H��7���Ƙ%86 ���񌎘�9b�p��G;��!���3;�\-��C��iV�`V�=�W�t�y��w�!�`b��k�R���s�Ygo�EY90M�{Ӿ��^�*7�tӷ���t� �y�c.H^t��ڄ����ܕ����w�K�R�������=�
��t�y;�y{v�]����8�ԛB�`�n�)�{�����t`ߡ����vl�k��Ҏ��}�:3��B,AG��rz�����ޞ��=�q��V��9��L�^r���p&�H�)��BsF=���Vc!{�:�9;ܹc)]u�S��h��Y�ày���r����ӏn����ђz��+.K�G��j�QҘ�"�{�k�������<����5��\�']r�cz���MtG�M���O����v�����a����.��ϑ���ݬQT1���V�������}����;۷��'^�ce��j�*�ܾ3�|]�s����[��H�:5D��ID�����[�n�N�',gg�g����{����$&�:�C�ػ19ֳ}�N�\��I���1I���Xh��������+.�Z8#ӧ�a���}z]�|�h~�[�?�=��v�m�m�3vs�� ���MjB���AP�� e��Q^���s�Hm�B�򖷤?��?���w��镯|�w��H͓�Dq��(��у��o���FI��ǋa�J�[����E�xvO3��qV�j�*5�$�9��$�5���`���7�"=�9?al���*ؿ��vdlhh�뎝+&��������?�A��m ��=�)����
�L'��Pڶ��:u�E��qR�x)������ޟ����r�������}B���~K:��mv�5��^�Nfs�%����t�?H��;�o*Lc0�u������ғ�|L�/vlْZ��Y+OVӶ���߹#����?��H�{�X��_v}z�k^h�q6�:���n������O����L+X�k��	�����v�*���t�u'��c�q��*>�_|��?���j ` 5�ϯ�ӿ���O?��K��u _���<��csxם��o���j��v�];�W^����/{zZږu�uX�v�D
��߳绔�������7��Z����7���ڕk(8�� [[?���qpUv��y�_���]���²}!����o���9m`�5[��m��5���(�/~�o����-�y�^�����;�fK�s��.t���瞫R��ۇ�_���TW��yn�L�7M�ұ�l�i����d���կv'k�+�FK�L2�@9�d*Qx-B�ގmM5f�Js��������@�@ �����).�S��uf����ɍ���t���Ä�Fe�0Ĉ���E�A��ʰ��7�t�O2C:���⃉Ԑ�W,;���#�!�����[3�ܮ���{�8�y�##g(~�c� =�����Y����t衽�k����M���1�]|ۙ��:Bǘ��`�}֊��e��iea�30:�P8{q�L�V�껲��+7���g��{��ťIZƙ1�a��@���R/8xwN��Xp�_Z�Z�6>ҋ.ܕο`[Z\�}���gυi߾�n/�+�}�bڿo�m�����$j瞳�X�Yimx���L�+;L���}G�l���x����s�MȏL�䒦��/�s�X����<ώ�fﭥm��2�ٰcV�%w^��s_ ֖��=�3��ڈE�w�z:��rmt8u!�Hq�&�� �m5���`Q������Ε�K�;w���&������G�`���ׇ������w��cǢ�k*����{�=���\��=hb���d��c�K�&8V�wl%؏����w���0mhl���Ǚ��si)�d��k"��57'�Μ���2G;�1k���dSM֎"	�j���s?�s����8_�?��F)��Ϊh
%y�E|_Z��R�-X@M�2g�8��j���h���wZ>�i�Eg\�L���.��0�
fw�u�1��א��pF� ��rSq(>��F��D��]�z�� ,Db�9���w��_��4K2غ\�X�Ԑ�@b�ǉ]G�F,p^ٱ����4X\p���]{�=�ܛ���Ϧ���<|�IO~\��T�ڝBkn/���7�wpݓN0#,���T��|�[���HKۗ�EoOW^uYڱۘ�;kvHM`;]��J���T`|�onM?�����祧=�t��%�\�9Č���QV�D�����Ӿ���}S��������fl�{nK���µ~���� V���i���ih�S7|5�r��5�S��.�e�ԫ�'nӦL"���@�+t0؞�����w��}[/���������v}�=�^�Z��YY�vC��m-���;�}�>����uO�:]xɹn*@��:i?�����:;�*ZZ���7nN��v�k?qՅ�k���pSHi��2��",Uǳ���Nnڿ�7�J7~�oS׮钋/HW_uiZ��w|���&� 4�b���?���a�f�������A��>��?�t�y;�ֽ��y��Y��<T�eS��L�uwJrM'[�d�!b�)l0�}���;  �$e���ou�x�^g��������<զ�m}�(㖡��vk�I@Dx�v��=F�7�҉�[���舜*�Y2���w�c�w�d�r�25p�y�v7C�(���Ka��FdV�YV�����X�DH�Ƭ�A�N>yI���P���*��"�b�����,�}`�1�>ے�*<����=���ƺ�����ϸ:������{�Ys�0@XXr��`���rE9�y(�G>�����t�w�sU��O>+������W�pj�d�f堟��J������o�f���{[��M?0��۞^������Zc���3]J�Rv9��D�Ů}�a��?�����|��I�Ȼ�yOO��S�s�n�Kf�\�R8��������������L�?K�ݷ��ql |iz�~%��ϼ8��Y�z��׺�I�(�L�կ}#������������Q���_���o��0�N��~�f��xT6!][/��[��O�����X&�~�^�^��Wÿ �&�lnM�3�<"���q�������|6����M{|�M�}���[��7�s�s�	%;s7��ܷaZ
� t!撾��/���_ߖ�}��3YL�9'���_�~��ޅö�g�~���X�6[�ϭ�ݟ��~{�䧿��eb�����_}ëҥ�{�=��L��n�� ��l�;�\��/��j�F'?"���l�z�����Nn�U�H�����D!m�������l6�p��}9�-�Z��3p~�*�5Z>���mm�}�<L)�j�i/~�En(?� 3����R�)+�4�a\��&��ᆙA�Y��|�C4�¼�ı�I!�ɟ��������n��
2��Um ܊��9Fu�̈��m�,���ݾ���s�1��N�}������ie��tۭ&�׾��t������jKS;��Fͥ� 	�1����}���M������|���L�_��t���9�r��]��.�[�X�>��/�>�۟Ɗ�b���}0H�x��M|��Ya��	�*nO�z�uS���nL��vȄÂ-�s��>����g~#��k^a,|��q�s��hB=�ή��o�bZ��������a��ᓷ�]g>]���`.9�Ф*ܴ��Z#������_�n�X[pG�n9����䟦�_v�;��3��L@.��u�'>���?�t�@�7X�̯?~���%�=1����gɜ��s�Y93�&ﬤ[~x_z�{?����E깣���t_z��h���ڼo�=A'��,8�h�Z@��u2}�+w��i}������K�Y�??�쬍���������7��`��JkƦo��W�ܟqM-�h�?��Ϥk�{F��1O�}�͝��f���3�:�&,��)�O;A�v^�5��[���o@�=+|��/ RMt��p�?��ϟ1�g	^Q���"ܐ}YF� �F ���O�[��F���َ2L�K+���w=���ȷ���/В�M6��cp3$[���H3=I$�M06�����G?�Q�j 3�;��_�r��}=	�@�H��I�A2VU:�!��Vs�=x�����T�r�	�����z�(zg�mw����~�Ύt�}�|���~�m�o{� x�c�z`-=��aS��H/~ɥ�{\�����c܇:���0=�qW��.�A:��!b����t�}�l��I/�k���.cav��('X�]w�7 YN�\�Tcaw{����ko��>��]隧</]{��y��84��P�m���xMZ?|K"�r��NS�/J���~��������[��_���-=���٦��KLwl����-y�k��ք�!�0پ�"�d�Ԙ�iI��, �k5�}h���K��ړ�x��{�y_|�9i��a�׮����_n >rf� ߷apv�ѭl�[ץ[{w�ZX^��`���M�S�v}z��c���y�����G0ƾ�.{���os{��2]asp�	�U�OI/{�N[{�j݄����Qz�������Y��'<)=��m���*�g":���g���j,���RK���w��Ɩ�t��ķoK�{����9w̕M���m��~� |��!�2f�i�9
ႍ����'?ُ�}^����U8+�Dż���o|cZF��������	����:�`��{�= ��`m���D���iˍ3�'C���R�}�.�8�\�X�*֝7���	��H,J�1�0gl=H���8���JkH4��g�� ˎ�0�hw�)C������8�$r� �
MS�����y�����_�m�/��I�7�*o��u����)�f���$�c�Է{^Z�Ą!y�}gүy�y$l��6�!�xki۲���*=���LO���.��xW(����ܟ|I�'/4�u���.�n0�=���%D����e\�F��^}�3|V�����H{ο��m�1�����Cv���HYIW_�ܴ���;�{�%��/6�Z�ݻ.N�{�����Ҡ;p��ֆ��+�N������v��f��"c�}�����r��@���u����⍴z���򫍑ߞ��w?�g���>���i���t����=+�֧�&d�<P���g�8�oH��zz�ŏI������� ���_~��ߡtnS%�X`>���Dx哯J���-����<-\c������'�N��T^�P�8/p�l�����g��o��w.���g��;�\uͳ��������6pX.�����级>���_�YyT~k������0ը!�0�#��+��}�2(����I�H@�d��s��9��h8�L����a:w��UD��}���������@(F<�D �+;��g=��6���"8
E�5n��g�
&�����d���.��ff�X�Wǅ�������v4sB�l� ԱNv�J̋��^�Nھ��OT�"Z�ӵ�ޖ.X����O	F�I�=�H�];�2}�C�P/K�lm{eg��Q{M������3U߫XFUM���6u�0-�c4,�Jc�;���o�(������ٿ9*킁ނ�gl�ۖWҶ�(���z��⒛P�Fa�E?���"a�Z�<-~y����bJj�d�K��F���a���:��AG�3�����+9�7�ذhs3�cO�q�� �ޘ��E�@t�r���X �Ѹ�����\n;ǎS�5M��������ߎthx��υ�<#*k�vb&|�&��\^X���HR��wβ���!*�fI��{6�6�E�ڗ0u��z���p��g7��j��/,�i��0H����ǀ��	��D0c���i2J���f�q4�'�/�Kc>�7��f�JS�lDՍPsU8GЖ!��髮��q�^B@ ,�p����O|�΂�5!x����c(�3�p�IB�.�c�2�����B�I�P�Vu���#sC�����%7Ex"Bc��#
�5����F�t����sD�{, �� �08�U�v�D�t��*�]�G���މ{��ȹDכ'�g	g�VX��.j2��6q�==��3���Ң����7�j�Q�x�3�6F��p��M���9
Ï��f����
����g7L�+��լ�z�_� �v[��67y�02b>�3#�k�G�NuN
���^���4-�H*�q�l�.�q
/5J�� �g�"�n3'-P��.���Ǿi�e��+@{�5<:��ϻ?O�i4��s!�_\1�p���� >���Z��3�e9���mv���|�x�:������{L{vc��2���Mx�z^��0�%7I!	��� Б�6XH�W�=�sm�p.�^�Jj*�?���I�	oZ�[�#�b�c|��͆$ŐW�m,5b�#���/8�&�S*�G�:Ų��=G�l�_��צ�'D4Ci�¾W���FŨ;���7�JE�}��^��-��0 S���L7�B�Q��6�P&��u2g(��RL^&�'5G��r̓���[�f���L��@Ք�TA�"���ey��\^s��Y=���&��7��sX�d%Ϥ#���d�qΞ�S�F�I��$�.�!y߰�S{!�ը{���+]]��R���L���U��笻^g��j.%9H
��f�E!��Ef�9�?98�zJcAU.��Q����]6��P�zmfϹ�p��� �N��M"Y��P�&��g�7g��q�\gѴ|ϥ�X��x\n���{��)�#B�:O�����:.ܜ$�Ru<>2���g�t-)F>�0��W�x�)��r[�[zd�t�"G1�U�u!��a�؇a��F��D\�Xs<H���`�0f�UL{�uaNf+B�8畣�M�n��N�iʏ��V��*�b��t�wѝM��8�m������K�P҇$#�JI�h�9�!G�	ozϙU�+���:);_:��C���R��%|�k=�^���T��=���uP$�"��!�Cf쀵�NYR����E�i鵅�^��KF&����L�t[��s���n��5*���-s�aS��;]Pns�j���)�$|�^B�r�aO�����'XpG�g5� *z���{�lm��IE�β� � �e:����R2�:ɵu.���z.VD&X��5�&�'�v���GUj�=��hrHk	{<�Wk�i��n^�Qo�4ʢj�q!�M�CNZ��Ir%�f.��I���M��>��p����h �n�
@-׻��0�#{�.4";�N�oI	�x�D�M �֬���1q�""���QvGͽ��l�)����"H.�2�4dL�$��r@�ט�[��0!;���R�o��T����#���2���C3`i")S�i���)��M�t��u״�:����sű�5�Nw��~Y�e"�k��s<qSϠ <+�i&��穩C��y�������۰�:; �IngT�3����=���f]%r�G_c^S�x��47��*�����,CBB��r��=sM.�����(�.��Y�tfdE��6�Ԕ���$�Y�^�jf��M)�
g�.�oM� �� ��2w���E:�Ng<7��2�\���	����!�^
�!^��>�4��dVߝڀg�Xv�G6#��lLcDS�!���Mْ1+f�>1<3D�S��Ĭ������r��*�̖9{M�mU���@���p�Fs��#�jK�n�@�����~�dU����=C�EaX����j��+�h�6��eS7b�����N&7��VPPʑ�C�̒�q�4Rĕ���}�r��\X��ISƱce����*���2�z�9/�6<��Cv�?�l�g��F'��>�s
��$�G6���#�g@S!rŃS��Ռu��V^�`2]�̛�O�z'g���Q�l�.<����KN�0��"C���^��9Fn2��{^�$g��ba*�>q��J�Q�g~�n�/ZC���$W�΍�C�GwT5�N=[*����ts͸)�T:㧤e��k�*MKw֏l fDBv$��~-�[<�2��%���������C;�k�i����`g^�ٍ����p���^������n�*�#�{a�5)LD�� ��0"�̈봰H��<�=/�΂�$�aE���q�e��Ȍԝ��ȩҶ���=Kk
�tHn�$�  ��v�\wOz�o�d�����>Eo���X�d X��r���r�m�y��>F��g�ts��<8IdP���۵�^�-<��	�����٨���B���Y8"ȸ�ŉxo@��Q1�M��XgR��}�����$C���:^"?���gsI؞/{?ޤv��3|�˜�[,�B/���M" �t���\��>��T��Ft����\E��M���~t�ML���7lf�tt�y�8�7�m!u˦��x�S���\5fi.��1�{HGf4�0�]Y	�cz	��n��9���.�Hɶ��7�@PW5�u��,m����VC�y��C�4�����HGd��>��[o�^���ﲍ��,�w��^�|��hG�1P�g2^M��Fڷ�J_��_��ݹ�q��gv�u��-`�ݎW�"��`�5c���ލ�o����`��)wi��<�t[���Kw�������������/~m�T3�k=s֥��͂&r&���<c�;߾՘���!egdٰ�ƖI���r�GUӕ�������r��D�2i &g�i?t���3�MXw�q[��WK����gբ��ah܃W�릛o�݅٨��B�*W�-9h���D7�l��6ގG������ʴ����}�f/���V΀�ٴ��g�
�1�Y(r'�J� ��fW�ą%C��n$�C�	9��7�!{w򵔷�#���i����XA�N,�m$w�͔>�ZβK�o��7�?�#��B���'�Kr��S�1���Q�ěUL��l�
Q򇘵� ��$][m���ǅ���ŏ ����r�ވӀb89�=��m'X��7��8�}��Й���O��~�L�W�{熬�e�z8ruvu�PZ\�xA����� ��>�ZԒ@ƌ�{�e���}���l﷍��[nI��r[�� �9�P�N�A�����%�O}�=�>���h.�C�����Pbp����v[q�{�M\{�A���#/0��b�������?8:��uS@��e1[�5A)OB�;��d��羐r����jb2�%�=�Ո}#E��[�F�~:D��M&W�9S��Yh@���w�|��/ _�2@q}�o6{��>�;���Ye۶�Ё���jj�i�K�n��{䐔�FԬ�X����~��x4I��X�!�N�\k�Z0��=':�):b
��4j"8����S��^��ь��{1�WJ�!67Ɯ1�Gژk��K/;Xxo�D0�^�4VQ�;jZ�$w�岀S�sa�!`�c�SjL=>?���z�hS����rn��x8A�ڜ�&9�id:j%M�a�;H����ZK��VL|�uK[���?�O��G���x�[p7�GM���a�p����Mf��z����7V��q5�~{#��z��Ta��\��0�I!_ل�\���jԉ>��oz��٫aj�7n|�e��a��ٳk�Xp)��3ہ�����/ki�ӧ��X��ςU�@pv����LaD���h�Կ������Y��r���5N=�ǽp����QB�"F�Q�{��*���%�b��5?�X��GS��Gp���'�0��������S鞋w���n��l<R`���Ю�|,�,���@�Ld����n���s���]��Un�w{����Z����XSfԜ{��G��4��(����^���Rs������h�ߏ��9 �@�q* �l��XI�A3��b�0#2�v/��1d��w:!�9�ܖ�N���o���jb�Vj�!� �~�匓ж	=���ϑ�2���8���{G����1�9Nd."��w���8��j�ۼ��s,sq,�u�A�I���h�TY\�@Q8 Sf�F�L����`rصK���6��T���U\x���G�>ua�p1�!J�^�7-ƳՐ���+��x���H�=/��h�?@i3�c1�̘��N���@|+A���JA�vm5�5/a8���hю��=H���1Y9��J���#�K�e*���Y��t�h[f�֖)�ũg�ոWl�
~��s,6�;��a J�8�iB�_�x�hr�iYu��;N�p9����X�D۩�՘r��9��\�����^[�c Ȫ'#�nd�1J�CɄ�* �9r�+�͜S��G�r�a߫�x��	�ˍR�Dݔs/s<�іMц�Ր݇�(%P��TH��yl��؝�8&}��'B�[s�Bu2��p����6��.&+��-bHk�DA\����?"w��[�s�#5��L���#���b{��%_�t���qH��a7V#Ou I@��,�*�VC�+7�\}�Y"� ?��0�}���ĉ>��}��sr2��h]��:����k`���53d���8� �*��QR��:7"u�Ȉ	�Ĕ�b�\O����֖ �+=Uc�
h�#s� .%*/��R�LD^��ƹ)�@P[��XR����%k0a��8�{3q���S\��=q�m�':��$p:��cqXI;;U�hL�s��#��4 F5���0���:�I���d�M���#hSϜN:&����$�P5��Ԙ�����ܔ�Ʃ�	�`�����M��L��27(^s�5^(l�$M��q
 �&P6���ƞ
FTV�TS�8U=����z�k_�R��`��_��t����!�>��O�}�C.T��q*�t�c�j�=����od���Þ<�3?n���xQ"�e/{�W;c��Έ���/y�Ko�7g��Q  �B�/������Ee*�v�, ��(�IsO���/SEÈi�q��#�aI���^L��q�k�����E��7��b�X$�@8&PPY�E?�'=�I��Y���4I<�K�xz�=�)OI��|��ԧ���˿�I���y�s�?���(����ʝg�?��������I�u��W��������I�f����1\MQ|����E^C�أ��1������{ ��C.U�2��DK%lm�0ܡ�XJӛ��*��6��=��t�嗻$�,@�_7�D ����(ō�l���`�0�TJ����C����5,�g�a�L�����O'Oi�qB\ęqf<�" b 2&��U�J?��?�c�d ��i��	�!���gz�`uw��{���2Eo�c�; ��=�y��7���M�Ɯ�p=�6�d�N��Ki�6r�
�4h�y������IP�O~�4I#$��!�)� 3�8^��:8c'�6��1 �4}�+^�7�g~�~�M0pu�PP����A~$�93Ό3����){F��`��׿�����>;;�tXva��x!}��캊C��<���y���M|Qh���&�NEQ����sc��pq�wp�FnRࢸH
�sQ2l���xj-��M�LmF���,���V:k��1; �L2��x�~�����Z�r
%�q];3ΌG�P�����}�5�y�)Z1L�����܄�S?�S���!E:�)8��� ,��"*"Q��`�;ǀ$�XD�:��&d�����jR���b� ���L>mo��I� �0]�$�I���x!9��w�N�����i����X�Vc����[aqL.��n�gƙqf<r��%�e	^��pѾ�����zM]�g��$h��`V��g��2-D;/�rNp �[<�A$C�6���	�I]vJc����;��p�!@G�MIރ�"q���'�C *�	R�/�5;1��b���Yc�A�5����s1�?�3?�Cy@�p�p���g�?�X��1[b����L� ����ڵ�?��\	�k2=/yP��l�;�+0G�#ӄZ����t�UQ�+־�&|ʣ#�bSQ#<��[��x�ށ�2�L�)�q�|N���XP�C�d 1�)�c�m�&��_��_w�x��L�G�>��Ϲq�@��Q���V�*p�錝��83�e�h���a����T �������{y���/Т�  ���A�wԵG�l;H��bBS�#�$��WҴ����pܩ��Y�+:N߉��瞻��7����2R���
n�5���q��7ߗTSz"����;���xA�U�.�G)6�����ԣ�<?���)�i�S7�+UD0w������^o�Xo��\������vѣS�-�H}����K�������F_)X@��W���t�7LqQ�E�ٖE ��M�7'ƫ�f�2�x�F���ٻ�'��EK9�q���1�=N���M������~ћ�E��g���ȉ�Y��thW*��A�}��w)DV�7��Mnfrc�e�Ek��g�ԤF�^�;,��i���k��m~;7y̽��鎿_W['S��c>3N瘷�Ol=�e���"K�c�����.7E��oH/zы�������o�qjj�o� ���
]��H�x�j�����6��P��贿�o
�We�Z��Z.�~�u8��skn=T�Ͽ�)-W\�nP��$V�<C��&A��߀,L��~���CJx
���u�sI��3�ڞ��8��3�f#��4�̩�*��i`��������W�ES�*��)�K#�3��8]c��?�<�Io^�d��u��-N���L�����b��a�Ҷcy�؊(�=��4�A��{D"����r�m���-A�c��锹=w���`��x����=�t1\�b�f�����\��4�T�"1d�����=�d��yX8������Όy8��:����y�{�u[�W��zsQ�<�Pc� l�R4t'):�ku�83ΌS?�懶Y�h�y�8��&<�'��w�=&HH�˷���C/x���2?���W����>�'"	��>�a%��=*��\:S>�U�F�_������M)D�-���\��rp2�K5�Q�1s'���*{EG���������&�8��b�����.[N�Zʠ�j��g�
UΤe�\C��(+��f���j��jG��3�Q��B�c^g�����>�>�6T��?��� F�c�P�� :
��_��+���%��MR��b�ص�+p@X�h%��!�Z��g��oxksĠղ]��<eY�]g�L��AZ_��[5�i�t��p�ܐ��	l�HX.�p�v�vM6c�$��%6�	X�R�e� ~,C�Y��1mne2����g�6oB�wJ�0p��:�������b��c>3N߈���f�Gc�G�����T�:`�����w;�3���%4b0 ����5`�� ��Z��`�2/0�a��e9�%�q8.x�5t�3֝����~ԅ^W�l�U+sm`l0O�}uX��^��Û X_Ib�
��
�}�P$1w�,��!;���m�]~�b�T�GP-�m��)��+J�#�i#cq��"K�c����ek
�9�Òs7\�Mg��,���3��3�4��bs�&z4s��z@�}1ѱu*2WE�0;���o87��%��5@�$0�2X~���*���1Ҧ{�]������5d�I�i�\vG��	
�$1��(���?HW����(�zh�n*'^ �j����3��"@��"�H��*!S7H�5�Zbk@� l*+���/v�ü<�R%�;�1uʀ	* �1l&a�*���
o/�tS�-���t3�ٙ��1m�әqf��!�Nb�G�cq�EU^�SU>��p���'{���wyf�.˱j�@Kam�0��`�I�>Eq� ��5���\��s�po��焩�Qi	�rFk`C���|��_N?��t��d�ét��3��S 5�����_���}2e_Aa��+8�G>��h�X 7�:��ɐab��'��>�չ��&[f�t8�,�ic�PZ^��h������x#M0����,E�Y�1����pL��N�tf=��������P�6������S9A��=����L���L�G֦��0�ΜxM��暡g��Bճ[���u*���%�ߏ�i9�֔3&��S�RϺ(6T�QlI����[�T����Q���\߉eY�7y���b�����o�yf�V�<[�}F߈�I���h>�-.��0�;Q]��6�G��BW�����ǵ4o}i�D���*���x���Ҍ��Km�M���	u�͂1� �	+�-�װMS2�h�M�>���2u�NVۛd�`����>������!҉UGX7�E�bPzng���~��n<���zP*���u&���"Rڳ��c�����`�t�[V�k���0{�ũ�����d���R��U����Pw=�Mҳ���	���`9��Ua�f�<|(�y��k4W��m�3��D��6��ɟSP3��kk.cXN;����q��0DE��,"���Q��q�ц(A�s��qbcƨZ�dc�dLT�E0�wb�,�������lϟ%�d��rZ�
i����k$�g?����磹��IQ����9"��ׁ����j�;�u��p���k�5'���	J� S�G���I怈����b06���ߔH�%0)��������	�;h�C��N�8j�e�=U9�����v�^z�S�꓃���r�jE�`q21 0��=��J�j)�Z�)<�X0�I��j������l�?h$�(��I����sv�z����0���4Y7 6��v�^Y��tO�p�KȞ��~z��Ҏ�.rޘ��λ�I��E1sv(�$n�MϠ%��_�U�aH����<��z��Њ��^��o�TF[[Խ�Z�uEO��'Q�n3�M�v[=k�|E�C�MM܌�P�5��ⳬS�[���j�<T�J�V��GdB����D ��� MZQC�@=G�T��U�a�1�I�K�����c$�T�ڶ����h�k�<\l�B>J�ҵpm@59�t�|����<��`Eh@U
S�	������o��?7�#!%�*�V:�q�*j�lc�䅼h�nf�D(�ݻ�A�e)y�Z`L��j ��&H\n��b�I=5ew2e�d��L����������mS�a:�3\�����0m�Hc�i�L�o�;�L��1?$n����z]S��:�ԫ�>�*�Yl��`p=<lm渨�����.��{b~����o/J�#1a͹j��D�>��f��jck��Y�X�|Qx�"Lb�z�\" k=H��њP�n	3�(x,�{�f���	7�Pe�X�@�)Е��c��L	F��ya��9��F�>/� �}VM4|F�s]7�M;ZC�5�sH�E!x2� [�Yb�c߸H�tj��� �-�^aN�_�������7��y�w�|E�TSq��xtsD�)�d�OV��^���Ƃ*�M�t��܄<7s0^-ˈ�$Q�e0	T�GRi��q�yO���g4.�gK��b4d��c2flG6�P0 .�1f�I��ii��a|Ua��h@�En���Y/���{�nV^�s��$�z���,7f������ʓ��`>����N�P��h��L `��uIeBj��GtrD6�g��1�R#�H�&�X5jM�髽�/�f��\Q;�J�om.]s�=��hֶ�1�:�3����Q����ɼ!����(��֠��.^׫=5�v�A\x"㎎>�qt �[_�2��������K�A�F��/ӵ�=�t :�	�C#�<�u�s��^�k��jFDavl�i�>�z�2ؕȎ�v3��Q7��Ҡ���=(?�
*��D��ő��a��E�h3YZ�L���5ǖ=O\�Q��h#/��*��Be�W�lA�vX�^����~�<�*���ʩ�%��Pc-��0e�,<dc��R[���b޸g1Xݣ�����Rs��m����ܺOƑؖ����D{�
�G0��#��Jz֑-���)@����5�_	(��~�di[0�L#�D�b�1����������"���~#co3F���Z,�=�q^%����H�p$տ�^۔��q�g�&2Ui���ccp�cQ9Q�eQ��פg�\D|���N W@�-�����x��=#	�h�kk���p��V��B7,<�A����ͤ?L�����T�B):,Z���iqkB��8��c�6H���&XFcy9gj�_~�1��������
�#T��Sy���T�̀Aẜ4N��ɣ& ��Ttlsv���y�����]6�v�T/چ���0�5�V���5�,@�T��E+�)՜��(�E��&&�+۶Y4*m��Y��)���H�"�^ڂ�k�����F�?F�(
�m�՚��x���<en�YM�X�����^P	 1j�p�f���5q�<j\�b��]ku=Q(�AYj{M귀���6ؗ1��D�� k�k�ه��_p��ڋ���Ks�&��7�)��s��k���#�(��υ=*&K��f��ؽ��Ә@;lʙ�%�WLL�Ɇ���ʪ���V�d��MK����~�Y2����<�ԫ|;e��~�I �669���ML0�k�m \t��r��oRx�v~�H�$J���.a�ndw�m����[�M���juu�Ȝ��	���?7=���{|��Ճ�7�;���cr^g_��������~&��{ -�=%c2��l��;�W�������=�g"n�8X�lr���[F�%������g?�m�b�Qk��]���Cj��72�ig�V%�Mt�I�s<� q�j�6B��vZ�A�^���CmU��(��@0���2ma�� ��ԧ|>�k��>6!ҷ�76�z�����tŕO�s��.�����'n�tZ�=�|b� 	��]=��\͢\d���(������F�C��랢�"ڡ�}��s\=��@����A�	��)tO�c��?�HĮ8�G[3�aװ �ș�b6k!4�����4��u��ۖ����I������P��a�9�f���΄�Xۢȅv�����\����l��.80�;������NDWTv9��1ݾ���$8��a��G}5�cM܎'n�÷[�O�:A�c�#ۈk�i�9{Үm;�D޾���Y��i8)����7��ඥt�TK��L�F��P��?�d;��h5�}�Y�
WRJ��mz���"� O�Es�g)W}c���L/����F5��c#��~��
9��%��h�I��1�F�$��E���(� ��Ħ�&�/ ����v��J`�	׳��3�]�3'%�������{}c--��H;�9�C&K"q��c��ʆ��8d�dt�������	���}��~>Cy[�k.�i�N���=�ԥ=�~�N-�����5F�������8M5}Đh�o�i��{m�,~�mW�Y2~&���L<'2�nY�ug�Ņ�-�������w��BtDck�EWgV�����N���q��#n�u$����M�	�i�$8֘�0`g�|	'�Ԧ�T#�dݴ<�s&�D�ƺo�����IAH�r7�5�5�6�B�Ū݇��n�>V���bw�����L���Hy]���T#��V"V�!}V&(9��I�#�p���}@�]�Ҫ��F�/;v:�� SL����C�E�C�I��X}&F=�L�:Eژ��ӛ���+�w�kB���Ę2�Au�ر�E\;8F6*| <�:'v*�j���
5�l�4�ߢ���#"���8>/=1���F�����8���'q���V?z��a�K���6n�ܱ-Б-�5c�K�m����ma��1������6����պo��b�|/D���ӛ�dUiۤ�����*6�1�8���Y�x�+��U�y�LK�rw���{{Z@�3���k�bv���7ꑳ�����%cT�9�Y�Q8V�AZ��1����<�����z���.b1Z��K�f�A�ًRP����� �z:F����,#������D�Y@ -u[ -�G�G��f��0&	�s�Ĥ)�����N~��][���!�nH0a:H��0�~h��|���&�T-6�1p�%�r������N�+����T��ZN���%��69�"����qޣ3.fk�7���':�i�� �g��9r�y�}�d��|�ќ?�D�#yH%��$��g,uyq�H0�2���Tum�ox,������=.�66UՊ΂�������0S ;�vw�V�c�À�t�}nBź�)�~(���zm�~�ϧÇ�i>���n�X��?�=�DK��=����D�`����n�O���O�s�O��S�� ��qd�n�8娐�]aal6JR�C����8�8.��WLWj����qS<qt.iHȡ%{���� 5������j(�����)�#��R��_w5i@�l�W^'���L޽�,��se��;�Pdi����l�84J��ݟ�n�u���߀�Wd��J���&�����aƵ��IZ�,����lJ��M�8��h���*��ˁm��j�J�m������T�~�wƹzjL� ��v��0}�;?Hw--xDDQ�p���jºJR	�m�.���V��`ˁ1սE�ƌʅ����!��� P��Z�W�M|�}}uZ��ҶA?�����;�L�{J��ô`l��R��ᎪQZ��9�7�\YN��]��z�Kd�7��q�s���n���-A�����t���0!1FEN��V��bYb�����̥���f|�8�,%��?�߀	M_N'S�;��~�@�L���p1@���y1��1�k�u�E֗��7�2���ם���\7L�*�;4�nB{����u���0�� ����`j�"'��lmM���v7���:5����nn��A<2X���p���)2�4'��ؠ�bw�O�7��"���Nt|O�����y���cl	���W'ɀ�$UN�}�xg�{,�I����e{؛����e[#��5�T/o�i���~���mE �nM�0��RNY.l3q�ޟj`�ks6��U�R�D��y����ɚ������;��=Ʋ���� X�f�kc��&����s�6��)��Z��_�q洸�O��Y��tNZ�C�QvTm>1���L4��]�,�c!1W�d����G �8��4�}�h#Î��y�M��L�Tbև°\(%�O9O�f(?W�U	&�$0������y2���a�V�[���iLd�{���y"�a��>����l>��Qu�rB�k)fi�1r��]��m����_��1Z���d맿[�-�o�	��G��9���6o���u��9��u���Qi��6�:�%�p���X��X	��G��l�:)���56��iNm̅�aSpP��&Y�����W��:�me�iTO�O���Dc`�s&��4ZM]��^�M8��,����#���B�Ŕ�U�����h���+;R����b�	�S<����S,*߶�	�b2Cj|���"C�"@�衎!Q����~R���c�� Gl;�,#�ơ�-%X̛��� u�a���A�P≢�Wl�1m��Fk8�kꘖR�h�l�u?��Ꙫ��0���$�'o����sM�T�"�3/K�w-��&�l��Hc��N�<dGG��(���4�c�fz}�#�DƑ�b4{Ź�@|*�tsD��^0�����D�m���U<�ei���:�N7~jT��&�v�l��V�G@d�!v7���V��no�`���մ9h�#�Rj��:+���x��r�������L�u�����H�_��fd��c�w��:����9�W�"��F��v����x���!�X	,���G��s�Q��\����$�(,�������	��E#^[,����y�n�+���{�N�q���	]н0Ѧ���'@����5@�K���Ԍ�򣻝�y6��Ud'���L�4�_�I�6�T�H�GS��ޓ��dAj����Ɍy ���^Lw�Sk�E��u���(-���PG_\�c@5N�y��T�"!�^�R��{9P\27�� �%���Oa@��dRT�T��Yu�Qy|-5T����^/�ncuc����:�~ʙd�T9!y��o 	��M�J��P�G�p�I��י����kg��l;6Y�Y�hc�� 7jc6�@b��N��"��=�(���,3II�:!a�d�6L�Ʃ�6]1�*͗�S@!0�RI	�lJa�C��6#��x���ڶ�vWLmg�"/2(*�`�fo�λ.]s.�+1�NS�I6��	���2,I�1�h?h/�Fɸ���z�a53KW�
w��S ڪ��w6��Dj��Cg�$�ǹ�(N�ͯ↹�X��H ȏb��~�����v��u]J��?�*mb�*&{t��^�$p�VY�`��Z�D�����b������<1��%&��6h�+��v�?-x�*�$�� $��U�G6&�������ƍէbH���3�4?LJ,����nm��q#����z�<���
�����&B"'��D��F-7H��\e
���2[�,4����&��M�I���d�8R������h��_m�ڦ���^6,˄@�͗,�n'�D�*�=��k�����{�`�f�I����7Y�o3�x�v�!&s|G
S��<���B,�?��3d��gu�z�h#�_���:�NZ�׹w���JA@W�����>K�M�%��
LU�ak#[� .����� ��w&^d���=:n#~8FDD�SL�j�蠋�(͙b�e_>��5���I [6��p,��H�3l�d`r="s�Y*dN L�4��Q5�P� �؄��I�	��� ��-�6L:�L�w|'���7\�"N��p4L+���F���~�9'@��.ʄ�D1e�@�M�K��X4nr-T�`_�җza ���}��.�X\1uV���e��JX����[4	ިsҘt<>���Ÿ��Q�:�d
�\ �.TfpV�g�b�d4���"�o��!���Wm�x�0Pi�k�Gg��c�7�=\{z�ؘ��y�s�u���=�s/< �c����a�3�换�:HsUx	?%^H�V�39͢SL�}�*Tx��N��<����Jh��s����ў}$[�Q�E��A����V�v�C!:y�J�W(B!���Nm@a��%���4�Rf�n�*�Z)��i4��J��:9i���������q�ur4=;�A,+���B̈�&#���ﴝ[�ʄe��is��U�?�J�߰c�븬IՕQE?��MI�`*�I �P��1D��K/ubI�a�tyw��D��l�3��n�U���$g��];��Wz�>҃I��Z찡,)����{ 'L��Efx��� .��2/MX�z�!�uW�ut8Z�{Ǟ����]w���;��{�ңO�(T�~;�,�n�u�����Jc��Ļ9���F�cˈŗ2�N�5OS&��6�2��#�i�c�� <�@���vO&��?��k�d���Yp��}əyUO�j�I��[͊��ȅy��h�P���Z��<g͑���y�g�bF���h�����o����J�D/��H)�C��h���Ѱ�.l�wsrVd�J�&�nl��=ת��Z�s�x�Ɠ��̩����9/SN��Uk"th{�u`*�L�2���O�y���[a͋��U�pL̐����Dm�\1��_��w�t���������Z_҆b�r��A�=+��Z�� ^1t�h�`@͹�.�@ c�f�TS�r�0�tSD��9>�E>���M�|�3��=P_m�5Z�|I��7`̀0�O�yL1)�T�0��"���?�gΆaҔ���=��H=y��$i��E����4�>9��(��=lz�!��*wZ��o�!��p=3٢�馆9:[�x�*兺�i�ôL�1��U5%�yO宭~a�gp��r1�ln�Vؽa��k���4*5�M6�Ϯ#^��mA-nsU������_��X ������<�)Ô]8�T#@�TN�p1�-�-^S}	=�y#:��(�I��n��U$f�Ţ3�OF4U�m����ǐ�-�*�2w4n
[���A���u��l�{v$x����Mc������8�Ԧ(%R�b�k�-ΐ�F���A>��Κ���[�>'��aqi0��5�}�vHEgf4G��(��C�x�|T�b�v����e���$�b��4� �8h֊?���PR�PÆa�M�UeF�b�0:α5�t��b���Ƕ���~���'x㼃��E�쓣�ǐ4�i����dw�_��88�q��ȯMHf�O��O��O{K$���o}�mx&�caC>�M��lBm��ZJÜ=t�9��A��p}H)�4 �L���Z��rvR�+��xQϣ&(�C���c4��{�v���fZ����V�@?,�P6�ҍq���߇+[���C�l�~.�B��}u��3���������>�q��w ٰ��qb�E�K��\�8T�W�P�{bќ�؊�@o+O�l�1ck�sN��b�v14��u v�k�|���Mm �JP����t�N�mJ�FR2�χ�r��gK�� ����p�M�����][O%�b>�u_�y��.��i�y��z�F_4)�N*&����8}�C�|h��ƽ�&4X%��)�1��Nt�� b4�|��^�����p�~t\WK#=?٤�7&X0X��7qM�u�>��P��z���1Os��ԛ#tA�ⰝB͑(\<,��y�*Oi�Ǎ�k�j`�H!l��^{�Ԇ, M2��t�M�]�~x�9������l;}�:JٹAhW�υػ�4�:����g>5��{G�G�Ɣ���{�d�pZ�i���M@�Q{Y�\�,|�(h�-��>s�b`@oB��!7�`�@-�i��ձ�w��;M�[�2�����0}�4�Ʈ��Թ��&�'`�)�h�ąцmdJ�7�i�;�e�.�5=�6�!j��LE��:�1BE�]�o/�dX<�;�V�X��~���u-mm��[�&p�K폩�*D�cE�m��+�q����?��7��j���E�:��8�4�ά��-�e�6F�`~�F��ɨ㭳&�OxM�Í�!��J�]T�L}e'������\rI��)4�̚��[Qsh�6�����g�"Lt�A�mW�;���zo��]s��*�$����7�ɳQv&Z4ׇ)��DS���ֱ�U)�s�q�O%���\7?u}�R�� <��~2�Z���:�m�V�7~��n�X0�{eI��#�M�D %)�lXn
�D-X&]]
����w�ˁV=Q#x0������XY�9��`?���A�Bw2ؠz\|�%�=g�Vb`���8�(�R�6�Z�,�(|�0?�[��f���+uw��g_l����R���{�t]=����h���͹�ۻq��c9u�=?-����Ѐ����f�O�A�T6��}C��{��k!=ɀڱ֣*RZڶ-]x��q�\<5GD�AJ���j�ʆ�EK�L,p��DV�A,3o��*'�5�x���4�bW}Ւ����2���lLE���)�)�9�Z[јp:M�a^����0�8x8��ƺn�ޝvM��R�J��봲dp��!���j��!�y�!��`�~O|�h9USv�����bP�<7��s[�;}/o߾��J��P��CM �φ=�e���w<CRp���ɚ� �u�z�f�Bz<D: ���������V�4�V��4�;�U�
J�z.:c7v��b+u����\�zt���+��Jm@= �/�ls���NX�ֆgp\�6R�̓��IT,#���>,���<�y@[�^�p��|�/-m706)l��ǾKҒTɲv@��L�(;�_�C<�t[&�!5aOEV7�\%�fٔ�d3Un��̮I��,L��t�������Ҏ��Vnj ���������Â�ۢ<�p�2F�X�=����x�׆�g_�3�k�N[-�_Ӊ/�_a��h<��zի������b��y	��M����Ǝ���Ƹ���Pg-q<�1�VD��Ą�cFN�R���ņqİ�c#�����H@�{�1���Z��G>��gs}#�B�S���0��t�B����4�)��ͼ�YX`���d��VǦA��)�dߙ�����wsY�����&��h�Mh�^g*���2�u��D��J��##b4J�d���W�WݎKQ|��F�_��z/��)Z6m������1fz�&�+�w;R���=�*�T���(�6����i �Q�����������t"7�»g�]�*[1�JЈ�|���&��;y��E�Z4f����/��/��U�w��Ƅ�������Ռ��,:�x��Ԅ����,7�gΑt���"�D�v�q�^�d�n"�5^��].�=u�Q�%z�SVY�,M&j^�E� ]4@g�k��t���Rw����NZ$��>O�:�l#;����a��`�k%{��D����dV�K�7�ܤeD#�Q�����%&u;Y!F>�ϭ��ܡ�c$�W��@�k�@�=8f��d���	��O#�@��Z��f�H��/��<�ǔ�̟}so�L��\J��d�x�4�Uڜ�:�����»/ w����S�{� �N�O�7\�%��漺c	ӹ��8��8����@�<�W����^���?�A�|���p
 g)�J �u��i�J�H��	��c��M�O�9"�BMg1��`��6��K</�=n�Ȣ�jL,�E����t^}��n7��G?�̤��o�V��?�c�H&Z^q��F�͖6=���m(*�Ԩx9�l����u9�B�<C�3����^쎿�|�QAP|��i����g����,?t���qӪi�X�r��QZ�.�=,�Н��۲�86�3�̞�&4������o9K�Öp�=*\P�|�|%�E:̋z���Q���'A�.�.��-��R��[�/�4�yf�h���%tt_ڴ�L�:�K�����I�'w8I�X�g7�����L�Ns�\�C�x�.,j~ǃړ��o�Zݸ���x��,}��ż +��a�~����{i�<G�V�g�o���-F��GX���7�A�LII�-;'t�Gi�9�	kZq�ZZ,9 ��Yeɟ���1�ͅS�6Bm\&P^c��̚�����o~�g�D'���
��^���ڧ,A�h�K]z��=�n�s�$%�Λ(;U&I��p��w�kE�Ջ��zS��'^���v!��n���t�Ъ�g��Toq�$�&�y��=���-��>��1Eԓ���H���~�k���yc��s��`S���v��
��9ڀ�F�^�"�g9/�}���ϫ�ql
ӈ�&��)}?ޫ�RM;?�Fvg�����L$��g�M�lM�����{W���4(�Q�m���A�Q&lQi���%��}ዼ�e� �o�,�ʠ"����4qq��1&Ј!�Mws����C��uߟ]ߺήڻ�34���tU�}���~��o�L�͂�e���%�}w�Y�l���#�_�ş�m=?� ����;�JzH:nS^�G��f��m���꺧e��X@��>T�	��I}j=��'�i�K� F�*�[K�1.�H�"`�#�=�;-��Ս�S� �7/��J9�tL�]�=���:���j��h���§�?��W}�W����� �l���=Z�a-�*b�����P��А�I9o�sp�3$C���%v�9
6j���YHK�cx�+W�){�=��ǚw���}�io�:d��VN1a�ӈ?����5f1-J� ��u}�����8�1�ڎ\�1tP�k���ph�f���h߻`r< ����1����ZF�����@�7�ɧ���y��9�G�gl-{+4q��x�w���K�?�5l#)	��d���7�Q_����m~�����?�áF� �����-�j�Z�	�3��w�l
�E1�Fx~�NjEc*�S-�������,�������(�n�A�,�n�<�ƪC������,�^���?��r�1�1�a���@��k0�<c<�}A0�LdDk"c��D�0��5�yM�,Lt�-��|�:9��ps���
/ԍ{���%�s\ �L���߫s1�k�ZM��v�=���:4�|��=~m�	>�ȣ}Vނ��*am�o�$(����� ]��DR@ee�עд��L���M��s->��S��a�Vh߸�bΥ�+�@�i�V�㈾w��L&�X��|&�'�-:����8z�� k�ױ��(���h�=Jm�[�='������c��1]ڥ�}%������������gǏ�e���0�X�H��������{��җ�z׻�W��U��^����BQ��:��g:o���q�d$�ϩf�!��x.��|��h<����Ɂ�s� �O&7�a�j���y��"i�9}�>�:4a&:x��v�=��=%���:xC��?���q�1ji��'e<�$��j���>��p��Ӳ�r;l�9��F�h?�X�z��Ds�-?WP���1Y��QےSЄ�x�䕽�g���|ڧ/O�>;oww�L�@Ts��#uw<�Q8�_�K�z�C���!L���.��km���\�7kx$Ր���i���uԴV�D25�!�$�M(��Arۚ�j��&9�右ԧ��&��Y=����ܝ%�G�8Q4Kj��К�h�Mb	UcK���I��Ej�q���ӂ�j�7^?S���}
D� �l�%�@t�l��؏�N;���4��x��;�A��a�CA
l:�Zt 7@ȿ����1�wc���xy��έ�,+?QeNy:W�T��A����tB~��4#t��9�����P L:~��++�k�d��%l��󶯐F=��bҁl7q;�q�N��ϊ�eT��+�Ep��{�찱h{��h(�Px{�U��bqXwb~Ѓ<�=�Bq��;��Z��p�l�V��ս�����xf�+����o�����u2�E�䲬e򢂗א����w�m�L��woHmE���JE$�;񼎜5���j��<���g֒�s���¡W^��J��h�v�ԕ�;�I*�}��M�����1�<w69���4ۏ����;/}�{1�q�!�`�h/�%�W��v��3t��*<�5nҿ`�t�%T	 0A,���J��i��dMx��Tc;+� �^F�X|�+^Z �����b��H��9��z�iDB=hh�uZ�	!��M�T8a7_t���/���MozS�����z����LQ��jٞ�w^=婟��M�>O~��.���uZ�b�M�	�ޏ�&͕�I�����.�&<޽��~0j�ߠ@_�}���{�Gy��j�m8]�:���e �յ� �~}/�����ﷇ%���b*�e*m��LV�{�}�V�Ϭe�����;�ɽ�N����'}��<n������9�M�-"���֠u/4�3�o����MGM}LD�g�g���~پe�|���򓰧r���w�^	��G.<�>f��$�>j�_��=Kz/�˒����0w�F }��8yv��P�x���ȏ�HyBW��ۿ�` �,kS���Ll8�+�`]�h�j����x�Mr��K1}����i�l��F�0Ԉ��-@�p�7m>��Z��08՜h :�����9�A�\(4��_X.╯|e�v��_����Mf��|�ה8a�w�աL�t�!�Xj�P���o/IT�"�c���"���m����H����E��P���nF��{:��4�+�t��Wڍ{Q�`^���)4���1ͥ���̛e�qn��/[��2Z�N�^��j_d/~��/9m�� HH�0�8��YZ��I�i�b�2��h!3�.�k���~˷|KI�b�������_����q���Z�8H0#����#iK5^1�s��(�;ڊks'�:���S1h/<:�4��0�c6�/� �0�y_�З �f��	W���X���r�(/��hDk ���[�Z8 �6�5X�h ��6���P4�-����/�i�&&G8/N%TƗ6���(lo�y��h;�Q��+���ލY��P�	J�ٞ;�5�5����.٨�[����KS��C�:�/��m~����e;�Ns�C�oM#��VǶ��9�~��eJM�b;-@���D�Mjg���?�Lk��U����#:ɚ�ʦt�?������</Z1|1QS�IF�Xl�yL�.�n�������n�c���h���~���Hџ�n'eXSDK��~o�-��xz�9�yn����U@5�Qn�tP�����AepM�BY�$�O�tb%b�"&��m(�#@�Fռ���a֧E\�(�X�Nh�=G�$��L�}�Jj�Bo�8�+�X�o/i�MS2�F@_�z_�1&K��q��@g5,%��k��6j���tr&��[ṿ��9���~n�:�l���f���f��c���|�*R�s���T�N��:�Rt�3��"qȓ���F�3?�3P���"w�A��:d���2��5f�N��҅k��v"<ҡ�mw��s�E���������~��>�O%��s��9�QXa0G [�4n�B^����ĺA��q6�f�GkF[��a��m���Ȟ�zm���J�-��1��b����%;���(�4����h�.�6�������<���L����G�5ړ&�0Q۾OF��IC�)��t�3�U[�di� �����'�(J���SN��c\>�
Se�c3U=��{�iE��v)/���X�k��et�d�&< #��%��ǝI������'A��zqqʸ��X|뫨����v����%�΃a
�����8P��z��Zx`V!~Ҙ��h��2��f<� �f�3L��c���Vɧ���������a:��߸D?L�^�-�/��{p�H�f<�U���z�Rf���Jv�25rѧ1�b'[)������Ak�{�5C�E/�C�r���]0�H)�v Ϊ���d6��A�+�*C���=L����0�Z6Q��M��K��,������OxN�b@�H�YZ��BQ���8���F�P�_��Хh�p��x$Z�֋�#JC���fm���a��br��,$�y(��)��B�~���8��|�s�j���%����3�+�n���9�`8�㏼[֝��u��M�މ
)��P����Ė�:g}�>�3���[�Þq�E30l pI�q�ŰS�
����WO϶��%p�=]X�e���	_�����r+���Y#�qյ������I**���T��SW[q�G�s�	̂ߑ���6�Ęm~�������6܏W��CJ��35�<��qԁY`ֹ�9m`Gٔo���C�?�UN����S�=�Gn�r�͵�5�>�f���2n@$�U�m�����0����
���Y�*��*H��Kj���gL�I���Jl!�����"��+�q��Җl4����Í�q6lٛ��sQ6U,!-�i�ϕKI�a)�c�5��4SգNЧ�r���;��>{Ϻ�p��!eF=���xnk�x�*ǷU��T��y�kA����P\�7>��ris�NI�	E�@;�O���	 ��9��g֥���!:��5�����3�#�d�C�ס�}`�:�Ǉ�qR+u�T���d�)rKj�5a.@g���l��$鷋�,'ʃ�ڎx����)1F?��	���5{V"ߢY2��t�O;-{�!fK(��]a�rl��#�mn�܉�o�yE����cW�����)��sM',�4ڥr��γ�x�JTt�o�(��Ӷ=ǳH�Ů�N^��]^:��c�T��������q��,0�K�?��w̝Sr�����>I��G�N<��?h�y+��ޠ�V�w+�![�崒���~�ߗ-���4��΢m6�|: �z�W�M+<����V����!u�S�~����I
�I�$��5g�4��ٖ���rF	̫�n���~�����RGc(�FU��~��wV�
M�,@|r����b#�$ d~.�m�(���滕�|��y�vS��*�=��׶�x�ss���5�+	���^u����oAz+[yb�y��e�����d�9�xf^8#�ڱ�f�me+[�����8+�x֬R7Q/R��i7�};�3k�.�q���)�-'���<qe�OhU�^�y���*���	�N���n)H1ۛ���>{��|�Q!q�f�el^Vg2hN��5Ӕ���6_�Xd�#��B��4P���m�t[9��s|���*ӯ�`�
�O9)�,���DZ�s���\r��N�:���C$�`��kȝFΛ�h�� �i��I0�9��w�sS�3� 3��td��c�M�����='\J<��O��Mg����+[���zG1���������9��[X�
jf�X@�x�6�ŧ�\�L��CLY��j9S\�	�)'i%�����}c�yN�e�b{�k�Tw��϶V�v�=�ռ2=xUM�z�;	\3�vG#Y��y���!�o��3=9ے���Z�s/::��r����ֿ1}��`�G��Ӿ�uuz�v�;Z�԰�O�[Y�F��Ew�����+��Ȁ��C�bn��dCԓ��6<�n���f�]F_�
���� |�y�8�:���R�:�cV�����LA��%�]�o�9ۮ��vzזF��*P>�O�`O3vΫIg�Zֵ3����cb�J ���Z�f蚒L:��ӁUVU�������pV���R�٨�����bSv�����G�8_W��Q`��Ǽ8`�N�!_���`�bd�d�[�˕�MZ��t�ֳ��|�C*�������x��ǣ�2)kJ�,�L9	���]{�8�D�ʸr��IB�����.I�X��8z'���ˤiR����u�[��B��Y��ZH���w05]��������(u#����N�v
��W�."�[*3ۚ����|:m�����H���~g�8ǻe��g?��e�^��GTw&
�%.)�p��=��x�41�G�����5A�/��//�Q9�FB԰���J/�&���i��d�{M7�,̀��Ȫ���4A}N~2���� �-s�%�U�A`�
��֝+�iL�֌�ɂBtn�$����Os�ӊ��|/bXn>�q�VV������g�
l�6�#���T��d&xC�]�Q��1�����e8�vvڡ:P�}4�\L�|v���^���y����BV%�C�MHV6��8jx��g�8��]3���W}U���5��k_�ڢU��~o���		`#TB�o�x�UZh=iO#5�X�l^7�s���6Wq��-w��=��K��w�d?���bCaj�J��~�p.B�c�t�*Mv��c>�Rp�0U�jk�*��Ɗ��������+|��e��?��?-@��(s�-Q��������F��=�tI�mt� ��؎x6���lY������K��-���4��<�J���'�̆}��^_Zg���AL�p}@͘	)���v�s<��NnX����ҳR�9�4�yMM��4�$�z^:��kgIĴ�r���E0�m2��ww�I�Y�d����}�Y7�Wi�g�\��������h��'4�t�%��ri�_6��P��$:��������= �`}s}�oJ��:}Ԧi.A��Jw�	�N�CǰR����̧����R�݊���N�Gx94TL^��/yg7
u ������-��_�x�7U�9���lYM#
�4$�cʥu���x��G�e�H~�����owQ�3��e��ŹG���zCG�Pw����7�U���w����y�i�o�9_;p�x�\���_�=��X��F�<Q����;w���j�75Ԛ�Y5�7q��ǿ�����:Kd�Eܟ��`Q� N4Y6����_��%�HG����Х/y�K��P����(vL>�x�q�A��<�X�+��+E�ĺ�6�:B)��s�^��3>�h�t�������_~xٱ5#��/�Ơ4 Z1+��ԅQ���c?�cE�������5�{<q,�����tXzVW˨�ض~���ge�N6�/v�M7GlY��Lg��рp���-F]�-��>�V�)\^S�zQ6���iL���x���	��l�Xn�Yvʘ \��&`s�L�Fv�6�^�ٕ��b���^�κw=�w��)�=Yx�S��;C��E
�!���G������@�����.)8:X\��?s˘�l�c��������n�)~�J.()�$�%�[K_���
YJV%��5��?�3N_��]m�F��>�s��������׽��2�%�k�7ύs�x�[�R��s"`;%���/,�g�b ���MHݐ�cxfϷP<�>�_��]��3�\��~Y��\h/l��áŲ
 �L4M*�&C9�2��5�8��b�¯Q�cJ�-G�dr}���+t�7}�7�p�n� ��|���>�w��Ґ��W���/;-�^5;��y7��zf���x/'��k�:��4�vV��Ѽ�9[܏5�3-G�_]�X���w�����~��q�i�������4%���]:&�Bq��N��?[.<�fm�N���:ۦ��6�� yw^0i�]m������,���e���a�q������������rZ: )!��DY�?���B�o��ļ���6E����j�*HI
RF%����J:�yf3}���v'�|n2̎���:Z���Ԏ�Fay=#r�C��ъѦ�+�jX���.8N��\�F���<��4�м���备?��惥G�4�<
/�>N��4.Z1�n��G�����ſ�e C�9\�E�x��ye�i�@��݃י���ʻ;�d0�H�{������®C
p��8��i�N#�ǃ���Ԇ���>���]���+�9$â�@��]>��� �N[���f��כ��N���V�!C����u�$w8N� Iڒ����zf,��Ay5n5����C���h�Z��|9�w�n��N���]��M~ү�- @�~B����]m��=5������:��J8�981g9�t�����__@���/��|M�������=yN�%�{��9p���X&�:F3��4�
$44(N:�o�UЇ�@�pV�*؁�����}ۣ�f��~gRUx���ܣ*�s�Hh��X=��̎1\�kp]V#���X�8����1���t��_G��L�N�m��k
p�A�l� �u���ɴy���Y����On��>�\��)��J:�n4���f�j7h�,�\2ل�/FJۃ��M���#�8��a��Y�ni�䈻����W��z������>�i��d�e���Q;�l�KS���a�8q���1��d2��kq}���o~s1ɐ�]l�@r�����jS9/X��"�����T�k5U�Ѽ��C&@e�WF� �=�P���8)#��r���� ����/��������.�>	@73��*����:�ZY����H�r/>�	^l����k�q~�tD{p�i��Og�x0CC�/������;�Q��2H���n�t�����1��A�P��4���e8��t�<�q�7���{�o���sԻ��2{��g~O����o?e�\ߟ�ĕѸ{����f|�����|�k˅����\�
�:�����y8f6�μt굝	����{�m���zj��]��|b7Jz���μ���Kʹ�׉Tm�֜焳�4����O�����51�c�#�a0�%���ó�w�$}PG�lz�����ڣs�߇
�o�D5��\t�Ч(C��I"R�ab���y<������*��+^�l�5쳨ȩ4�ǻ�#r^h�!�ͻo���B�uhC���]��`ؓ������9�;�Q�K���R3���0$)�U5	����1܄I���te��il&4�<&/��{L��FE�̣%��	Z`�v���9�yN�_���=�����z3z�Ϛ��?Ҍ��E���pʝ�v����f�x������
���9��X��ۚ���m�#�q���'\9����֠8=:�|��<���7~����4���;��4�?��?o��)f%m�IY:w�(�3j:Vs#VM����F�߹�2�є�������KG��[%O$�w���]k-��P0���
���j&5���� �;ᤖ�xp14�
�bFF�E��TԸ4�O��O���~&�@�@�p���Nk�q(�߶�J���f������E;���bAx4���X�i�H]t���<��Qr�#�K�A�5	��������w���~�����?����K�S*��iY'�����9ٽ����a�했("��rOs���6�Gn�kݽ;P�>�5�����DUtϰ�<@�eA <��jċA��y	q[ x 7j������aG��l��~�fr��4�w�^�R�_���i͍eȽ�������Ȣf�+>����t�jN�vP�Ŕ�İEǄ|�� ��2՟���Q󹧑�4��,�e�8F�4�Ȑ6R���<4f�B���!�.s�����G ����/�Ғc���1>0V����x�:qG�v<�� 	��ul6b� )�����ީCv�"�l�ߘ  ~ʻ�1���^}7�19'AY`�U�@t�\��d�!�|��w,S��\jr3��t���u2��Y�o�3��/�� 1�~���^������ ݶOp��xgtown�M8*�o7�G�zFɹ�l �f;*�C���#����>�eQ����B��17�g%�n�so�'�EHl7��t��$����7�a餱�\��\fB��aB�w<�a3�ԈV�9�<��"��1�E��v7X:!���Z�GbÛ���%ݘ�ٱ.06���s�S�����^FE1f�d�b)�S
��/@C���q�w͒��J�»�1,0\K�� ~1�LfW�y��� 'k����d�3o��t��:�lR��S�0'���,1�K%�a#����?��������z����^wa�&�>�w��J�/��Bw��x�1��]�7ˊT��g���g�����w�%��j^��� ��r/�'
1�=�)�c\�3F��YF%ԭ�u�6m�{���[!�#�5^:2U9��s%�ΏԞ3�že ¶sj`ϛ2�uKԚ`>_~��+�4<FM/#C|��}k��e��mb"�����$ţ�{ؖiu�����?#e��/���:���A4M�gU�}��h����3�5h������0�B!��+�����@�ö3x�;�b��h��ۖb�c���}�� x����m��ѓ.<Dmr�8�;X��$n�JD�X�G͠�l��>��lP^NS�I׃�Q��`p_��t�f��zp��C4K ��d-�bH�P�1�GC�D[�[��-l.\-q��$`bu�
�nw1-�=��Ym��g[��ܩ@k�Q�f��iw���s��<���!�u1x��>����Ӄ��6?�aT��}n�V*����i�_��q�#�E���J�vҪ��g�#Z�z��D�tg�*��E��`	��o����A{BG��K��E*p����g|�gM8�\�
k���f��Nx�N�����r]�cn<A�;L����ދ�[̎�����w}������9 �%-�����< �/%���h��?���+_�ʢ��Rq-@��~��=Scs�_k�7=1j+�K�r���d��~���Ƕ2�Ƌ���
��
`��j��<˵����h�]sZ4�/S��� �{���(��gy�����֦2ʡ�`yέ�'����9c�gE) ԰���ӌ�Ur+�?�Ll���m>Ǚ��l2l*��N�U��E��!dFڀ�mԎ���}3]�������Ԍ2�j�M*�:8j��j��1��.)��������F�x&�{��dg������ާ�|��|�ou��e
1�B�X�,i�j~��p�,��j���� M� �C?�C%<��D
3�S���?��'&+�I.����h5��w��.�5��:Zby��?�Utџ�����= ����pˍo���FK���g�9�3�-����V���)�j�L��0I�0.+��>�����2Y�{�[f*I� �IOhp�s3��J��#�����7��lG�-?����׼�5K��Tz���$�E>���b�
m��m��K��xi�Y���+~r="��{ǳ.(tp�4���`��J�7�s�< �����JQ�?���^^Ƽr�L�/����g�'�Ά�g��w<�@�Ώ���7�����*����'xȐ�*���w��;���4���}t�'W,O�TKr܈$��YIY��~�k�,i�vI9\�p�����V�yQ�0�?�5�^ĤP$8�F�q�d��i*譺f�}�l�xUƁ�pnJXg�7&ΝP�Ƕu�:�y'	tL���	��.�i��iZ�e�#ڌE���T�Q;�ְ�KL��{<�[) ��Ǳҡ*����^F���3��+��F�ʚe��D�v�],/�;�|6o{p$	bV�B�������i�����?�3������0�LWE g'?\ +�8mM�7�́�F��1:�t��y���=�I��a�mh�ĴP��輈�y�c���%h���+�2_�K�`1���G��iz�F^*��c_��p��w=o��%�2g{�U��YD��@ƕcV�ؕ�BVQ(�~�v�"�P;M�0��a��t��r����n�\f;�FX9?�#?��Ji)��:pI2L�V	�i��*��H��b�p�n@��P���Ң�br��Rk5ᲂ�g���U��'�������_�P���P�`i9�\�T^���2��5Ip'�k1>��P{p��1=���P���0��h���6�`�4�u��VJ`t�`;4�v��zƢ��h{��}�"F٠�>zTz3���db��n�i�7�V�!�b�!�����k�.�L�̶\�ӆN���r�]@�	�x31�	Ř�B2�`���w9���y����`&�P@m �$�[�p�EN���#���a�o��9���7\.r\��W�W˸�^
T�b����厵��� l��.#��;�]�c��e��y�}�����>�++�����e/{�T*��@+f�#�5	-�jD4*�5M��#�w������YrţXƲ!���@j�\S����'��m��?��&R�?��m9���<�v(WIŴ�a�ʦ]�UTø���7:R؇�rM��x`GM���M�0T�,��5�=���Ti��J{���&0ƨ+�1� �L@��z�s�*mRJD�L��ա���=���y�UϙV���z��h�EΒ���������^�e,o0j���Z�]�\kP��0���;w}�8��Y~�t��MтKxǨo�v�.+&B!Z.��I%�C��$�����,�+\H4�����E����y�M��AZ���k��f�[��҇�;)tA���i-��I���P����n 1�;]��d�,
1Q�<�9�z�C��@It`M4J���I�i�w�.f;��Ш5a�n�!:�se\i�}e�{��P����Y�6��&xL:�,���P�K>O�}���j�h�W��ssFDʂ�c��]ES\6�՚�����3ӄ��p���3���W��ʈ��s2c�3Q��Q{GjJ���Y��*|��M����琚�����UERyO�,������W�m@�O4_�MF�a�؋�D�Mmap�Z@֬~:I�^s���r׃�����Lh<9 ���@,�cxʺ�آq.�!6���>a���b�y�ա�X��N�^�>Ԫ�k��$�/�|�ŐI7/��6r�Ӿ�p�G[�|T�cvx�2�}�G�N�p��ֆ}������ߝ&m����;A;�]���7�H��5��^�]Ԑ�� 컬Ɩ ��S��[)����T) `�A)(O���ݖ9��Ox��ؾm��Eu��;��5�ub��2���;F��
E��ǭd��4G�z4�A�6v���vz�����]c��!"�-������_������DD�������DN��vI��(���J9���c�t�[-z��i��@� �7�םE�b���,i(5d;_��E�>L��:�Nt}
P�������n�?�9}bF��`::-ƣ��8�BS�`��{��y��OV����5̪y{-�L��_�М��:7�`x��]����&�f�qK6��k9p\�LS���˘�����s�H����0�����8w�ü�>�m�'_,�Ej�#�k��r�X����/[zxe4d۝Oh_i�:6�󜩮NNk	g(�f���]���4|Q-"'�I��z���8�?]�y��U�g���}e���6��� �S>��T�ѡej4
c�N	������ͱ�bg��eb���ye=�G��e��KIj�Y��Q�����V���gu(c.5r�F|9�etD�\��2�@O�i3�ޖ���%O��h��q��C��@Q4͐�Ԇ��o4oz�p^��#��Ϛ���y�� ���i�4��K��K�c5wK��S�`�������\��2�����bD�h��|&�F�  ����ʙv�K�#�A�I5O���%��s;~�0�q
�X3ƒ�ZL����bG��[�8VoV�<��c�;q(�����G�;��lMO{�\Zne�|ѓ<מ��6"W��I�ϲ�O��
7.�b���b��ˣ�~�i��Ѱ��臅9n�,5�a�m�.� \��aw�r���e��K9��n�䖘�8w�-)��I�֤SՍi[+ֹ����\��px��"��H� �n%�'��Lx�O+[ >*�Y��{���;� �Q�[��i����� d?�ղAT�tzѧZ�n��δ[!��!7"M��,؃�1���5�1��\k$�&b>hz�=n]�M6P6��D�"�^�,<}�dE�-o�Š�6�C���D%Tl�GD�FC��v	�}a���ۅm3�I'̇�����/'��B����$B�\��E�d}zɉd�~q�p���=�p�kE^��o��>���br͛>��p���b;�|2� 6����@�����������PD��!�v�����-�(��89�R���;u �R�����ùA��C��b'�\���4�hy'{�2jkz?3�z�j�E�[T�#��Eq�M�}�F�ѣ��0���Y�}�B�y�_Fß��S�-���:= ��5`�~���.�ğ]���xt�˄:ᤗ�#��0~�>����E�r�3���$9ae�o.�KI����n`�������Ҍ���Ck9�"�5zo�Ծ �D�Q	�BU���tgֵqLn��l���b�"�f�+�#��!�����q���06�Ś$r�ir���p���^ic�ϫ�,��y���5�d�<i�����}P
�+�޴_P�r����;ݻ�'���-�佾p�Z��� 0���$�� ��|?n�3 ��T�m�v�9�>�P}gҗ�$�����C�4�A�b�E� &���N��?G����wfJ�����H���=�f�<~����3�K��>w���,��E� ��O���L:�c����\�f�p�s�#<�� ba��n7�`cD����y�~�ﵵ[w9i��]>���Z�����T�<��r|��i!��>��n�	��^�e�|���yNrKZ�A���dY��6\�Or��4f�
�6bC��i/��ݝQ��b��w�"���?���w�u����'�3k^��Oo����ь�ԁ���p�0�@������=�KʳsQ6l�qGjMFG̗��)Q�W������/��Z�?|w��������,?������I��䈗V:F3�z2�u�s§s�<��wy��Z�~!��	��K��i{��/�}�jR�s7'�׺�%�!�Y�s�c	8�6|�½���IVpN���g_�&w�?�2+��"��$%j-T�uP)i8-��VM%N�M
"���m���ȉ <ߝ��	�1�o�C�Iz_Xo��v��m�Iǭ��Q�� ��: �
#y�cް��n4��N�8�s�\{��������']m���4�Ϛ��^�	�V�\����i���v��� O�uϸ�(�1!o	��.�Z�?$34��QҔ��4�����f1n�=6o����������h~Os��f�kÇo,9��l��� �@�X��Vk	�Y$E�:'�13��u�F���@.ԙݥFc���,j�	�j�����#�}e;Y�H:0����ZD�]�<�@&���t��/J�┅Z�BI�vͬ��\H|9Fe�s�1}&u�d�Ny��o���8!`6#'w4�!�)�|n��q������C0o4و	���`^���5���;�+��i�;�=�u <jw�G��7����o����G3��x�B�̺�8�+�;�3��<�#��֯Q�yo�1�='<ҟKi��W���qs}�j���,?�9���^�����Y?!M��:����	~5P����?3lP�H�tq�>Qs��djvu��<��J�El�s'H:�k�C���j�ׅlՂ��B���Ͽl˚]v�Q�~�����ĢTH�����\��K��9?Wj�w�B��4rr)˝���˻��VM�H��M �)���~q��d2e������}�}����
�ģ^����op��Bmt`�N̄�=>lf�Ǔ��mv�����G�R+�x1���f���
��;K�[,�s�{�f�=;��w�i����'�&��u��i�Bi��Y������8ps��䲉�����f� ��[J��Y���L�o|�hC��vI߇��{�+MZ�	5/�B�8 "��\�l�Զ��_��"Y�~��h��
㣎�Jg3�vG��K��M��']QYb��E�1�]�m�сK�7����M�aP���o����(�8�(��!	��,6y�^�]��i�;AH�k#S����D5L�;E��ܝ�N�j~v�Z�쀁Jڤ��N��G�C��I�7��l�[hD���yoëa^�O�JUƄ���3�#�ݻ�v�ּ[�g���M:�e��B�Lk0犝INZE
iS�\���F�Ms�|�n��H�I�$i 5�z�y-a?�HB��%��\���+;�����.�%�8�|������9fy��M�q�9�.�i���RY�]��x_����N�����H*��?Z�Z�\�S��R舝����qK��x�����g>�����MG� ��>��>�������	���Ex�z��M��'�w�]5����گ����4�ɚp�{s;'S��` D�:��o�S���v]с!pg�u�2��R�� x��h�B;�Hs���=�Kl_�lT���;*�w���I�N�E����vJ!z��I� s2���}վV��&�hN��$Qp��U�e���,���_u����[m�;��&X�;��L3������,�z7��zK:�8���g�{g�*��R�|�צ���5��`{�Qv����tW�a��S`?���
ճ�/���M�E{r 2�a}��=�䗣�R��偭t�dc0�͢!�E5/F�d@���|��k�v�-��}ٗ5�����R��S>�S������y�4���I�pߑ�i��'�)`6kv�t����$:���������6����N3ݙ���ʼb�K�q�媜7m{_簟sS�B�m�
�/F%�uP�.��,�:��R�S���2���a����i5��&D��I-+��UϷ�=]Xұ�.���;%A�62�$�$���~�Gf昚r}Q�I��#>na8�����pQ�8����He����X��۫�i����2�aB�)�d�L�y>nK����fo:��N;\4����m^���u ���D@��Q��t�uP�	UbB+6p�m�8��������������rr��. �M�m���B�,��Yq��Wq���i�;m�A7�4�����.���%��D�ᜦ�{�-���=M�h�(�[�7���^���34��B�L���g���M�U��i��U��8`O0������o}�Ȫw�%��:�v��V����,���*Kc���m׋��'}?��Ԁ��s�����)��җ����H��,T�wql��
�DBsF�d�$wJ�e��%DGt��|>k�by���^3� Z(+����̔!�A�3�*������AU��N��1Qu��hK/1�x��P���_~SQo���Tۏ��ਜ�j����̫�O�����Ng�����o~�E{���[��:��;P������������%�4U�<`	8���;8������B�4I*ƶ'u�Be����hĀ1��IB�B	g]xNք��j��3�ǣ^�EM�Q��}������=
Ʈ0�4B��3xd�EB�&�AS)�J�~��_] �M���Ƨ1�\f�1u���[��ǻH=AIRnոv�/���7��^���BD��C��98� p��Z�d�ִ�����hJ?�B*��	㬫�
�ˠ#��a��rŸq�F���o��  �8IDAT<�Tf"ځm���0��[���#�#<�+�u�t�����7���s@@������r�g}�g-CI|�4�.#Tf+[�ʭ*��|�(k�����1��~�`8b(���~"�=h8l`�N��p��ɗ�;:s,������I�LZ���7t2j�%=�{�:x �z�]@j;s��Y��Pb��N6VW>��>8����#/~�~��m8�ʩI������l�NK ��(���r��}�k�e���5�w�,�T�����"�YsM}N��3�;P�4_��k ��U�$�����9��\x�p;u�(���7��~�}�'�:�������Yіm(x^�u�4@�W Z�i^�"����%������s�G�u��	��2ƶ������܇�D��bf�z6 _АZ��V
x�N˄��`����%�ŀ�5˥22�c�j ���,
���K��&��ɧ���-/��ݴ�_�E��G�kK\kF+���Z'"y�	�ѐ��Фx��^V��[���Y�X�X����7��7�r��l��9�7���w|�w���/� �@x���%��_���Zǉ-�&�
�%X�ߌ��c��L�87&6�
�������	��S�_�҈W:�,9�ڝ\)���X����I�z�Ь.�+�aŒ�5��h	V+ N��<��f��ߒ�6���[��V�N1�
�{��{
�����/�b�-�jf�~z�DVN3٪�H�6g,�a��>�]{-��gC^f<N�����S��;���N�"܃���馂�1�j�� �4�2�����_����T���%���|��}]��w��$f�[Cs��L-�bH���L��<uH���V�陕����.q�Dc����J��������YW[�P�Lٖ"UcN�0����:8Y�,���>���1[�m'��A�ӄg��br6k��%���],_\�4r��Y�%�=�43���2���46ǲ*q/�l�]����5��R�[�V/�R��W������r�ŰS��o��o]�����I?��?\xa�1�ŐUƳU�bUVf��U0ӿ�gfg���h|�i���|ҩ���4�~�o6_`��?�c�E����T_�H�p��2كP�Cd5����IK�	w�&�U�LIEn��[H���*c*�"wB�me+`���"�o��-�up�8 ��1�82��v-A,q��\�Y�ĲL'g�s��6��������.�H?��фǋ�f��7tܙF�~bfn��d����0�Y��!���;���<�aú�}jv���G�c�
	�:u�2����h8Hub�m�D)����W =�������:�M���`��q ̼c��=��J��
^bG�p�ω�H���ѩ�d>8(qo�A�b�2�#�������.'1 JL���^J_*�T$�1/ $�wӎ�C�')�/zыJb�;�����A��?��%�.k#wJ�F�$y�e��4���
���uի�l�N7�k���ې2/�~��?�ap�}�H9F�Cy��%b�,�Ԁ�^�{qOl��<�E�҇T���9u� <�L
'Oˍy����J�i���������v��� ��FLа� jf�$8Ǒ����庿�+�R���ჸ�O��O���[��vq�����z#�=k�[�\�$%�8��.h�#j�y�o�v�c,`,���H����g^���{�W��������*��C�y��=x�&�3�����Ek£�ɂ�����;�� �GԼ�%/*�����Z�&i$�<��/G�9߬:���9נ���C?�C�Ꮉ> N�Q�Z:��ِ�ŝ!��N���mk.[꺳��1�u���lǭl�v�������5b�`�%m֬�e����峟���(ו�����k<C���!^��6��]<'\d�� z��~�l"�����R��*`4/'��Cb����2��|�;���w��h�hŖ�C�u���3�3���@�u>5��'��� �I��饈N���[�����ϭl�v
 ����D�*�H��IOHk䄶RR�ϠM��Jk4i	�Ȑ�/�!1��#ΝA�l�g�XM�ݖ*���}6� �����/��n�����aš6DF �2 �/�JĊB���x�;�F��I 2��r��gl��w�hq�9Y�5;~�6�񻹘}������s2�7-,���=ϩ��u0V�#�Fw�c�N�,c{�ql�VF�tv��oDQ��qj��o��ͺ�j�uq���V�������}��ssN��E���ķĮ`=
%�ό��1���=
#�FFP�E�"�5�%����e�V6iܿ޼�mo���tB8xV@چ�Ù�j��􆚜D�(������K��`K� br���D��u2����;�7�r��sq�kC���1�.|Zr��c�tp��ǖW>Y쟌2��>5�&��C#mr�U���fƙ�Mnt���Y�ܸ-ʼg�Iw�B-�*�?�����'�z-[���8 L�b�S#���kv�\������:�g�t�u����l����?��#�[���t�E�<^���v�蒇DtX��J��a�!�u�B�X~�Ŀ�:Y��8x�>G�mp���p�R&T`�3:�B��Ӟ����;�io��a���0���$˰
~��c�mM���m�̳�U�;�ᣵ��sX2���(�˦��+RR� 1�Nm��;� ����	��o\Ì��C8���N[@JCw�`6�u6-q�t��6�z]V���	��4_�� R�_~ZH�0���LM
����?��>�Bl(���S ����Ǧ��h���)a���$˪P�	�����:���83N���[��2�O���'_oi��ՒTD����C@�Vn�ASŇ��"���.�ck�Uy��L���n�P�V�����P*�����r���v�1�Yˡ���>�3�Մg�Cs�lO9��sf�������QhN��fϹ���P�P�"�/���Pǝ+:���,j��+�A2�G�2���Ƴ��L��(GԂ�ГRpR&H��jBjdy"OK��vK u�d��mm�Q����8�9�F�d��}�{�of���;��P����Q��,J��q���2����
��#k�Ǔnb�݇�Eg֌8�8�bjV�F�\�n���P	��Eٱ�������F�3w;�l�����d��YR�uPІ,2~����`�@����ȅ���\͊���̫�3��]��'����r�d;ٞ��Z�i�G��s"��a
 �Fm�
�^W�Ns.y�[�;��U���cbP��!���$~^Y�&�|s0T�o���&�/sV�ɲ�R3e9)�Ԩ����N�8�&#�	W�1�.��!��%s�����9x�^�PVQjA�'��馆�3�6k���\�j��EZɶ�|���C���%WK�'��ɬr���K��y�_���r���s|5�#�A)�2!���5	�i�;U����4��R�]�R����Vd�^����m��~��_��(��v�9��`������t*�J(Hy��k�����t�X�����8����U�:	�j�`�8��LS|&)��RMi����F@\)J�E_�E��=���_�Ņ�$�	���>j����ٟ-��'8�������O~�G�p�ܓh�/��/)�d�
R��>[�q<B��ù8���?�G��	M�Yu7�--s������\o��*�-����F�i�;����9��V>Xƨ�C.��'�*0�O.�����$~w^Y��o��4�\��t.�1��̂�h8��p�2����㽒FpM*'c/�(\\��<v���J�p\^���w�� +٠�����Xw�=I��ⳟ\��c�[�1�a����'~∖Hb�ԡ�������<�9��#��ׯ��M�茉��a;��՟g[{~M�&�+fy��A�\��+�ͳr�浪�k9)S���M����k��e˺{��K>0=��<���Ϡp&h�
��L���J�w�Iih=x�4�r˗�����i��} w��2�vff8���q��X0�S��Z�E��aI��ß�q±V1D��c䀴�kh���1�9|�3�9�IH�c�A�A8�>�$�#���	�F�
��!}*z:Jk�RNP�.O�D��l����7�Vk����.����t���'�"��QF� �9R[�~�����{r.&*�I~�~C��ⰽ1w�(ը�q���f1~<K�;mHf�UZA�*�Nz,��m����IL6��	{-�<B]�P}����w�w����k���; �FIIYƃ�gL*ڷ�]2��O��1α�c��ˤ���w����H^���s��+�z-k��p
I-�ּ�9��Ԁ{���y:EM(� �4��Pe�0ǺK,@�Y�ɑ< }ҳ:�QKKm<�ޘ������[�*9λ%��2%Cǵڙf~�������~D� ���G �L�1��G]&�p.�e��yܗ�\Is�9:c�ύ�ВJ�t�j�Y���3lS۳NF��͘�\(<&�U~�S>��o�����Z�����*� K�S����.��v$�Y��EI�Ey������('�geC��s�F�A��	S��4M����-	&���~�`�4�k��s�A���:�z�5�Z�C2��.p�v+o�5��0����ukǩ�K:˱!�����*�z?�,A�E��������V���Nj��LJ���'>m�u/:E�b�7��k�YtrH��>Y6z�2v@���1�N��N��V�:�x���H���Ni =�H��1	�|D+v��jY���I���#��W�hz� �O�x���x����xԴ��2�;O�Im��ԨS�κ"��L�3z^��˒��6+7_W�������]��T�VaIM���*'^Ƹ��k _��%.x���Ό�'�Ho��7������\�O�o���E&c�0�:���8��PA��M�8���G\�8�D��ƩV0��� �1�P���t�5��L���>w,q�z-��'��I��*�OC`�����9�)x^���B�b�j�� �v�SJ �tw�����HW�{�3��g���4�l:�\rK3۹�z��<�ݥ\�l����E����OG�ٸnM��>H�8���`�[x��ɚ�hi��t�|���ef��	�p���s��UrA��v�Zc�T����F�{���fD%q�$@L;F��3� �"'5�V�-����w���^ku��U+���T�L�������2P�E��L�zQ�컼�3�OGlƆƘN�|���ZWY^���w�s���B. 0sE�2��2��4~��Oȅ�~�����N��'�����4���v��ݹ���{��r�nI[p	"�2/d�<WhӌyA��QIM�I�LS����� Nэ/��//�������'b�d]��$�Ok�KG+���ns��}?�>ۛ6��t��-��9�)��Pg��� ��D�	��������` R�/�K�3XX�X�l3\K]��JC$հ�$�w%��ꐷ\ 385�4��G ^e�
����ч����>�<A���@j DRK��p����XJG~Xm��E:-)�ia��-L���_�y$�`������K<<�s�g|�{�S
�[�tM�B��^Q"�S?�So��N_��'`��F��]�\�cn�mG�Ō����W��> 7[6�������/~IE���ښ� ��S����~����J�4 ���w$L)����%��/���{��	�����e�y�M7��r~�Yo�B�/9Ư=�ؒ�-Z�@8If�ġ-�R�Z����'�������>�nU:��j-hS����[/�d�ߵT�.Gj��P"�Y���5��x�L�I*$��y���~~������!iiy���Tº9ʱ�!衇J��ׯ}�k��ء�q
�K�x����QI�^�E|��F�7(@`���������e
A���x9 ���Z�A��r�8�[z�\}����>�SK�#;k��`�g����|тY�ȼa%�;���=/%��r?�Nxӛ�TJ(�n�V'�|_�_P��k
�9��l�U��xܛ�A}Q:ig��r�פ�>��?=R�����se�E�J$��=�yw_ϡk��ng�^fA8��4VDS�v�n���gc@q-��o��� X�TIJ����N�MP^j�`���v|$�'�@�@=��Z�H�@
C�Pm��pN�ǉ�%&A��oy�[�_��_+������%��X+0�(o� ,�E$�0Wğ���^���<P��^h�(��/��pٸ���&P)�1�+l;��M�Ox�S� n�$�x����Լ4{=�>�`���K�����<���/��/��|ei|�C�(���ȁ�N,�!��9�~k;^�nǤCE�L���8�a�����2#�`zd��r� �9��^k�h����\׺��,@[�<��Lzhk7H90��Eӂ3�,=�5�Z��:�2�;�65b?CR�^E{(*�akc�:��������ƨפ}��Ѐ�!N�3�s��{���s?�s��@��uH�� �@�{�mso����ŌfЄ/>:b>oG�Q;�ﴺa�y��>��E����������ұc\�������.Z-ׁw��0s`���W�������������u�5��ۿ��vr=���`�I��1�-�Ef1_,�Y����>��`���W�H��m�sZ¸]ہ����:h�<��a]�WϺ}ķW���x�+
 1���hY*lO��0��p��HWq�5@��K���\����1T/��T��	|x��_]ޑ9��7�qI�!���! �Ջe���i_��_ۼ��/l~��~�Ȃ��8ݠ `����Y U�2$�y(����;�8R�����^�L�I��:��p��Bf�<�'�q����bGs�Q-�FD�G��]�h(�;����
Au�4�4)���q�#��'I�tZ^���[�����ɖ�v��mM��l�hLLV)��t\�Wڅ�-��q�il�[/9�����4]M7	��0�|q�*][��W���	���F�6���^#�?3��Hϫ�jA�q���ь��]7G9������?+`
}/�jz�g�*v�Y�g��B�s��SN���P�xVh���������£#J�·jF�U���"X��qGd ӎ����P�<y9h	���
�'Z N3~%�/��\n��},��8�J���&��`�rq��g�.u0�q�d�����m�3=�I2�����dMm���{�+�fT���ٛ8'�r1��9�%��@���1� J�/�̾7�\^�qa8b��9�~g�U.� �1�>�4���u�k���ƍ�"�	��������jhj��,U�r��bA �Rp��4��d�{�myN~�b�9y/���vHŅ�΀W��^�aT��Թ���xM����vԍ�7�O���%R�/��/����� �أ!;8r[mX�I�ՄՍ�	��c�p��ꒋ1"������t�����!W��˭M��צ]���`�M��}��L+A 6D-���5���9�����x߭�:���e"��$����XT�
C>��`� � ���k��q�5���Z�
�s�I4�S��sƏ�w��~'���m�F�M�彩m̽P��`�u���=$yӥ}�
��O@5�����5�p�C:�td���� ��f�Z9D�ݳ\�&܎ǋŌ������%yHwS��r���ꏨ�f�$�J&�/�@W��x���vN;�ḁϲI���X��$�L��<Y���Y,��4j\�;��_?��hP���$t~~��T�`5�w�����$Ƿ��/����C��U\k��wU0��r��ߌy�_p�������,�c|y�t�^ř �o�����Q�Q$�)���D'�ǻ�.���,�/?mCA�6b�ءu�����}M���IR�`,%��Y+�Q��X0b��3�ɚ𸃠Yߐ��t��/6��4�SK�������CK`��R�v��0� ?9^���gpX�����zQ�Y�<��\�.,.����`)�.L(�52`~+�#u��N4�c�Ɋ���N��ܼ��� �J�;d�QFZ�^��#�d��?F�V�L�b�G 7�%�@��e�C�N�x�Q8(@��M�1�y3yV ؈��`��}w?��:-���W9@ՄYDT�2cϮ��Ԁs2Oǅm.qjM�ǒ�WV��<���e��ڹw��X� �+�����?���\��\���fŦ�����^aޖ`������,׋��]����}D:M�m�6t��5li'ʖ���6ʶC(/(
�UyWw#G��DH����43J&3��Y.|�Id4����^�4�|R�D�Pj��9��h���-�R���f�$�2��:�8(�����k��۾� ��~�����A��$�+��
O:@]��R��`�-�
�]��7:||<�`O��0�:h`�Q��R�e���f���������+��e_�A���(��� `��P3�s>˼yM�;Y䆙���&j�f��r�:<՘�����r+�+iN�4?1�	äo��˘Գ�Z�*mڟ'��B�T��7p?(�l	��?s���� -�3︟<�ڦ�8�7b��!��I�x��Fn�u��E%CF�K^����n��2��cwIg�JMǩH&Xg�"�[Z(����h���2�#�N؆��E01>����_:\4R��d;��A`�[�<�,�#�*�*�i�I=����Ⱥ�C4��PB�<����|6_:�)�����M�IN���{k	l���Em���(c葤ҩ�<I�J�	�1;�8s���"B>ǌ�F�.U�5��\���u��h�@F:��D����9o{��ʻ���>����P2���]��<3eP�W�+��j�$�����g�3��L:�J�?��c�D>���IZp�fzVYi�?�>�-�
���IEh��j�?�L~�!<0Vd��42���nI@�M�G�Nq�����=�@�=C��`�� �3������6�e�7z+�#�8a<耡cے�I���* ��;rHUf(�	[����w3+O��s&���q�Xs���*�������KA�����N\'�$܋g{��87���L�������,�����b�3D��YT�Ѩw��j�b6g�l'��h<-�0�>*3��?��J�����Y� )�j����rMz=��㚬pi�	@\�e/{Y�Q�F��Ȭ�Հ3f�,�W���������P��uO8���(��*���'��i�M[�3DK&)�4<J8�ag�(>g��%�̶�?����1����jق0���6��|��*@�ʔJV��Y;ƨ�\�|דD����zы^TƸad +��Q7Դ��-Fy�y~�s2輇�6-m��E�� '!�p�>r����k�	�%��N��� �>�����q�16.�A�`ry)_F�$7����А�wr�v*�!�y�k��C�;���0��?�S?�ܜ03��(M��e�y��̠2�Î7
BK��� 1aP�`�Y�t[�\Y�	�L^�P1��΅$-!�M�C[�\��Q�I��r[$5W~瘴l��� 67x徆�ɍf0�OJ�N�� ~9eD�.��8� �o��on|��bU�) 	�5�_���F� ^p<ֳ�������Z���%X��y�p�����͞A6J[��R:����L2L�O��Oj^��7ׯ�h>��?[�4���1�P**�����dU�=�Ƥb�����\)%G�Y��%7�xa;T�G�k3���@����9"�nQ��J��7*e�W�ˊ��N�\�5!�Y�G�8,`�NS��K���[���%#�$�o�"B,�W �����sė.�A�2 :��GY�s��	#�1p�`1GTPL쑣U[�Ӥ�zj��=�q���|S���Y  MFYB����u���
j�0������%>ڭ��ƿ뻾���;���e��1�F��rQ����,���r����Fb����5
^i�̦VM\����LZ�����a���d�����B�JY��O�����q`����6��%f���T&~�`��>v�&�⬐�X.iBls�r�i@;�lp}�\[���5��jIj5���8�@|���[��!���B��5r����A�t^�Y.�~�w�c�t�E"ǔ\*���sF$�J{dd��ajZ�|f�7c׹�U�)I�<+`��=�,
�S�V����=`���������u�ٗ���<�=�G#ϑ{?*�M�j��0�'�xtu�����_X^�	~%�Z ���Fc�Γ��@ ��uY�seup
�TMm��1���s@� �^�Z��Y������iz���j�i�aj���).Vj�75b@�j_��4uP'sMMX�~�1�Y_�- ���7���R���&�dn� ��s,�;[j�9�� H�$����AQ@Q�XY2V�_��Hh	C89��uZMe�IV#�|� �r�(��םj�<�s-B]��rĵr6�0���q����9��a�R���RM/�h~���<�h������bL��#Y�So,�Aʳf���������4�\Y�h��O��2����߮�6��(i�;Y��u�����Tn�%��EMg����E��4߭6|�Z`~F)V�m�X�:��R3<����  cq��q�?"˛r� z.�)�����e>����DI�5����\��ID%'��8�����7,'�����gý��wJ��1*-Fx���蘗�U�ח��y�CX��[k%�yoF3t�	�3q%�B��.��8�Y����W�Q_��o}�[�g�z�;%�Y�p��Sǂ�W��;��;CE\��m�d�K�!�J}7�h����!���?�>�1Ъ���-�!x� ߂��K�iMI�S��T�b_e���r,> �հDnnmeqr^�%�|�'�����ź��^�X3�6钌D�8Dʄ��[�%�㴐O9k�q,�<���:�sg񌭷x�A�0Ϩ�F`@�oJO��j����L�B*�=������7��1x;Tt��̧C
s�!ӱ�(A�����6��3�:�ģQ�D�z1��a���d�Ϡ�SNX��n ��q�vЛ�o8��9�,p#�ʨ���q�p�[	w���Ο�{ Tm13��.J-1N�qo|-�`h-�1�8�9f� (f���%c-w~q����_����n��c�z�'	mF���_���/��k[a��q���A8,�:X�?�EF����+�˱�k�$�������x|I!j8�\yv&}��^�sZ��+�������%����-���m9a���@q�M' �j�)ʧ���}�<8�L���Pc�����Lj5�h�	C?p�Zj�m+�c	��Nt���'����ݿ+��$p��4�jpy�:
�I�ǹ"`"����%�u9�,6��kX�Q�Z�>���~��o��r]�b���vQYWV�(Ƴ���F2�X ����S9�����` �)��iY�FP\��Yݝ�c���ɝfہ�������`r,A@U^�%M$�a!�& vb��� ���}�W�t��ۮ��b'Y@�Z�f5�����t&X��N�೚�C��{9RO��Y0�w�&
?L*�+�i�,��:�>S�SMm/�8X:�̮�Tz ��,c�}7��3��g��vN�$�/Ǡ�RF�9XN闬֦��u,�mq�,��s/J�I�A*ù�iھc.��8�xN��N��y� �Ĺ.��nz��>IRz9��,a�������&�ф�����軓%#4L�*9?8q&�+sZ��[�X3��)�#ﵕ��U���p�Ϛ��@k�&�"�R���C�{�/%?�|5O�RƔuX�_��{�Np�P�E�c�C�;D�X�`O��Ys�1��o�[`F?����*`f�|i��'��nV����\VY'��(�ssQƣҿ�ч�H���uWb�b�fQ��j��R#1[��;�ZD������V.Oj�A����c�!�t@��zr��
��HM1��R4�����ȥ��G����s�i��ؤ�q�=�������1ƽ���:M8ۢ�<\���(�~�����*�Z��(e��C��ƹ�dg��]܆9�(N&$'nz�kn�E*M�Ui+�:�A�OXT-5��H�B�֨\p9�T����:,��@̤���\�	��Ka��
�z�9�D6�Y�T�ۈ	�I� ZgY;Bz�{?���=�(-��Ƽ��P����2��q�^����c�&�n��� ��C~M�;�6�E�9�
�#F�j@��A=8�<�֞��VҏwI���-��c�41iUHZ�u�0 9F�u,���Z�TcG�㽾��ݑ[N@�FEj�n��C�{fVYf�%���]8�gH��\f�'�h�7���n.�g�� ������p �5���w; #�N�Bm�d�4�2?�ZH=�:u+�'�8F�'1�>�`� ������4r�[6��u#�w��Aҁ��?������+_j"�[()?ñ�ְP�Mm^P`��z�e(NIH���+�
�Wq��%�h�+5�Kq̝Vj �H�U���� ��Ť�T3�����ñ`VyJsP�N���H�' KG���/^�n����yV�c� sg�?�O���cܬ�5��rH��2�<���&/�q(S��2ؑ?MFk��*,�`|�r"/f�3��EM��#��}�� �`��"߭�b�tC��sn����\�V.WrqK>���2��H�7����ke�ǆ�R֞6�غ���9��v�����@VU�y�ȵ������PM'��s�C�;<6kN��:���JXu�Eʺ{]�p2O��-屲�1w)�d]U3�6	q��r<mb&��5�g�{��I�d�a2�I�)�U�����L��&��ˑ$
?#q���n�Ԥj�Q�5ـ1a�+=���6���ƕ#��qh��,Uh�E�.˙����sezr��Ҏ�t̩A�I���6$�$	������Eh_\4W|�ս
����6�4�ɸ%A�d������ Ð%wp���.��z@Mذd��9 WZ��U$�]}X/}�KK}
��	��Q�p��ʽ�61UD�\���ǥ*0m>��NI��o���/��|�V�c�=L�ɰC��^S.?7�o&��l�1`�	7�x����W�$������L4��*O|����
�l�U�;�l�[��)�Ǜ�f+گގ�	1?2Hm��'Z����~�k���e�;�ȝ5���*�H֡ �~��8���F�P��1@d�7��:/���;e >��3�[R���D��hՀ�:��G>�4qd�L�����_��R���g����4,/kf : 3�ٍM]��/]h<��f�fX 2��u�S+'���h����P���O*{��5ݐ�+]��s�� �i$�kG�O.� 3���Ea���u�+;�ґ=d�x�[����/�r���^��ׅ�$Ȩ]��ec��z�q�wX��k��֯�t���B�!�@�?���`��SǍ��u�Xx��q9���t�w$����K�dD��R�H�wr�逳�+0�u��3N��05A�k�E���o*9�Z�!o\�qc��J�*m�~G��̴h��X���:�d|��D]bv�aAr/F�CF����h�:2"(�Z����Va��#(4�3�E���g6�IJ�~PЄ��O�ce-'|p���C��bC��i�Xn<�	���E�ç��{�!��f��"/(�MU#4ƕdg�׽���m���7ӎ�B����z�j�j_f��~x�x�+W�݌;���f��3lĸj+��+y�ޔmۣ!Grq��j<��I�k���A.F\ۺ���1���ܚP.Y�$(�=���M�w�x,��ϡ{T�=��I;��G�8�������~��e����sj��t3O~������Sk6�LcK�q�x�(�`��;�V�����U�Z.����)�j)��\��I~����!������&Ub�r_+�Y����(�jÙ�9��9��h�`T�Q'ֳ��;��-�OGts����ޛ ݚ������t��!	�$l@.*�6(� �BDEL0�������[7Cݾ7�R�U^��X
j;&�hd0� *�DTEiA���3|�������o�o�=������~N���;�w�g=���4G���p���zsn8F�W��k��?�K(A��X�Y7t�L�=��O.������d�������Jg�@�T0�w�wO�Uy���������'��Ex�x0��d���K�����;��5��N�����e�s���>��W�bȓ����U��f��z����1��l

Q��I��@�Ș�$NA��~-�35�ǲ�����4�=X��]=#��X5'4��Ve�-��1WT�E�u�Y��H55�� (��/(�A��>P4V�Vf��#���ۻ�����\���F��3�)�ڎ)��Iyű�#_��fO^�A�7���V��؊��1l�]+|{���]5ƶ�b7�J����]߮&�����
�-E��*B�΢H;��f��#`r�z���������A�n��Ğ���G
l����,���:LT�Z�(�ۋ
���},�a��� '�,���9�sk��	 *��6M���gx	d?���}'Ha4�Co|��LD��r��,T�"� "�GU�fi[�E� f������e�Ls���-���w����.|��r,fgϻl��EH^\ೡ8�Af .+; ��gb�a�j��;M��	��K_�Ҳ8P������9���;4@�Ƚ ����<es�v-^z�$̆vk��\3������U�yl��O�y11�r���b��J�<�iO+*�z���7�,��t������j����z�"J�ű����ѽ�6�s,�@#[S{�^i:��À�.��%���/��0�j+2L���l���,lT;N�=��)@E�u��h�`L'�0��Ƈ�Fd���J�4�\L���	M��/���b�ӱ�=,��o�!� *���Y#�%5q%��Gi�RXr����q�(#ҙ����؏��t�2�r�P��"�ǋE�?�ma�f�/��S����l�rL�*�jM�j��J-s�$�4c�b���Y���ۄWV����䳞�����|�����:|�Cz@>,� A���Z�0P_�Aa"S�=+X�V
M�"��U*�c��(Tā��3)���p���8�m�'kH�����Z1�d��DӪt��չ`m��D�h�n#L���X�H��qW%�}����2OL�}���Mۅ�f|ޮ1n�c�b0�>_ބ BK��.+�ȍ?%~��$���c��Sё����4K�\�	�Z���s�8�M^�M��z1�o��V�	��	p�����s\{�E�
�D���at�&M}B���Q��R�L�{j.�A8͟���*��h�����q��Ak뭀�:?U�VWNs+jB�����<���p���8�`x7yP���v�+�+���EG�h�߻�S��.�t`���p�����k��%ӯ��������ӎ�;s�3�4md�����N ��ԩQ,zv�B4Mc���d�h��plB�9ǋ��mn���ow[��s\��"�[�h���X���7���T��N��b�SV�ct�)ɂ��ղ��(@�����\,f9���{k�P�z~֙�3tK\�g���6^�;}'�d�ۜA�~�`l����9��W���1��M{��z���]d��L2���� �)~�l�y�D;	���Eă�UV$�icU�h��u؉X�AԬv"?����HWAC�M������P��`�9��Ύ[*Mz�8��w�h6�S����6���ȏt��#���R�K�㱪��&B��$�c�H��`Z�k|��O?�я)����G�3���w��	�V���y�4���`�$�D_��ѧL
����3�!U\7.�f�H���q�F��lc"�4�-
�����n
8�4NI�.���~��F,��\�}&����U`:O���D:�;�09�w���Y<�ߐ+h�FY]��-����b�����ћ#�M����Fsթ�J�/�ˆ�A8�0d�Y�B�blN<��AxX&:Bt�Ȥ�qH�
����Y��o,�@��6�;��`:�cJa�6VQ��ɐ����n�v���X�j�B�	��� ��Ƞ�2ݽ��6�K^P�.�BȀ���n�i�;K��RMN�h��Z�g�i�7:22I�K��+_���=�cxG�Y_8��y��w�}�k���'�3�k!;@�P�\h>�}Ӂσ�%��q�]�V��'���:��3g�96���7G��PV����0l�P�����I�]疓8�aVI2X�ϱf:����0
B��;�u��7xn�3z\���H!4�j[e���.s��Y�=��7��Z}��L��|��2���e�l�{��a,�w�Z�?*���U�y-2��^���ٽ��,��DE���U���dY�}���s�}mҪ���~�g�h�|���F�#7�]6?�!@��_�C�r��aH��A �!�-��R�4|-ې�ؤ�L�0��(/�ى�2�'�^���5��/W#+si۲��0P������k�f�'I���Y:��/��0�����ogz�3����"���6�Ӆ	�&�&�D���03Q�N(��wm˽u>�6@������~� Nހ@�?�3?S�Ђ��L�:��� d@��K��<^I�\����F�K?DF������4e���]3ID��?����<��uו�c�E>`�@&������a��)� M���KS��nD���1��ʨ�9*�\Ͷ7�J�'�c*U ;6���������]>���-���(��,�j��ʢ#�Wņs�_���j$�E�μk؍�&�"X����*���1��ܓ�g˶�*}�_�2��q;w�t2�L7�dL��ݰ*�h[�\���X5��`a4"���P��K]LˮwP��E���F�(�(�^��-� ���_��.�i��o~sɠ���^f�M��Yo�vQ��v��?�M~��ʶQ�	�-�0�o��n���ډ�����X��)ҭ�R�@Ⱥ��!%; ��9�/� ����-E���5(;���=(�=���U�h��L0��Ô|�Ȕ夽h�_� ��hpb����#4��H��Ʋ�4Ҍ�=��@''<���U ��(���p=
azR�e�C��W���{��	c�	�z���9 ���E-�23
�N����N��R}+�Vy?*e���y,�	��[y�o4��&̱A<��
z�賙v~�'ծ���F{M�W.O{&�p����;G��_򒗔�#I���
��J�o4��{��.�S3��(�8N���R��a9��ن����k%�l<����`�C��횒2���?H�4�X-0���B�������B蘧V�� ��\�UuI8�įx�+J�Z��܃,6��sMl�fM��g�d��R�T���e��<�����i��-�뭴S��s��h0NW�;n�� .T_���<NQZ�M%�	������d����
c�;�!���U��&ev��?���k�gr�D<���7���\���f����na�<�ϻ�գ�������6����A<&� �Ǥ�Y�E�E6�Y8�M�����"G5fA���Y&�M�RF�)�c��(:�ع��}�|o�">�o� ������S�f�c�MԨ�>��h��r��-S0�{���)LxV�k����*�u�ݍ�zt �T��P�l�"4B�����<k��,B8kxʼzD�CN�ݝ׻ݽL�2���T���.�%]qFB�餃���R�jgdڻ�}����{������S%�����{
�#�����׷��嶟7'����v���+��~�n���"�����#$U�4���Ѱ���D���0���|�)�L�wz�H��KAݠ �j��5@q��F3�<�U��V������=�3�B��I&�B4lL���BK��6i �}S��i�0s�e>����~�b�G�^Ď�G,�� 1�Fަ��o�����^]�e��n��]�J�C�)@e����O��v�Q��ʫGgPro+�$�ێ��(�S�;.��i��e-{��8�����O�Y��/�՞k��2�D3��&v����,��A���pVPf�}��ש�h��qg��eV�jw�I!��f�x�W:��\h��wF,��E�y�����6��5�<��ܡ���%h�nLR��c�U#\���>��	��w�q�c�&�c*g��>Xm����J�i�I;��"4���ͫKt�g>�?�9�
ܜ��e`�D0�v>����ʕ��_��W��=n��꫋�x\Rs�tG�F��%]W�㤌M���z@��5�J�c�C�6��s�E�{Ht��̅ӱ��@�z�T��m�ud��, q^���] 8�{��ģ�a������ݑ]8D��v��6-+#ۅ����e/+�e����E%���!J���[M���S��a�G�Z���1�����\��SI�Y��-����	S�b�5��}a�6Cm�G=��%n���G�:�!�>(�/B�L94ˊ�	"���H���/.i�=&>uEA�T�'F�X�D����b��B���b��R���ksE�zҧ��ʦ��k�v^�7mf��QL��;�%师L�]O&�1� [�Y���A|�pD�����^�c�
�y�!� ��Q(���zU�D�Tl$s��0)�.L��Fq��F1�,N$?�W���V�>چ�=���1�R$��}��G�?�%������kvw� te�\�3Ep"����q�dh��"�R�[��L
%�9�)��r�������X�7��=>򑏔�,jU���U�z���/�ʖH�Kq���:k.B�ƐH �U��y��[� ��S�{��Jb-�=f��� $*��|Ϝ�t���"!� cY+�ۨ@��A|F���r<s�v�2]��y�5��(ؤ����,��M�Bc��_����D*f�c���e)Y�� %� SBa�[@����枤]�<�?�pݤc��6Gee�N��-%yb�D��続�?���.� 0B�,��at����A ����P'&�c�Q\����F3MWۙ�<M![hCU]�]�N�z��C0k�f5�bW���/m}�������B)l�SC����S�0�R�[)��ַ���[��"8���7�s$Z���b^q-�^��W4��?���LJ-�Ë\��o�!��;���M<>�������Y�/��/ԙ6�����ۿ�|�h �gĉfv-u"xVk##{�~]�X����h���g���ݐNw�D�`�@�q|ڝ��I+���Bx@�Q���&�s�O�6��qkY]>��/��-x8:,��
F��3�nR�v�D��M���6��Yp�O�QR�J�!C_L�>���ժ��n.�.�D����t%W}��R�Hdz�k��R�?�)�cjB9���5���(��Nt��f�|��8�����qJY��y��h�F"���\�hv@����|���)�!�)"Rw�ܛ>@���2������E�z�օ����	��Dv�!�耢s#T�5`���?C�l�Q��R	E�ⲫRЮ(%�u��Xcu����&HT%��4�cݞ����!H�ņ�I��G��o��b��ZT]���<P�5�3U9=��t|����"��v^��MӁ�c��^���)8�n��v>� S-t�o���`3��cR�}
��Qȝ!8�H�x�32�4��_CHQ�-t�-���)�W�)�ۍJ��`����h�����o�뻾��0i�*h8ܨ��%s��ұ�9}�s#G �`)���	�J<2�_���Q.����uD.��)��;�wW��JO�����>����ǉ��|i0O�J���5�#��]��0��~闦�`Z0^���A]�� ~ғ�����e�����#�fy�Y�e����<���y�9�	y�Ь~��T��\����'��K�~J6��o,��Ŝ�0��O����
#��bYF�ٽ�mo+�F��s 4�!,�� &:	r;M�鼭�$�W����q�")ʠt"" _f�������E����W�(R(sM^,PԞ�gʫ4:N.��$q�M�m;�:4LIU��ϕ���;褁�(��Ƴ	��0M���5�3�-��=�N�qڮ.��㦋�?���q��(h��;�EW"*�~���A�|��v;,�55ZH�� "~V�[{49��
A�����s�"D�%�a�-��=�g��X� j�̡4�%R�G
մ'_u1��1���_�j�T?P�	j�g�.���!Wڬ��a���bǪf�}t_�e������A����Ԁ&6e&�d���:�B4�ݗ��<Um���&�r5)�Paw��8�.K�b�l%�ˍ&2�Ӆ#�\��ϟ}��jW�h\J�w�!j[$ktk����O��X�+�fP��v��-��l��KA C��^��-37,b�KI_L��]�W��2�%��Ō�v�d�vv��������B=A���v�"h� �xf[iFМ��]��,@�%§>gdM�}ҡ��X�tGw�#g��hj0�]5��l��kj�I�Ţ�1��y�����h�B�`8�ť,����K���N쬧��s"c`u��(��03���:�����/�1<NT�����~�4�t5W%�ۧ�}�E�9zs���7��|)�0i����Jngb�_���6���Rt�]�4ϔ��|'�~���(��b/���rG���6�4a�Ӟ�'�iF�(�t �����^�"��xv���6k�'�%Q���ފ��޽9��"�Xf)�NR��;�	���g�-�� ]�,5̀�&��6;S�+�)�y�ܺ��i���,9�ߏ�v���*�j&�E[�_��[�id�k
_��)��T�S0�7?�"\�s4�n����s��m�o�t%"�p"Z�1�t%��e�>Ʌ� ��h�Vi�Җ���b�j�U#�e���J���,�(9���P�}��"T���lQ�z��E��������4�=}�������v�&2�kߏ)[��L6��!��<��|�WVS�f�-Qs��t�mH�q�/�ڶ3^W3�Ϻh�̣4�@�5_��OZ,�WT)n��q�6�>&�?*�i< �_j�[���ߙ5��VЋ��൬qꠤ�@�D4mx/�;Zd��g��8��g��Y���^S�Y?�(��e�Mڹ4٤-�g�g��يI�?���z��皕U���lm����W����LP�p,�{�>����e։��&e[D0�(������E��ϑ߉^�l��\�����Tצ��Od%�QH;o�
��i�NԘť<5/�R0j�����z{�4Zx=3�fQ �u|'�)��I>���=����{Q~���_.^8#{T���vA�H�[��Wzڋ�9e��B�n�p��z�R
�X(���T-j�!c�ex�� ��n�ݐ�\]�1�M2�� ��|�'���>��ƿm�!��iCS�7�s��u?���S8���A�/��E�6u2ʇ�s�ZX���m�hš���W�Q�G5n���J��r��v{啋���>S�]���9n�	B���N2R��%:�{��˩ۚ�L�C�Q^�k������	`��5���;���9g�f���U)s��Hj��>9��h08}�Hx8,����7L����[ؘ�v�^Yo��<;����J�ꖅ�U?\��xu:"�.Ls�/��m��-J�W`��9	jЫ<��|�(�A��\��������&k�f��j��j�,sRM�A��XMl+��^iphǃ�����N����ś����]^@�����~l,P��]�{������X�
9�,�(���@�xU���Җ��+?�b��Zjx)�Ҷ�ɝB@��e&��Ț���r#%��!�Ŧ(�y��ㇿ/���K�M��a)ۂ�^q�Q�#VVze��7��;U���W}�_o�k;��&ج�.i���$ۇL��C.0,F��6��w�@�E��*`S��d*�tl'����v�ʩ��DE
�p�B@�L�oE6�(�>�������!(0 �ͧ��\�Y⹇��t۰�V~����?�R�����0��֊ݝ�V����F�=��U� �[�M�sͥL���!��妗YQ�1��4�ɳ�δv�e�	XD5*�-j�^���IJ��m�Z�M>��q0o���0m�|��q�k�igتQ�>���"?i����]r	\S�%t����n��6���\!|������ŧ�����`�ln��'ڎm;���}�U͉S��yV��<�9�f�<t.e�O�5m�LΧCefW>�w����&�H�"�v���
X3�,b�03���J�n�"�SX/r�uۇ��b���R�+>��`d�Y2Q����.D�`/��������+��x��;K��,��u��w��޻]�A���ܫ���-2�a�p��=�����j+�vn�N4���#�B�����Љ>3�_��9���=c��
�=��%: �(�+�T@��m���C~OM��E�lw�-��kB���q�N�癙�TP�w�#Jfo��������������<��>�*(mY�X0�w��m�7ƍl��6�Q�_��<�1k�[t<<� _8Q�	a����.#(`�,jz�K�j߻�xgb�U��	��YE�Gu&��QϘB*2}
&'N2,��
��#���
T�B�.
]�*��Q��1��S��~�{��ez��B.l/%R�kʊ�ET���b۝h1�Z}p~��Э�쵼�}��f�s�����M�$x~����Ѣ�m&H�]p7N5�'O7ۣ����[��k>��ϵ���| \��=6��x��V���Xi�<��$66P�q�P"N����3�{�
�ź��l��`'�� IW�RX�9���k��e��A�Tf��o���ϥ�'���Ԗ��0s��6��ŏc�1���񿌜?��~��T�a�i�>��n��{p�w~k\�z��fY�9|�ӓݖ�'.�6P��qX���2��}m)pMiL�����z���m�D�aJ��d*���믟�.�`��&U�e�d:J���aS4��ך�]a;&&��|��3,C�&�'��?���/E�a������l�����Ye>� �F�w�£��o�Fi�y�9gx��XG��h�;c4ǳ=�Y�5�}̣���<Ӝ���f������|��vY�G���k����<�-��ۅ���͕ts~�b���{��8�΢a�x��#�wߗ��Z��@�0ο����h��O�Q����UĘ����}�X5����$+d���2������ȗ*f�����t�97�'�!��[��N�;0��^(��s�1��1�L~��~m��5�����/x��_��_�.|o��Tx��	��w(�A.���XC���:����$�7 �Iz�t�R�m���fj��n��mM����*���vyQ���(�/�R��~��`wh�ߩJa:����#�!9��� 08���9�( �+Ì8a�hv೓���A@�L��炥���h#��>����	R�fҊ��x�ϳe�	߻ןU��M��`� Y_�Ew�B�h�h�qeԎI�]�Ϸm�Ex�9��;����~�X�&�/-/��yT�4W�n5""�'�����>����~\�ܱ}�U�K�PD?#���'~�B9�w���uP��)���.�C�]6~jc���F�}���@Q�����f��1i�E�r'�e��|�3�Yd�;����ۿ���w�/�����R_�
6�Q��� y�<�AQ�S��]�R�����q-�sG�]I��+��3�	l������U$��oM
2��ЎRhhc���F�S:�� ��R�w����=�!�(�e�e��e�P�Iv%��%�禭++Q�7���P6h�E��̕i�Y�U��Z��2��6hW��z�3�'×�3ĉ��]sU���'�5�|Xkm[��^iE�U����볛줟v������jy�-kZ����Ҿ�a1b<W[�^8-�w`E�h��t>��4U�4�i6s.��N��hU��ڝN;�N!�b������W'sn�OĶ��&�;��ֺ���3"@���}��1���d$��Hǝ���h~q~z_��fJ�6#Tv��H�3��#O[n[�>̰���ꇚ��E��Uk̼�J� )&2���k�����!|Q�0=`�0�	"�2���_�I��P�.yL�<2�q�m��O鑌b�8�hXz�N����.���ҟ8i'כ>߰��J�ƈ05�o���$��L�a	^[��V���7�9�(o��֬�֊ѡ]^�Ai'�N�R�BL���s����"�ü�ͻw��-z�}7���X?�A��&�Ź�%��g47�tS�� &���1̽Պ]8�؇i��|�L��ҾX����eqWO6����9���
��z�)�^�$�r���s��PG� _lS\��VɬF%Cw1�/��y�<k����x�.�K{�I��Ьg�eJ�O
�����c43�tǉ�@Л��p,C�G�yI�W���N�a˞8��Rk�j��o����kMo@��N9��|�R
�Y<Q/�)h��Z�5�ݳ�"_��˜�ۜ'���e���_��c��� bh��ԴhLp�y�F���%K�*�5A�#�Y=��w@���	�ֶi騿���J8��r����)��N�C�U���i��A�a�����a�bl�f�m������l���`L�搮����Yh �LM�PD����:��eֽ�����i���f֯{df9h��[e��qZ��>�Zi�ޤ��j:����M����iX5ū5u�y쬿��,�t��� ��E/zQ�z	���# eK���ۈ�S����V�7��SKT �N��W����	���m��6ڝ�{mD�x�4U/8�g���C��ԙ75z� ^�4�{U�/�t�0�N�����jd�Up�Z�}���,4=��௙d����H��5tI�x��X}�.ҽ&�����V�)O�����D�p��¼ԗh�3�r~����y��^�ۼEt���K�*H�-5�8�)�&M	_�5_Ӽ��/-�  b^D��	�_����#������n��פ?'�(iZ��Fo�=�Ӗ{��c����	��1.�	Qgޘ.;�Q����ˈ�!�9Z����f����P�e4O��b�Y���N�E(��e�E��^`�۾���wfo�%�gԢ��T�����7,/2��ʫ!ss�����lM�d�]d��Z4��T�zQ��w�~�Z�C�JS�֏��-�B����w��(ur��~���9S��h�ܹP�����g��&�ű<L�+�}���s7����(-3�߆�X�^��f���?�8�D�؀�|��ߘ#>��UE�'g�X������y��"J�j}�A�<�;o�^��R#�"�g&�C��{�S�ؤ05[n����1KfX�p�����^��V����������fH�ۨ���K�,1�O�� ϲ)׿մ/Mf����z�����"��:l�K�/1�8�	�\��FL�<�D��g����6�/J�Ub��Od�>ZieоW��!j[#�sDz�w� �{P���}u���N�'RP�@)<�	OxBY�f�5�H�
Z,Ę��؂Q-�jA�`�+���v�SK����M��,;aݧyݬv������f\%m�B[��vnvz�6��IXk��m��ˠ�v|G؁����Aqᵂ�x��乊�btI��y�z�f�f�2�s�WW�ټs�^��j��"g�aH�W�V�ٝ�цMK�j��Y�7?ב^�-A_��P;X_/��hF��[��k�hgP�K]����n��������N�ґ����<xE?�яN�T���h��l v�uQY�}��t�����p��k���.2o� �>�'>��0YM���MR=i�Y��@0"ǳ �����$b��}�q��CaWs��ZG۹^��ELX&NТ崇�w���������4=ܭ3������I2�,�h֦��JU��n=��K������,B����nF�ԞX/μ��|s)Q-h�����^�ѵ�^;�D˰Ay��C�E����HL�ٝ!�y�i�R ��[��LQ�ݐ�=$V�v��;"H�'Z(�Ȑ��t�{lF8��7��M���}�ו�A��[��ɟ��TF�j�L�x5S�
]�ߝ�Y���`YQmy5ҬA��"��m_���<ٮ<��q��k�d3ȇ�F�j���|utD��f�H��2��!� S:�2�54�/"S�3�;�b�
�4�X��A�ٸ�����r-�d�Qf%���j2EڊP�Ǆ�/h/��xle,Rz�y7>۾6������2,}ɤ�=��Q]����λJ�Й��������R:mP��JɐM"ن�D1F�8���x` o�dʵ-/�E>W�n?���<ِ�����U^Ÿ�Y���"���k����M�y�{
����y��)r2[sY�h�\��0��3��̴�+�%1�+��υެIgh����xf��E�u�����2��H) $m�ޟ��N]ն_HЗ�X����3( �e�����j�S@%��]]�(+�)���+2��+M>H2]�\|�������䋿��(G�xP(�Zv���(p���I]�9 ��5r G+�Y�r7[&�s����X��s]�|��y�4���l{d�=���n}�G��eә�w˜.E��Z�{w��8q� tn�m��z���N��7�����Qn�4��(�jd�����V��O�������wi��t�V�V�B���|+�g55���u(HL1���� \��1V�Ԅh�*yV��!�3Y["͌������z�)/إb	��h��}�@�� ���y�\uQ}�D��!�.�q�K�Ej3i2��)��W�H�5���T@)� �m�D�(�G[M����N��_��_++*�"H� k�9�yN�Mj���R͟g���Y����Ⓕ�tY�&pPUwl{�^�k��.��R�rR��<�h��dz�5�p���_�+�n=�]���¤��2<�2�^,'Ka����8�����]dW6�;eLh\Vxe|͉íe�r�������M�Hr�X�9��7x������-:͚�FiG�R4�9e��B�ڿ��碑%S}>�Mm�9#R��ѥ�ڛ���"�5�P��ڃ %�־2?WP.H�P�P�Unh�Ȩ�Lh�����G���##��X��j�LS�A�DW�0�Z��&U�\� V>�T���&��*`�O��OM;S��E g�@D���m��Y��L&�h�{�*��".�q�r��$�x�h)LHg��c�J�QSH:I�N.�9�]h{��Y��[��!@���9�i���}�k]�jd|pE��q���cĿ3�)��z�_x�QmW;�+�Π�#��X�{���1�P�k֡�"��p�:s̶["��t5{h*��꼁rA�9D�]���	��^����������� P[��L���vhb��n��g�1���[�ȹ�};�~�GG,�'�������1v���f��Pm�H�,�a�h��a����ud�h��1g�2I��b���� ��i���\]s���Y�G���+�ղ�}:gr��{:F]XH(H�
�<�����a_om�0���ń��.D�����N�s4A�͸�Ψ��Y)���NwS.qÍN`�ž��#�7�C$/U��1�Ij�R�Q�m*D)e��X���s�\�e���^���ҧ /��9�����b߅�g�,�Bʸr�����e1b�	J��T#��o�ʚ	�j9������ZDN�;�>M��Gp��ϊs枳�����!'u2\��$(䤭O(��iO{ZA��z���+��+eP�v�����"��,]�=;�P��D�P)�Dz����<GT�0�ڳ��(;M	N��;�6gU,��ue�e��_
���{��p~���Z|�GeM�h�����[�IGc�:�.�}څ}�Ef��˽
���/e�ܔ��r�M;����B�6��p�N�.�s-CN�Ye{�.��{��N�E�<��gKg|���[%��p��/������r�Y���H$#"DЖ��<��!yuTJ��4�j���R�M�x�����4L롧�*Q�<���D߭˩
��4C;\]DPt\����o
9��5�)�'���Q,ЬP��j��^D�z��hK�p4�v-��
�I�v��L�k���Q;B��H���P��
�,l�ئF�t�jt�n�����-���&��m���λ2�<2�t��h��>z&5��?�-�A���d�	�V�����p�Slė2�����^�M>5N�hj��0�\�S8v	QH�r>A�O��(��U(�춋߻ڂ%����8��TL�:|F;��>�k��v>EE�ڴ���9� ��s��B�y��_�d����V%Ul/͸�֢sk��O5�U<U�o{�ۊ�Fx;6=�ڗ��t��b��	�����g���:���~I���T��ez�#QWmk��� �h�n�����=�jh��`l<�d�L�kT�.x�q�[���k������@a-�^�p8�y��F��C�u,뱆R t
�м�R�L�ؕ�=�G�]>��8�H�D��x�͋_���)OyJq�s?�I�"��L:�dSon���<LԿ������s�S[8u@�fd����P"Vn�=�F����Fꕖ�~��)�)[���
_h?��yt���4N�m���w&;p7:�,ҥ,όZ����[�����y Ӽ���E�%�XcзU��ַ�=X���B@S_BP!�U�.k�祶�5 ��4y֣������R�ⶻok>��6w������Ul>�'٬�Ϫ�:�h�����I5�T�ۢ�v9��J��$����E�y�7)��w���σ}�t5J�t�u����O� �2���1�"{��V�yx�m�]4��}i��j�Ӷ�誨IS'*�*1�S(���^�2J�b~.��Y��B\M��y�Zi��4£�e��Y����2�Nc��[�~6��vK�ܼ�&�M��_p�K�q9�aA�<��z]A�~�|
[Mځ1I�����S����e�i�ά`���#��hsí�R�l�����D8����T���p�ݦ�Xt��6v�N �ź���ric,���܅�b�OA�^�+��f�ʌ���[o4�s�pυ�.�t,�5^|-q�r��dw�@�Z���!�4h##������y������<� ϸ���7*��iW��v��}���-��<��YIw��������OpW�e�?,]�4)�>�É����5��񽴷�����l�w����d��y�(��D���0��Q[v���0��cȘk��m���a��/'�?Zj�Xf�Q���X?Lx0KlV��A���Mx4)��Oa8�3�F��E,8�i�o���qͯ��U�ƌU��+
�Ġ�@9bA۠��ݬ���e�_:�2���zj�I��7��w���dS�f����]F��r�ڬ�+�n�E+Ee�V]Z�;�����-ȳ��kHa�M9ߧ��Aa|�tX��7��㘳��ڂ35�cY��ΰ>� �L��GQ�0��u�	K�LQ�暃N��)�ks��ze:m쾬��ԟ\�ܹ#�,cc?!��(6b=ތ	������'��~�p����3��#��a�'�2S���2� ʪ���'�����[D�c�"[^#�-b5��a͸�	#�<��7M8˦��	SE�Wb�.�8 ����/~�#�����N�$�R�	 �;�9䠂q�����A:
JA��m��2�明<K�@"E�נ�eg�Y�59�FK�#.'��z��)#Q"�6�E��2�3ge���A��I�>�@��d�Q��F³4;�`���s�w\����1��e:�h� �}�0�=Z
s�tJ֛H�|�s҃t_P��*!@��=�n�iɐZ��Y��g8��i�.{!��D�ڈ�,6ߥԤY8�����R����Z$�����dĒ����^��xt�s�q9�"a8�zT�.C�VĂ��fM��`�ti�|�++�e�4=d�nskqw��A��Lz����.{$�l�3��(���YK�e�N]�X�=��=H� ��-k��)3T�4�oC�F mpt��� �G���W����]֮XF2��8m�҃t�R]WSD�,�G��eM�4A̪i�`��^��0dQlw� �(�y�Ö���j5~�#�K��N�3�򸖉%x��u7ǝw
O�@O��-�Q1�1�n��*b�Z�Z,��?큦�&:�Tt%vͦ&+�s���O�B�X���7E��	kvXa�ο�[.����g=�\볟�ly���}��ԧ�xn§���չ��Zͼ~��G���_��e�6�~��X�Q'+�j}A����ig��ǔ�F�pj���Ju2�	[1�0�e]����u���S@]A�߅��~���wwW�L�L��N��v��`K��
���3
����������˱0E���暹����~��C�^L�����^َ�Ҝ#c~��/��	QGR�H���]OO'�&]����~i/�X��)�ԏ|�#�lN8ⴟ���6Ox���}�c�w~s�F������2&��{�W���r_V6d�~�~�,z*�]�X�RO��E���GuD@�-vM4�Lهf�AY;���4#~��`,��a����yO���l/�.6|����y�K_zA�^H��w��쀮V�M��Me�,��q�-6�u�u��L1���C<:�I��")�f 	1��l�����&�Գ�W�Y<\�Gx���!L�!��gU~h�������w�5KU��qYr�@(���-8��)w�6�ߝ�3��c���*Z���,��g��1���?��JSR]�oY�.�ܭ7�??/"3��_7��><�a�5��nj����<7�����٘<�n-��b��\lsOC��eȚg���u��a�������i�^���ovmI�0*C��=���뻦��D�	  ��8��H$��=*r?����]�2!�dr��
=�e��d`�8N
�Da�f���@��x+jy}���+�Nn��/����_�����Yί$c�	'��.�ۏ��$"�V0��\Y�hrh�ews�r�pr��Yu�_}��g?{�N���N�c*J�T����+['���~�Y�A`$�U[��� wa�w�Ff�~��8��b�
(�͢e��V��q8�D��s?�Ð��>5:$N����~N��W�m�|ge=?���^J����C�9����sKV���r3�.�F"}�e�p����	z���wP�{�s]l�hkɷ���P�U�Ml���]��1���D�����`��,b���P�P��-����?��He����-������� ew
8(��JN�܄�3��}��Y^�.H���18�D��#%���z��D�j	)DT�sgm�:n�Fѹ�0��6z>�0�dͣY}4K��f�Ft	�d|<^j�ٮ�C~ss^(5�	G����l����D���D�:��oc��un^+�v��[d�耓���2�L�JS���c-]{g��9T�at��ǧ�`2!�q�bR}��xGE6��N[0�0�Cާ����� Ƴ�Șŏ������|���k�A�v�5�R��9�g�g�3������|ڥc��>�f���O���J��K� �3�Ф �G<��g����~y������s�|����s Pu��ϴ�g���s_Y�v�絉ľR�+�E��F�h�j�-��OԶ�h3��^��q|VD�����s��ۜ�v����{,�Q�1���p����&,RϫW\d΅�E^�d���;��LD*L}򓟜��yԤ�K`1�;����z�.!Z��mևN{���	C "PR��!Pm_��W�sElLZ"@wD8�������"-=����W
�T�^� �DB�ig�G��ɾ�Mܗ��?��?�jg�+�Ȫd�k�����;���R�3�#�+���s�M<�O��2%�c��3f�A�"���[�G�Q���f~�nL�ᗾ���f�����h�pck4?ad⛕f�4���V��±ߞ3��KkG�o��x߰��h&;4􇹡�{뎏N�=�sVBp�"Wk�뮛2h���e3�*C��V����t�pkC21�a��z]�r�Z������Y�&K:��	�E�$t�-�w��%��g�4!dZ���6B�2?��?X���C�6M�lV�cr���?��?l���7��G����YD�=�=9��p�'=�I�����s�."Q���o>m��2�|��6R�xj��4��~��ӟ���ܐX53B4q�9:�k^�{���d����VB��dK������*��3�)Z�&�vv�K�0G.t�~^u�aj�ӄݖmͧ;"��+�&4
�f�����q��^�"������+8e�D�V����Hr?<&2��C�MU��J��Q_;횵�Lov���I�9G�� v�/b|��V��ޞ��t��6����
=�^���1��z�0��8`���3M��D"8�ːp�gد�_;�Db����өC�E�w����ɟ,h�6s���H�tJf	J�r�]�j���U;K�gJ>�\�w�jG���(�:�Mb)Fnm3i\iZ�MEq+x�F�oƂ����u��|��R��C����=�Π�*���_U�z���j!�9�"a�y��;0�,A9w��x]�Ʋ{�Tx�|f�i�4�B��n���&��ϴ��c�� �ڎS����и��+
ә7c7�CS-���&���h$�h�UՇ�8���Y6��]��[��NmNgf�ʛ��ߜW��g	��P�	߳�9:�ϋ�!�	�~�}�N��p�}�!P��ឳ�!d��9�<���u2���
M�sʕhmV�LI�W�0��=o� �����<T� h@���f���:B2p��`QbrY�6�Q�i�L�,�I_�r{�e�i)HLڊ53d���g�`���r���§�6y�g�������l�;�<��7������ʃ5�p�#�򾦨�M�}.�5_�}s���t($� �Q��v��W�:���2Hw8����>lrw�r���� �������nj��,A��9�\���Q��ʛ%���.�!�������jXm���ѿ�g��o����x9l��`9���:�>�Ut��G�gݍ��{N��B�{�Y���i.��I;n�B�Tq_]��}�B�b��3u�^�1�Ye�� �\S;�o��1�����Jm�>��}p�f���N`ϟB.c����p�ĩ��#8���ۮX�G��_��E�m��0���Ɵ'N���:El�z��C�[�Wځ���������O�o6��@H�
(��#���^��gQ
�d�4C̚��T#s���F3��,L��U֪?����xS0�M�߬�����57�!f<�QR��]���&���|� �@�X0��(���-.�i�2t�"K���Zf�5������E?��,�̉y�y��xl�.:(�Nw���vk��lU�MlX��c���5�=(��{?�o�3�><�.`��x`,�/���åJW�g0�H�K�Q`��[����x�rY%+�O�i��N�ɬ����s-��~��2J4m4��`GmT@&�M�B�&�	�̊�j�p1�q��fۛ��\��!�+�k��7��}Ώ��E��������?��D�T�Jy���W6����y �v�)�3��1�:��@�_5�4�0�,X����J�����(�r9
�Y�9☣#���(Q��nc����u�f���$���Ex�&��oW-|j�ϴUVz�?��&4�I57S}s�s��~��e"�ݿ�w2�5g{2 >C�2LG�Fĵ��ZLG�舮j�D��h~�F������ʢ`C ���O�8y.���^N4eg��Z�ǋv��s�S�h?�<J�-��<��գ���?���������FG(|�9���Q���-K)�چY��5A�)B��gj��>Ke2�Dg ���K^��/3�Ĩi�)myQ'"lGC�	�"���U����F�������Yk%iq���-�poT�-�r���������=G�f|h���8�d�X`l^��;�SJ��=7=���f��ZAo�ۋ�&��	��-T�^�{Eo����/=�
*l�L�.{�#p� ߯��B2<�'|*�ʈ�&�Z������o.P��Ԝ�����e�b0N�������O���t�!h�P�i���<�'ٿ��d�x�[���t�ME b>��k�����k^���6�Z�֋�NJy�y@FZ�}����T�1��L�X(k�A�_�ѧ�7���T����˄�t@�2�|�䳎tqBԦBvT�cy���٪� �^�R0#����� �ڼ�v`OA1��>���
C:og06?�W�5~�}�v��?���bC����N�-�$�����P:�r¨T�m�p��۾��u�ٜ�F��o,�h�(�XC��y2����V$l�En�äE��2�H��C�d5�ְ*kB���>�<J3�Q�}`yO�^�	���-��@�@���f����@\s� �T匚�|4�v.�y�.�4M[9����7�&��O��V۝ʱ���s�����#�A �!ad�=Z-6�V5;�z�[� ��I������pТޖ����j����V���V�A�c#p�fפq]�`bׅ��i�Ө�=+M
�����h��*��I��@��G�o��h&���� kRNM@������M�]ǂ�W�����i��N2�j�Ь�DTƣZx��07�
c���|hz���}��i���f����]��a�ɲ8g�	G���?��X^�A���w|�\B�R�m�s��yF��3���:W������3�Z���w  ���,��u�ˌIx����#�mv�X���j��;=�\r�
���b�f�����l�����6����VVWoﭮ���6ۡ���������p������m��j��+��S뽕��5���i�;;��#�7 `�A2��	�l2���5&�G�T_p���*�I
��x�_}\�cQQ��X�t�+���ɿsҙ��9 :P��j�E�u�tMYD����O|b�7�aϹN^�Wۍk[�~��㢌 A00��ء�i|;�n���	������_�*~��#�_d��\� 7�P����r�"�f�X��v1R�b6�Y[3W����Dۘ��&5P�
f}]�އ�%��9��bѝ�H�`^�"��k�g��m�k'��ub����S:<q��m��S_X;ٿc��~��Be{pb�3ē����G�Νy����Sw67?�<zg�������U�Q���';E��q`Pj;Q�l)���t]A1KT����S���*t��,�嗿��͓����0|�[�ZTP.�T�W��_J��I&���,2�yf�!ϯ���'��֎Ό�p1L4g�jީ�6ե��%��Ї�Ї
o��u�+� t��c������O�g�9E�:K�G{Ws�}���'���?}"��'��yâN^��m���  G�\��d�A�ӋBY��P�m=6�����@x�I�Y���w������^�������m���W=䃽S��sW��~����}��Woͺ��7�w��ӟ�X���U���Ǐ���g�~v�̝�\��~�a�!�ع��g�_��Q�dK��yلt�#DE�:�p�Y4H{h�MoFmReco.���;<ݿ�˿\�b��>�,�js����p��F�^R��tX^"�e����?۔��*o�ڋ�~�2��~����0}I\�/��/�=E��vJ��K4~�߂��|�0��
Jx7��E�6��p�s���31Ͼ�[��h� b��)��
��=�s'�o��oO�AF�dx�qҡf1afTI�o��!����k[�'O~~p�C>�y�U�>����g7��I7��|F�י����������?_������o�>�՝�����>��1��Xg�G]�&�A�ƫ��1�9�����_}��W��`l����jm.�����8���>�,�(��o3Ѳ�/�2����p���z�긓>���x�R���ߘ�@r� �qcƯ��l���4f��� �g]5�״�BڬYl�M!���E�"�se֣ a����0��PW�Im��� ��"��	��`Yσ8�<Nx�<�茘Ҟ���<-C�O4�VV7�n���֕y��UyO�a���O���es@������z�?񾇝�����'���yp��ן}�7��5ɬ+�dҍ+�MPڴ�İ��F+Ӻ0�[Y��U���:����Jʤ�;���
�Y�9�<8XP�x�ɬ�ʻ�L8�u/�^���$����\}C��&�B���{�)��Vp���l�"{�bV`)���ؤ&/���3��50�]_d�K��e�R�y�o�PTô��8����!g�S�z�э�ŝPCR�+�^XD��1�e����>���2��S�G�	���˦�&G�.K��y���P[��h�����8��s��݃��������}��s����?�����So��/6���hV������+7��*4h���v5�W���_�����f=,��$ʢ�g�����ZA��ŋ1�:��Q��D�:��^&m$��«�C���6���Ѱ[!L�v�N��2R𤗹F���Y!j�'_���8��Ƣk{l�7Qp-��]��y����1HMH�X��6�d��BH�b%������)�B��O��O�1�
J'S�^)�f����q|�jkj3�A��f�5zh?!`�ۍ �������<K�]����C�e6`nQ ��^.�z�<c��9�6:"i4���������t�ݜ�m�������_y���C?��׿��8�������/~�CkW>���F�ίYkzW�{L�Qz;�����~��8Iz��W�cw���ʇ4ḁ��l'[����؛`2P,�N�y�BF#��UY'�s��ܢz"��&�\��
�+��d.��ȝlf��f	���RsrմL��2��3/{>��
%��k�~��R�ÏV���L����/�2 �dLX�+^���~�Ǧ��2痾���ق�O_�QD�=��y�5Ρ��,��c΢��B�9��w�wO��C.�5�����/�����i�maԻ��	���l������s-�:u⏆W�~���'��/nx���1�-?��}�i�����`�����\��5�vm�[/��j�;�bP�K,�����|Q�e�7n1L�BH�Gm�fM��h�+91����w�|�+���+���#g��.θ��L�]"��Х.d�Ѭ����P-������\HDU�%�	K�"��^\􋠂� 8ٺԾP�����7�\�ז�(��HQkk�ׄ�y���β��"a�-����x�k^S�jS�AHsJ�f@栵34��X���Q��Gl.���j�_Yk�������[}�G�u������1�����������7���w�����7�|F�>ͥCc9ܯ&�pƼZm;��xFab:�TH�1kJ��^W	[�{v6ÄX�l�|�:"s� ʁ	ͱ�`�~��KFcEO[�ahV�X~���c���}�s*���lbR�Ǽkxy��	� ��Ř�)a&~�@��)'��3Q">����j��BV�<@˃�A�%��>�N�����%�A�_���xz5D��i7f2i������훠�᱙#�Q��0Zoz�'ϵ�����?������>��+��k����:�I+۫덆'��z�qt�Q�+��F�J֞� �|�b	�1Y��v�%]�|9k������N�L`������L{��f��]:K4��%P갠K�RŮ�(tXD��<s-�<A���sSP��=Hm��P/Y����wY�s��� m2>�!�KPt�9�O�������p���f��F�)Q�O��@^KM�P66���_���1�>�~�0�ߏ��Go-�-�ڇ��F<�/����=�~ss��7���'����GW��9�[��~�~e�k�hX�hkL� յpxY=M䒔�c t�������EH'w�5��
��|
g�.*�Ӗ�m���1�����.aH�h��P����&lȖ5��:�vQ�)L��&<���}Qɩ����6�%@�
�.��������9>��@����m�s�B����z"�Ed��@ �`$�>,�98��>ۇ��h%�$�����տ�Վ��3X?�?6O�x�'������>��kk�>}�7�����`篍��2
+X�{��E{J��1q6YMlĮ=o+�&ֶ�M���%9X
\���SebtCdtr-�I2�L]�EyH��ѱ�%��`wCxX0x.P�QT����R���j�zm�?�Y%���+�.�c�V,ͺ�ـ���O�I�L� R����wO�]��귄���h��)�G�`d��،E�HF�:7Zլ���|��˽<f�7,2����}��U4e����Y�F�n����룍Sw�_����ɵ?k�c���_���'�|���A���͠z�'���kE��}�c�⢎i }� ����sY��\�A�;�
VO��vf�>�/�o�����ȝ!pȩ*v���\��Q�}XA</�������2+�������&������"�1%���a��ʐ.$D�5Gl�'�$�߬{��?&�5�a�8�ۺ
A`E3�&!��I�hl��qaX��25�,�!�b�@x��n;�����`XP01^�G��&t�q�c���� ������\u��'�z�؂��7���a}�����m��k�VUMV��N769�C$���K���-T���:Hǂ81�����b���$�)�c�Q�Ҹ��yWgse�a�ߨ�˖1u��lzk���IO�hٰ�>�$Fp{\?�2�5�@�'Nxۤ����!?NJ�������ctpZ�ŅqY���^��F0�k8�ue�H�X��E��'�s1,cK袻m��rA�]D����������_�k��5�3]Y7��a�f��7h@�]�ɺ�j���?������X�MVȲx"��{��8������Bxp�Lo��.�������k����$e��++��N�E��~oog��a�h0��������V ����1eƆ�X�(D�M[��ݔS-�z7[B�s3�;2�B��Y���jS���߳��]��\ՙ��q h�:�U;v5Na�=�+�<�XQ���gϻT���?�JAg�%��u��l4H��E�3^,���-��@ծJ;�����,���R܉�Y�0� )���h<n��ŋD�P:ʠ�B��VމYw�E���pXPh'Z  �hX���C�7{�:�4"�D� X���w�I����I��^�J�������-�l�ߺu����DgO��w�ε�{��{)]��:��	1��`�"��&Ӹ����)@a>L
xuq,�P��}3�����L�aT�5�!�,���.����H��:׈̐&"�ﮓ:��tI���sml�81��=�=��y�ѥ �]XV>+�8�9r1�8XȌ�YV���׾p6��q�Oe���-�9��|D'���G>򑢲c�!˫�[A�+���H[Ԋ�%����E��FD<^�f���C�-`Ig�<^��M���nIu�<����\�?4��W�7����^�k.�nN�������B�e�$S�����%h۽1v�3X�����3 Z<��Lm}���3S�r��tҩ���`�d���U�d����@�.��䟌Օ�k>�o*��%�f����T2�jDs)�Y�M�x��������3ĩZW`�"�w�g
/� 3�Q�[�����E`cG~ӛ�T�0�������8�>�M�k�4���j.�>�s��\҃y������C�����u�ڡ�f�����Ͳ��C�{2wj'�QDAkG���W�K��Ѯ��;m�Μ���x�7�AU
�*Lt�9b���d�����ΰ (�h���  �3�|��nGt�(��1�Đ�b��,�D�n�.Ѽ��i�E�h�캚�!9FX��\���\��k���)�J�J)�ٯ<��3jf���������N;���#2US��A��A�8;3B��R��{�w��r���cN^�9�ݐ4CE�.X.4���_�Q
�@�w�K{��q_�s�>H��:s�r�>����oIZB'}���]�Z��8o�oj�mtP^����6gϟk�7w��u��n���X�q!WhQ�L�<�o��Ewjǈ��w��3%�8��f��	nXS^6������4mc��ն��K���ڜD����J��մ��E��T�Q�=��nl�p��U��1�Y��EW��w^�WcsQ,�����k�(��.�FZ��h	(Ζ,Ma\/j�0�9#E���]n���U)����0�n%Ys�*0���67�5����Q��.vd�?�wv'�`�[K��Ɖ�ϱQgF(�\�Ex2�B��PX�nD�N�L<Q���N���zO/z�	���qMuZ�bׂ�5�3��U�\�ḿ�lӌq)�$jS�@��*3~T!�y�ť��86
�T�6@`q=�-�s!y����F�i�{-{�qHZ~Ja�(�d\\d2�85A�a�^�v�<94�qmHm�y�}LܨX�;}<s]��vv���/e�;� �V;�KK��8��Op)�n�C��B2İ�ӻ��n_��t�Wl�ﾲ]OW}��h��zŚ��u�9yb\����얦��k���6�O����Y�r�2�,y��X�tR>�Ne�I�3M��5�)@Rșƪ�
bJ��bemUX�>�̉���&����'�Œ1�
)��M6A�]�KCyF���(o�;�S�)L�\8���9j�>1d�J���|�}��rGp�s��!�O�N?F��8�|��WM=���!&��7�����"�;�`�~��߅�-��Rk�2I|hW��N�-K5�щ���ک՝��lJ!��}u�l�b��=o�����iVڱ�z��f�?.a9n7�_h�����y�U�ze���kǵ%B͑���~��D
�Q��r3BU.��W�WK:�ꠅ��頼_M5�f��~��|�Y�����ɘ0�uT<�H8mԗ2�N��3����i����C�{�!f)D�Eϩ~f�L��-o{�ۚ�����X򥱻����L��@�E�<pw�)of?)�r;yy-#0܆`f?��8=���:��ej�fa��h$�
ND�vk�Ȥ�Y�&ΏI�(uo9��N�ܐ1���՝�W�v6�����W}�E��}L�;mek�-nX'U�K_�vƥ�餭���1�	��i����|3l�J�vONd�	��L[����)%ӊ:-��w�I�'[U�+��Y"0e�E�:Lތ���)��>�L�^tE�])�:�uĀ�a3hG�8�$`{��ҟ�fι!���󬝒�D���~5H�l,zj^�gTK���"&�s׵�Y��t��4��?5O���Y�n۴�-+eN^��n�������9������P<���7޸2��?bo�����G�b8��XN�Tk�V+�W��ca<)�Xl`-���L�� �T�e�E6[3������L�a�rɕ�Fl���TSiY|kR�	�ʐ5ⵄ⥎��t�9!y��+��LB��/��4e9~VJ#L��<��$�m�1m����?���~�2�NH���z}ۇ�i�S"���t��Z�,���0��d�q�K��~����9�1�_γ@�7��	�T_�.�M���y�c�C��o϶�̭O��x�Sox�g�n��G��[n{�`�oX��z��p��S �v��={g0*q#'Z����l6'N��
K:[���n���&		&�� ��E,��'g�&�B�(�(��oJ�0Y��qN��6[���ښ��7(٢.��3.)���:4���������^"�4}1$< ��A#���Fiy����B�*�3�7#���1P�1�����W_����d�l�u�!A�fO���:�Ut-�ʵ��_}�u��a(�Qɳ9ޔpg�:V�(hA/�:n�Ȋc�z�L��k��Z���湝ǯ�{�3������o?��t�����k[i�5+��IWK{�������q����x[txr�9��hΞۜ&R����|`�	�gr�s�A|�63�3@���|O��QM�U�Yq���t���`ڃ���q�v����Xe.�
$���}�R%�!ǖ�s\ja�3[����a��?�X�чSM�EC�|='ۚ��4w�	2"Pڥ=^���w��S�UѪ܍E��-}������ c(�ǟ�n�s��/#���ģ^q�"vX�E,�cBA���KKZ�K��^��8�4�L���7��S����{�I��g����n�����ǭ=�Qͭ�]��u�	+Ý+Vʆ�Â�K�{ㆮ��0��j�`�!���:�ew��1��wu��g�&���2�67�p<dc��Y���r�6+����</�-���٢{��D���y�g���R� ү�ў�����1���@�2ce�~A�6\ZO�Y%b�����{ɧ.�6X��s���cjU9?D�"�j�P+�gN���A$��G�8�wT~�\��Txjrr���>�*j��'{�������Qq�x/K8�joxf��;�y����x{ȁ���D7޸r��_����OY�����!��m����R-Z��C���v�J��F���V�����g>5a�a����0�^��WM�����R.7�j9����ľT�&��ZV�ʭnCi�K��3�A�@��0���,�d�/��,��Җ�,��)��Dڼ3\K�flo��B�q *�%���X�y^�6�ϐ*��M���وP�
CFBh�b7g�0��n��E�Ĝ܇ҕ��sσI�~ꧦ��9A�u&�9/2[�=�m����<ƉyTk
a��}'ьs�����rG��h6Z9vb��Ki� ��Qg8h6Z49��z��]�|ss��w>����^ks�
�}⎧������{�z����ںN�I4�8ך���Ѷg�}��hՉ�v�yc!Dm����)�Rq�\}3��>�^�Bȩ��(Ԋ56��`&���ht�Π���&`V��v>m��q- D��/�lE��_L�h��?j;fF)ty�DN^���A���O��6�'��6��ΩN���H�
��d�M�cY(E�)K����v$1�!\��S ɬQ�T�KH�����nsDQ{�0�uY�uu)`�&�v1�0&V6tN��c�X�O�*��Ѱ���ޠ���������i;u�
�a����gn���S�������7��?>���Z|ݟ~�/����/����x����+(K�&��+po�LG���]��v��y�7壘�D6�3�©�����Pb5k��P*�#/��mͲ���|�̧J)��ȳRHUJ�q��j;�1�-C�,C�	��6�@��E����h��{�Yז��ꈊzLs��̞T���3�*I�1Ρ���uf��c��9W�N����]�]���z׻�Ü���ٮ\�R����	�r�1��t�M�(�u��i�����4j������[]+[����Q;N����͗��h�;9>l��۞������������w����O5G@W��3'N����in��[7��E�v�>����:��~ �����}�mF�gt�T��.�<�Χ?��� TO:�dl(F]T�ļ٤k���0��&`��L~��ɉ�3&��E$'oz��=���p.��E�BB�f9&GL,�:*C�xT&��M��qн��on^��וJr�%���X2Ь?�׹�V���o"<#�����|Ԙ��Z�?�ݖ{���aoeg�26�kK�o�� ���ŃV�g�;E4���#���z�+v��!?�Ʒ�x���=D��k~�M������o���7����ۛW���ۓ@�X�܈�"vx������͸��|�T��F�ZO��R@�z�]�ݵ���|f	���11E�:���oR��!Q�IJ��	�|�/��5�����늶1�Y�1��yη�LEN�./Q�6����}���0��~N�0��-oi��ۿ�b��pNa��w��1�sc>!��(J�v:��6y���< ���
��;->?�vJ��x�L2ϲ1�p����J�P�w{p��w>{s{�����#����_{������������s��So�q�\󹫯��/Y��5w���[�~j�mQ{|����~��/���wƏiGU����Q��\1]���{�ʉb�if�V�J-"m�NLQ����N�����$���[Ln�M|���,^��j֤�oC�f	�㶩gy��\h�q��(�4 �%�[�N܃����#?�=���ȏ�HI�f_<l�V�s�K�dF�8�� �9����.��L��j���7鷝�س���6	�\�l�����R�E��e���(��IY�5��Xȭ�H���P���Z�w�k�޻}EsŽ�w�=����W���˝��w��_���w����o�f�8�~�n����qjcutzx���z���YW�u�3N�{���g�y�����~����vo��=��`���a��P� .	��������6ᬠ� -S�t�
+
ΐ��E�t��愫�&\n|(�y�Wz��&�	�S)��s쑊�&C!�4작���A@3��]��k�p.b���&RDș�,E;y�k����YD_�a��������[+��	�Bg�a:��o��X�|����Ú��,�T�ﶝ�{W#�Q����gvg=럍mV��b#C�#%Ĺ���-nV�H(\r@"6HH�K�,$�	�A � !���(��8��z�;?�U�{U�zjz{v����'��������W��{Մ�q��ѣ���EO��VU�*ݒ\<�[Q@X\۵+���0CceB�W�3$I��Fl�ɭ���R��^>*gO$���hddf�HrE�M.~�o��^�i[�Z�<���e�I����C�4;�,5�'���Q���PF���=�1.h�%�F������zh����XK"&t�@"/���m�_А��2�]Q}�MQGD�D���K/��E�W�ԡI���|$ȓ���(�>}:'�li	+l����Z#	�ॲ������Y,��PG�:]J��K�U�����}��j�zA�H��G����9�`�$�'P">t�P�lI��,(ݢ�IS�lH��Z�u%�S�oBu������ f=[ȹ�S�/|���$���ρ4�'��0f`�`R�TSHÅL�D�Jq����+6� A��D5����cB`�I�U+sY��(�y
ucB��\g�h$u� �WR��P?*�a�@�u��4;��9�� C$	3C��^;���`�Z%��P��,������/�B�Ӊ�}�a�t�~�!_��gb�'$�F3>DqUg��_��A�����&w|����'o"�$9�h�$LsT_Ɂ%D$�^z]�*��"��(Ġ��_v�����Q�#�:}#$e,[tLB{}�b��%�*IȾ�M������E�/LH��.\ )�����bJ2�?n&ѿ�8y<N�Z�
FNC[5-������a(u��E���8��x�ep�U_D�i(�Lڭh7Ƞ�3&l��ք�d�����R�cf�"�����+�2�5;���J���\]F�垅��sd��}�Z�_�����>Ń%�$�~�,|H���r#h#m�&�N��0�=�a��!,w;$5�ݭ6�+vOKܓZ�:$�:zx=P�g%�Ǘ�}&�!����Ɨ:'�Dj؝4���Ȉ$A$Q�u�e��qHڤ�݈o�l���y�}Q�j���^)�|1P�on���߈�I�e�쓳��`t����Ե���$,���|���b���Z��w[O@��Z�yh�PYG�*k5qKP՜%7�&�/�<=l$L f�����%�Ђ���V��q�q�Pd��R�}x��5/H�x��$2�8k��*'����q�U�4v��đ�L7�V$0r��-$�����m�{�( �M5�����L
 M��TK����#�@�
LIe&h�բ(1^�ܶ����F`5;ٮw���}�Ң]�o��ە�k�B���ۤmc�7�� A��oޯG�_~~�?��'�~�����I��\��]�>Eg�S����Aq�A6��<B�R�����?�䓿y��W�R�UIU���O>��w~�R9�Jh4��.JH�>[�\A2t��Z����1�u�"�J�
͜K4��ƨ{�&p��S��њ{i�Φ�i�X��y��u�S6��T��>�|n���k��Xa������_-5��
�@�;���{(�=��r�F+�(6�.L��t|��͕�F�ïK(�I̋1���l��� ᓄOt�ٞn&zIz��z�[��F���|�z��I�4"�dgMs���o=����:���b<~c���v�>�0/���]��X�F��z��'2�2�vY�ב�2�% �,y��ƥ��:�.��y��2��WweŘ����M�Zv~�4e�KR�pz�!cf�f#0���s$L�������Ҷ���TM�r��)aI9S���U��(�߉9�7�@��E+�L���O�E��v��(kk������ҍ^D�Ϟ��Mb��r��e:ύ�|W�2K�A���H��<�*�&���bؿ
D�H��x�g���$���^�9�ƛ���H;m�MYzTe|�F(����d̝����a�bFf���ˉ¦҉��L��W"����N�)Cʖ�P�v)뤬���|�����+��|��׼������n�%�N���&Ν�;/B��N�|?љ�T��0c�����D����̩+� ����H��fLnI��&�Z�� (кo2� a����:�A������,�{���ܢ�����?>��S����떂}�������?|��Q�[z>N���1�b{�*5�!s2��*"R)j�'��b�~��v�Lc]���c���-�9q��'evQ;�w�~��V�LsI��/�'�hێ:��V �$cn:͊v_IG�<���V��� ww��(k$�A����3�aK������0Q�D7C=�τw���|��=�Û	mgV�/H)�LLL�=r��/���9v��ۈ�Bv�ң��S"b��hvi~�j�>[��x��1Wh"2C^��mA��r�1j�ʎs;�k�QG�H�K���F#�褶p�ɮ8�J^H֙�S�Ga��J������LKnE�|�2f�%�F$(�k;�e�ۦ��u��J��󗤺��-��k��i�Ӽ��n,ȵ�����p��E(�k�����b���;�Y�!`#��>�j v��|8ۯ��Q&�o$��h�Qy�x+"7ȹ���Q�V�-�7���ܾ}��<v��^x�O6���[�OO+��'��F-�}�+s_�K��h7�<"d<�2U�*�@sM7\(�y%�:�� �I��u��I�ܑq���KA�+!gn�������a�0k܆�]L�2W�Z/��Z9�K[F�Y� ʮGm��	[� 8|]e��i:�U}�ݟ��M���r���3�C|��Q�r�5�g:�	�`^DѲ��(��qeTF��
ɭ����$���x��M�<@�ve���o�t	ig�.�Yv����B�le/珅�k{֑Վ�g^q�U,4���E�:W\_��5�z��}tٟ�A��Y�.��o��Q���j�\~�#���FGG[��M��?}�����O�����_߿�={���=�3]x�[7��g�V}��lt����X��iV������{Դԉ�d�ⱝòt����p�t�)T1PqUe��E.�a�P�]>�9]h��k�/����IRvS�	\�)��C	Fl4��}���FSm��n�.5,����r v��͐�� �1-@�7����/
	�Ur%��@q���r!��mvg�င���+���(p\d�G"�*V<�Q4�rҍ8m����92r�Y9��t<����y�N�8�nvS;�l]�#|����,;?x�F�V�یu�a�y���=����x	ҫ�j��c�=V�8r !G%�T$�2���E\D:DR�}^�х��l��,�����7H�������;S>*��r�A�%��|W�D����D��D�8�@����^x�"�v�DĘW�	Mb@�}�����d���Í�{n�̙3l��>�R���f�:���7>UK㥆N�D'�v3*V:IAք&E��ɉ�<�D�I�0�x9j�Q��	���$uǪ�y�J����ߝ9>=���٩)�N�T��s��_a��W���T~�����ۋ���v��N��u��g�u���Y�_��SǻuuvV�LN�=V�KH��5���|���LMIv�<:=][����L��Z;Sz)br9fzeX�>���
i�d/٘�Sc�gV�G��2�>g�k$�s�ߥ\Xے�8M!���Gؿh;� a?�}��ӄNT���+�J�b8�D������_����x��x��ָ�����C�ML�����Ǒ,�-c��Eh7@�}�СCOMM̓���AE��y7HV��z��M
RfN��Q�^�a���9�_fl�������M�k6��l�������~���͙����by�w�N�=i٨2]��S�ɖ��,�-���I��2�!&3���]#��X�ZjT�� ���Qm��e5��"������A�w�n���V�&z?������20��(����k�g��Z���R%�@����Oq�ʝ8��@r���
�U����0^,I_(��r6 �
��Iv�����;w�Lϟ?��8q������4<��U���v�h6Z���.^�����{wף�0ȵ�H�E%��@0�SβD#Y%ZF�8 	��L'@2F���r�w�Q���Z����DfQǑ�*"IϦ�OQT�<C:��O
�Y����R)k'i�J�T"ɡd�h4�������������{�l	oA=s����W���.�-����إ��y%޶��l~����6ν��<y�d>�1	�t�Az�F �-�	V?�kl�0ξue���NS���N׽�� �7`+ ���V��V�]�q������e�!k ����v��Į�I�ㅙ[���/�����!��������GD��F���w���p0�UL��:�;I���ή
׶/r�'��ga�dgaa�llafbbj�p8�R��hN��҄��


	*2.,B|J�?���m�X0g�?x����sJh PK   �Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �X�r�44  /4  /   images/863c2d63-52da-45ba-83bb-7a6a6689309e.png/4�ˉPNG

   IHDR   d   9   ��}   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  3�IDATx��|x�Օ�;3��h�43Ҍz��fY���c�M36���ؔl��4H�f7�P�d��n
� I���t�1w�d˶���h�M��s�X6��g�?��Y3_��=�=��I�w�)��p&�:��ˏ`(
�$��z�e���}��Qz`�NP��G��ѵ
�A�>�r�J�]�g�w�8P�c����1dG�R��\x��w�%u���F'��
Y��"�g|�F%��]wB��DE�n_}cN1�O;���_�|/<B�(TJ9��i�°�PI
qO����nY^�k�t�5��~�g�svf4�L^\(�s����?�*E}�Q�@������@TäS�D���Q]h��5>�9�?�!4���ͫ�i�<��_^ZJP���:Ep�5ӽ~��d��	�`�l+�1~7~:��P ��.��S�s��9lǕs�q�e%s���W��p�!gM��?� ]�ii!V�Y�P[�����nTv�
�|/&��e��}e��جor�C�;�*��e`!ir7/)ſ�8��&�}O�| p�T�Z���OGj �t���*|���P�T[I�!mΙ������	�� qӹ�d��G�Ɠ%֗f�+j��{����Y���ǭc�[a��^>&T����=E��yXO!jw�@�$��x�eȕj��t� jܯ���JFU؂������5���(��A�'DcC�N�y�)�s��!��	�|�4FEY�EJ�
b+�;��+�R�}њ�f�8��d����̪ʻ�-�����RuCI����|�`/$=������$�������/���d۬�#+�s����b�@䐻F���eѿ�A�H(����-L�gD��n��B��$�2�
5"����h��`k��������y�2�����9OX�Iw\S�T�cʛC
t��ARi�7��J��j1�<��L��d5d��g��8ֲ�9r�[D�5�)�����I<_�рeF�u%\.7�V��"b��#V4h�Ȳe�
�U+I�!Dt���9�`�'L1���c|݂"

��'�H��/�/#�<E�7�?G��$�(���N$B�TF�v�� b'/^�X8 ��HR4�<m��'�ͦqER ��a|�6�t���+�V��'�|f�p@�A�����FQ`FA�
u
���E>��߻�o��I������'�3����y~&Ǣ�����������wl9%Y:8GZ0�҇y�@-
��)F�>�B���Bԯ��XF���</-<gƖ1N#�a��\,�E�4�	�}h�zI�{�Z)�5�k�E�N��t�] 8�`xŲ%�<�E�F�s�è���B����rݺu8�x/������3�(	��ʙ�	������H�y�#�����	�pP-���r�Q���N�ؠ���z㸰&��S���8��C�D��+�?���d�x���� kw���f��x�|H��a��p�c�c�ܹP*���Q�Ø]w�uhok���?MI�����|�y{N�v�oc��koEn�py��W�X�,py�E�yQ��	�Rꠁ���M�[�����uf�On��bƏ|j�����
��Dq",ΚTUU��/���3����,(��*d"��(�'5Q���o�j_����VA�i� ^;ЙB��oFTE�J-�;��N;�dR +_"��oqd������<o���TZ��M�ҍ_��70��;|^/)�F�[̄�hƌx�c����� �zb��Ā��������tĲ����3v��e���$:yhҋy�X֒���3�*�;q�kB,)`#�l�zh?�C��S���v�ۅ�'Q3�6��$��`�*�/]������V�P�)�!�I������7�
"ߨ��%s֩��Q`R����1dg(��Ŋ�w���c�2g�qiES�	\��2�U�f��#�i\r�#N%�AW+'A���N�kQj��c������R� ~?N;���
�]N�ƭ���>�˖.�/<�+K�bW��`8E��'�;Z�q��ƪ����� �Z)f��J<P��)����b2,��.�ß;�����Bzz:�~�pOl���P0�)��JE�M!�lAwg;*�J�Ν��m�aL���)��ͺ|�`_F��L��}>dR�(2)1�bA�ݶ ܁(����=�"/����IԖv�l�$��F�}^�fc�W��k�4p�4�����j�~����7��C����e�F������7�)�����E��+(��� T*5V^�
o��9�W�o�N�+�g%s�}��ВW�)��Z��#�t�)�����ra�`���l޼�BS�ш8��`���Ğ���}>/LYYE^~��RҚ>����.��t�p�4L�O�w,��gqe�\$�bW�OI]Ϙ��,Zz�"���ꊳ�td���:��o����q�P\��$�Ŭ*
Kv6�/[NZ�౱�ͻd�pYa�S��%e�O4��Ks.*)E���8É{�P����6~�"�^$�G;�Dn�J!�}I CȜ�8B�$;{���&�&�_Y9C���3g09a`�@l���*��Ҡ�����I�� �`�sOa.œ���c|��W��'O`�(���B@"?�K��bl2_Y}=.��F�Vzm� �O֓I��K�_7] 4���b!�����t�l�.�I����F#N="<+���MX�d)��3�>��f�8��2��G�h|@�N WGrM:�`3v�'B}1j�
	2��$Ԓ��L'3!��� |)�ϲ�J������s
Z�����r�r{J�����Ja�,�X�z�DB&C\�9ز�)A�c�)�� ]&�R!�t�1�2����%�����1��\���n,�d�V`��BPȂz�X����[��;7�2�3�s�򑝓Y�D"fx<n"5iB錦L��*���"�"���cG�,�b���فI
i�S��,�H,�1��ntQ�����3�U4h�V)ā�cx
^�.��#��jo���G㑏�P��j�zb>��#3�(|p��������=����:a���hAqf�e��y|��b�윂�,7���r�%M+�DNmԋ����Zw'�&3���0����
�0�#j|iy�Р{Њ̾w�Xq-�am��1-N�*�I�0�b��o+)V�&1�y���dJ��=���3���B(�yy+���̹��IW ��Z��cd� 	%��1I!��:`���WT��wv����^�.h��f��i����Oz{z��W�rr]�6�$��W��KN�'	I��V��].�8�9�.��d	m`S�)�$�AZO4�qU����/���d
1I�͚�P�D	&۔��tp���Cم[e��D}��<�^?,ᣨ^����{��9�I��)���i1k�uDj硁�x+��@�l�#9B #�ᘪDAQ� �c{�V3�2�bLF�R")<��]�^`���M��I�՞1��c ��K�2ݗ��i}�P���Qld �;z���Ѩ_8�i�j՜"QYe�ӓy1K8���щ��V̞33f?��q �H��&?��^�T��w�!��B�ϊ��P���gѮ9���	���n"z%T� �nC��N_'�F���ï4���B��@L�?f4�6�|%��~�������K�!Դ��U��O�j݃�0i��/��ȋ��~,߳�-6���XT8>�������X��*���`o��hr��͗����F���Yp^����W��?��y�l���C��2r�Z��N����L�%�����8�2��3M���`�P��?��$���l61褿���s.q��QR;?^b�3���pS���{�bG�����m;�}��~��<`PZC�Ϙ��4���Q�{�cO"2�K�6mCh�����|ț�Z�gя_���:���i�-0�y	ƌ��\�C��_�dMza��=�v��Di�,����
��I�OL3-#K0���r��j�gj�0�,���e��qqɣ�V��V��^w窪����2
�,!QzP���N��+$�>}u���L�b�\H�y�<�,b²��Q1kQb��Ufx�J�p��*����B}!�w8Ѝ�7P����B�� ���<�
1��}�a���Ԏ7���	dK`n�QSoB^4�!ˏ����z�gI�ggg'$r����'6�Y����]�Y��%���'�Y�����5�a�������I?��>Dy1���W���_�1�Y����0�)4�K�@m�	wL �(c�XRYY)266&2��µ�<
l�FL��	-�ɐH=>�����,�b���z�������潐gW@Qs9����- ���F��z��߃�������S�*�AQ�Q� "�g�Vy	
[O�zC.~�-J|e����"r^2�JX�S����.�e�21����5cnN��Y$��$
�X^��P~��рk��#��./�9�cH�L4.�&�_�4���Ξm�L4�eegB�����tZaI������
��k��F���<�e��&�͛�3T�.�J�Qkb#-����d*�]yV=|������~�4k6���5��5��h:�	J�(��� �7���0��� -�5�DT�Yfʧ�����t
ϗ)���D�ٳ¥�C�[[�-@a�c�`q��������,��cL�6,�2o�(�m�w\5�^����V��nBiuV�rQR�AA��l���(۲e��G�5�&w"�I��~vi����j���E��'~��X�<(c}�~��,*J����ɼ
O6�qut��3Q��Z����.-��W�&��@oKZ�!BVu@��wV]w#��0�4�BL�%\�P��]�h��G����0���d�1���z
˫�;�����3�:0��=P�����v>j�t�Uu�#��ijlZY#�b�2Aң䛴�������d���@�� (S�:G�o�+d�!t=��S�#(��:0d�O4V����dYs_���.,�n���߁i�0�>��4z���4HcMV�.@��
�nW��u��,��=���)�j���,�p�}��}x��ڬU���++xm�(�Τ���_�(0{��[pb(@�	A
Pޕ]�1��9�XW� |�p�_�\��()d싲��0Ҫ9%x�O �$-v��i2S0�+Ri҄���Bi���'1d����Px�W��H ���r9K�^wH������h�L)�$����+1m�vm	s�A
�u�S#��;���`��	��7���k\)����BSh��'O@`3%V�8m$�J&X�ܢΥ����Ʌ@�\M�EE	$���GCI�y��� <h�$�E�E����\� �(S�N54v�)��y�9����d�=����]��u�������²|,ep��Q.� �4J11����H�"�q���^�7�	��l��0$�-��#&���$ֺ��y�;:�0Y!$u�"ˁSD��[8JYLd���I)"���9;�M���b)�?&���a�U���L@(&�i.r����{OS.%�:适\$1 ��sd��')�GMTB#geTa�����_\��>ڇvM9ʗ�"��s��	غې9zO=}
�s0�܂o�d+���l!�L3���1؍QF!�_9f�z�|A����K�|k&�Q��+*��k���d���v�-�>�F��- ���9��47����w9+Qu��x?u��Z��2(���OI������L� K,|E�1r�
��T0�߼�(ܦ�ۗ(�%��"�|��J��q�z%�~�?؊�<tV]��.�mw=A�Cn���"^��|��GnENa6��V�^�o���6���h�Љ#��pO��v�S�_T�4E<��!�M�Hq�D�~�ɂ��jQ	�(��<��=6���K�%4\�W�_�o~�q	e�s��"�փvm)�0�S�<D$ȉus�닽���C�m9K���o��7���^)V8�HnJ�G㫎ܻ �������Rt�$#.C�$���P0w!����	lcƚ1����T�YJ(�Hó~s�)V���=�W�:��5uH/�F^Zv�I	��QS���	'�X�#|���2�������47�c'�(��/QX������J�t\������i�$|5���t((�����;�S�J�K7��軐�~�r�	[�nA��p"m��c~���m���2D�>��;�Цù�E4X�bK�
G�LB4A�D=m���Q\.����Cޥk��m�J��^�j���~UC�Ҹ���˩�����?z7߸>��y�k0��	B�c�h�)ܩ��R,��e����m)�Y8Ϲ̅�+I�\�R|�`/�񲼌�����C�/�݆��mDp߳Ȣd1�e�1�B��|ь,�y$�;ȳA=�XZ�ZD��4��?����bW��8>�	Od��I�.��D�'5	.�F�U��W}N*�.�JMZ�
�ysp�=O�'�[_ߏ�;B��P/d Vk��ɿ�^�;Z����H��EE�y���2^4���$A�S�YX��.�p�,"ީ��
������U��>WP��n�
'�I:#��5��p��ID\NH�܌�-P.�k(I���;����1;8����<��Y�p����|�m�B��,^��4�Kg�CC�;F�|�������08/��mne������m��P��XY�	,�f��df&�C˵E�y��>�%�e��M/�	a��4���8Ո6��!{�Z��0��q�����GD�Wμ���)����j�~���~���bԉ��s
&�!]K��owX	M�'
|�YrbGG����4-,��+6!��g��rW��S�j2 �����%_O��K>��7�ʠ���Q^�x�4�� �6!ߠ��99��g�X�\La�T�%ظ�a�o��8t��W
ʑz�����d-:�@�澽�B"˝����e��Ƴ��U�C���D��TY
�Y\*�����3��4Қ�	�u�#/S/�Ѭ�"��F�IPL1ui*�d������T@,�p�Y����`�L����i����#�ټ��%e�a ����8��ٯ�Y�\e���=��N@9w=B����10k���3�"6ы�Yk)菡��|P�����Mz`1�aH��51"i*�e��7 +�s������)pM�t�(^��������d�2��@!d���� +�4h~�9�����7-ǃ?݌�T.[�XY"�g��>�yF@��o��`6�đ��G�}��R��d�xu���`���i�ub 'ljb2*D?wu1&�8�}��F��%#�:�
`��^�ko�d�W����L�)�V/��V�D1�\ (eX�7W���Wq,�Z4����5�"�PB�ry|�+��H��������
�|/�+uzt����1���[��k���;g1s��)!�B�cmm��J���;����ԯL��=O�;5!���C~�p-�nzi�������������9�����mCv8;Jy��]_+��Wϊb%���؎^�E�o�6��'EP��G��"i����q���o�EGn fD(��S"m�iNo�#W� ��}����ta�~4�O�OMvW!�w���.��D,�;��~�$a����̫��{����3�'�͜9�	d"�wܺ

d������u)���߅�C�I��'�a82sK��?}�'�(!S�_����,b`�KM�}�o�9��=�	�<BLEM0�CAt3��fӗb�zX����Az�W%�Fw"�oL�kj	�/�X� ������F�kW�:.���T 	�}B���9�!*�CSƖ�j1yH��!~	�,M~����3�L}׻����Eݦ9�V͇*o��8�@E�>�ׯŲ�7��j���ڄ�k����1�Ï�ub��^H�4"g���Z3$���m%P�L���U����4�}'�,�i�C�J���5���g`P(�4�&ڊ�'���vA)�����7a٭?¡��)����x��WXIC��.�ȓVC��]�5��U�>c����������7"Ik�@�ϛ˫�3<w��qՊz<��a�_�()���C��Ԃ���$\�}��P��?���rL���+�W.�Ǜ1nWb�=�0����[̿��'�DM�kI�YĞ��G�َq
�栜>����#Ƨ@��/�X(w /|؊�
f�S^
��9��#�+z�1���d����Ԋ6���)QOc�;�+���1��;���ޞ3���*#�k�H�AG��{�R��u�E�v�oOT{]0���D��^�����"l>8����
1�GN�/5A���E޴�LK�?�,���ٙ:dN�ύDi������&�$wc`��U)>J��B��^Q# �6�6��5��4�eaqu.:��o���?윂I+GN$����+&���<��ݎ]�1�_���L�B.�D5�v��*A�2�w��!ƒG�H�`�Ab��j�f*�:� ���.[�`:��t��n ���>�dJ�6�K._���q�?�"#�Man�aU܅%�_LL�104�J���Ct1�|�#b�3��D��x���?;",���!JV$����cQq/��J��=�E�a���� ��L�q�� ȃBN1x�I" O�w���Ţ*3x���]by�b�H?���@���r��a<���`P��G`�������X�B<����3��hǰ��
l=<H���e�"������;�E�M$�=y����q�{'���Uj���UF�Nq�W&0נ�Z3�g�&qiu�(���rj��r�aF��g�)C>:=�ݧ/���c�������MGj���E�������7�5<���Sw�r�,k��r�D�JC�l�x@�����. ��
*D����	vŎKg�����I��׋�$p7�MLL�47VTs1��)��V�����h����xK�{a`` ��'���/���&1�L��*��Qh����'�6�f5
u���$W�F�Q���i8=�'��|��e�;W���k�~��k_�a���O��� -��A�E���a������E3,w�������.V��x�¡ni����c��)�J�G����L�#X\����E5Z�L��B�9���K����Rּ`���Ԡ��T���n�9v��w�����N�˿S-��ݙ3g�5���)�b�͞=[���\�뚚�D�(�B�|nVx��? �r}q��"0E�m2mAZ����:��B�D|�NK1@�DE��Cl�V+@X��������?��.g�ěs���6��=�縮����s��Y,^L�6��-Vd$�u'l���ķD�e_�EK܌]�⫴�tOu����o�i����Z��������]�f����]�X�� q��w�+7(�j�R��6��{����������P���vu����E�Y����wZqM��8�:J^A���������0&+���I\7;#�b_��	�X� �{��>�z�~�.M����^�߃�,�7]Z��3��<�~�t!�q�J��u��!�� W1C4?O��B �g���$�=�nű��T):�T��[ԭ+��7��E��2��X�ĆJ�]�0�ǓǂJn���fƂKZ�HB�м�%y>��k0�"7��*J��i1�GŨ3�����8;]��r�T�g��Ti&fT�=�F�c��3HגˇŠM�Ϩ`�7O�l��̺?-��:�ڡ��,���w�=�a�|ihr��;xՅ��d/n�I��S���8Ol\�_l����	������WH&W7��Z�ǣk/)�A#	an��X��G�����Be�d���`2h�����zX ܨ7��0��3���Y �tr�����H���m�!�'x90g��@�K���ꪫ��w���?&����)��R|I�`ԫ0<��3�]Ƙ�HÓރ��M���'It�՚��7�8�j����?)��%:�����4ؽ�h����2Q�W8;({eM͚f]1ц��B��%�o�Bn��#S���1��$)�3����9.$Af�Y p���B�G <M�,�@��;�qK�	���=A�^!�I'Q^�
O0������6��W&���u�I�?�/��?�2�	����-�����Pd��N[.?O�'ujŻ'G�;>��<:��������L7MN��s��؈)6���g{Fq�g�Q5ZǮ>O;c����n ��T�
w@r�߃�,����
��77vG{ݓV���m�}3�t>���|��E%;����|v�\�ae�Gd�<����߹��e�;Ш����v����w!
���2ds"�w��U��h4�]�,�AJ����.��\��x�oi�*0�4;Cpgֈ�A;<�s[�t:��Oa�#C)}�~~.��\8� �d�H��fJ�U�j�:�V�"i�
v�A@M�rV��310>��M��N"��}�Z��㏧��qLaZ�A>ɺ��n��СC����/�In`��������=�PJH|������>+�2�2u�_~vM�^�����M�I�'���	OB����I�E�`�����{p.3#߈�h|C�x�͇�4��u����,��OG%�t�^xb�>�D��.�.D��?˘O}؇rY�<�y��h�y��������6�B�����)��Ţ�ab-U��9s�@����c��3 �9�`��F���͛7����𹭭��\E"�(++���?��%r57��!0��|�?�2;^��kPQ��o��6�P���'y�<v�5�i�6���6wD�@��bԫ2�z'��7{&.ǰ�x~+Y�aېC�![���s��a�Gm	�T�vb��Y���<��0�r�%yN��&���Nʝ�Fy.���yByy�ؘ���-��o|#���m�X�,�dl��W^y��7�~���rޣRTT���~:���,��۷�>gww��ǔ�x�l�:�������ؠ�0����8q�(�����4�[[i�|�/�������/�\���ф��®�Ax�5�[���+�'��?�8K�:���dͅA�0,I��KYbc�";�6F~v�X�QPǶ�����8k���늛)yR@�J�;��Z)�ׂ����A7ɔ�kqR�����=|����@��D��<8���D.�����g�K,D���y���L������75!޹��E����'9|��(*.��9��ȊE���ŏ��)��q�bL(��G,5�l%E�®kIM6�orh���v�J�);�nran�O�H��8�1.6�3������"-V����z�+ޱ��3J ����7)�1�܂�+����b��(aL;��s@f0��Ş?rG�K$|�$K���$#KY-=��A=%l^�{�ݸQԲ^=f���D˰O�,��<��ݰ��_��}���%�:��k���?�>a$a�q;v'o#��`��%�����~�áV��~�79pkN%|~q�D�]'�9��$eӓ;ZŠ�t
,�2��7����?�Y���c���©>	y�
�/���~�l#ӿ��kp�w�ũ�y�`���c��`Wd�#OG�3�E9�ĉ��$Q� ��`2JZN��#��� 'K,,<���KX6�ρ}��E+,	�7���w%r�v_�T��1�r�3D�UH$����M��=x����3�>�<�}g'V�XN���a��#��	���������^0�����:9�n��'/��"�&�Nn_Y�bA�-C#������z�
oS���mV1�	wr;��h٘���CqWǉ��D�τ��
]&e�!Q|�A؜>�R�	E�K�N��S5dA����,��������� �[��M�6aǎH�c�w���쿹��L��[o,�� +��p��J�:X�,��m�݆���ȕ�����'�r2@���=ѨLt��&lB!�J���cb�P��:g��&O	��炰}�y��ܸ�\Px�o���㯞�KAym��wBq��t����4�����<���#Ҭ�y�p�B�1{���s��eӀ'�]�*����ՂOs��9�F#��S��0��+�*e�[t�*��صkn���J��o���`Z�_~�8���ڵkEޑ��7�½�ޛ�i�ݻw�{O?�]!~�W��U����cZR��٥�h걡�4��"�8&,l=����(+/<�b�PX|�ꚪ��C:?��|A)�ca*�-'f��&B0a�2 Y�JL�|����Vʝ� ���^.73�Gۭ�ʊ
��\���'�d���+f���;0I	S��5���6[���t�ZFqm��ܗ�yoG*�嘛,Q3h��̚.<���c�&� ���^{�S�M}��T�%�θ��Y�g3`�s�5����N|Ŭ-��5b1'K�)�[��[��~��3$�x�z��lv�[Ըea���-N�1��ely�_hFسX��~�p�������{bˁ�}_ZP}�m�ό�@�&���cŉǷ�o��&n��&|���H�S�Ɠ���Kf橡��������!����bQ��y����(����t�bǅ/ę���ڹɍ��v$�N�Gc�8�������Z\_��Ms���BfN/��%��c'�y�w����I�:JV�%^���������67��O�+'w{������[X�Ȭ����$޹��g�,$� y�H?���-�z�����w����Y�ܘ5�߸�2셾�����ՠe�p��^��R#��^c�N��V����q]��7��^;B?�!ja��;e��h/Z�'E��-�፠o2gL�)�3�E.P��jc�`���r�6@�1H�'JVe	&��0�?�r�����#�uӁ��⭤,�E��.��}�x��P�N-ULo/[8o���f]�����Y�^�kGG�0X��T@xs]��3
��-��!�>?=��V��Ma�3x@QKQ%�,�B0���C��']��LBŻ�2�zg��V?lubo�K�a�Q�o�Js	~��0��#�sR�g!⎢���P�0%b�؉E���w0�� ������ҵ��
#}oZ�    IEND�B`�PK   �X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   �X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   p�X�l����	 ��	 /   images/9b0fa5df-c9e3-4cc5-abbc-d39b3818cb07.pngl�g4^��u!J��]�Dt3J�!�ѻ����^"D�]���$���e����w�u?�g����k�o{�ki�H�鉱��HU���`a�aaa�<!�O�3֘������êc���l��屰~�?������\��<���{���^�����he�k�	v�wU���d�i����n�d��b����.e���.%�������?$!*��ea����?6R1����z�Py/��k�}O��i�U�{���y�*r>Z	HgT�bN|���M[�g��A7	`B.`�l5 8~�I�泭7E4ou8�����>������(]����4�Y<��8ķ�-_ �n���!�c�;;!����_]�}����oB��z����ׅ��a�w.�wǑ�[,�	5Y]^�Y��/Wn�>��u��<`�E�;>L���U��F�p=�y���ߦ]��혎��~����(8��kr�������<�A��އ�&��o��o�ܮ1�C���d�w� ��5��(p�J��l��P��ڼ��}o��Ǆ������>*4�� ��.r#�6�>n�Av��H�6�����I(�j2\�4�x��<�k
A^�Ս�c��!�Mۏ�R�0s��+�v���sEs��RR6���	���wk�k�%ߙ۝�BUq���H���Y����>|8��6�� �9�],���.�2=�ʳ?�X9����5"� 0U���Y3���e: �R��;0
���9��G��ŻȪ͊N��B�p���P!�B$3��JP28���Q]��l�Q����6�g��0Ӯ�]�xNaB�!��m�X�?�0�0�c�D��V6�<����R|b���ƪ�oq2��2(6~5��|�}MF�h\�����=�.����ɿ!KhR�#x	C�j��;:��ÒB��d#we+�X��d��i[�nW��,����q3iRa��=��G�+>è��Ȩ`�%���[�~�d'����i��і��r���;,!;`nN�1�j49�V5�1Ts'��W=s.�9ʲn����<H@��:s[{7���6����
 #A�i��I�5nN><��:�[eV"�*l
�Z;(R�I�A���g+-��"��!�?>0��s�,l|�C,3ː�/%ᑮ�?��t�c��|D�<�"E�'��!����7ϧ�
9�~c���S1N��i_��cb$l.�Rރ(���TN����W��j��fm��t8VT�{�vDA#lMFBل�K���D����~|�5���4j�s���N���͠��&QAe��д��G�����V(@��&�~"��T8�* ��ɽ��K�Z��(:���X�qHM����3��?i��\F��Ÿ�o�X��y	gՃ7I����2Xw�$��
�A��42Eå�RN�%0٢�Ea{U���M`HsL&n�aK/|�����k"n���Km�Y��2�HY��$0��Z��n�.T�?^s�V��8��f+��Y�M �݉ �c`C���ć��E~��{+��`���"���8ɲ�f�v�U���!���Q=�ӯ��ͯk5(��]��1-�������
�7�CZ[��^�>��7��1$��q�N�Z��ĝ�[���Ҹ������~M�n�כܩo���~�����q���"f̊�K�eg���#+�5�B7m�䁯��)i{��M�
�Mq�ތ��ے��ǃ�'F�A15��M�jװx�b|�{I�h���)]��_Z�����v��#�r؎L��Kɥݣ�Kt�mv_߭~�ߍy��M*��\���ʚBM�~<c��I��Ge�y�JvU��v�'�ZR����[��m��ea�o������	aH��߶t4�<Ȍ�w:�SG3~`,�ʻ�1��'gi�-�����h{8��r��5RL@{
Dk^��L;_|�*��p�����D5��ON�6�JD4��ЅYT�]ME����`�)kԠ����Dժ���72���x�]�M��v����vb���3I�k��D�\3�{zo�I�(��c�I�=1��N#nFZst�u$�"�N���lMss�J/��\7Ȫm�R�X;�7�M��wL��n��!�6�}�GD
|�G��*��%����5r@ �Kuq�Uvf�"t��O�.���4�=+�NGH8YL���1:���#�P��g�NMa��KsR^�4m�I���a@�[��4�6R��*S�C�uW�>���Z���A+�Ӥ��VB��}<ٻ��i��SH��A>��3���"�?�vp��6�6(�HW}�-�ID�{�O�G��H��$�oI�3[��t�a���)���&4%�t񔯜a�(bt����M��������Ql����yQ��
��
����#����#|����OC�ɒveO�;��&��i] �"��8��y�bk1����ʿ=tn�y��"�I-���m����y�e�q�ʜY;�����AShө)����\
O� .��Ǻ�V��_�j1���S�`Т�y5?/`� 9o*�Р��y��ު���b�M�#46�/ڜm[�~�b�U0��oc�ƻ�d�#���	����m���e��)9�\���ㆽ	v�m�a��������t&���7P�Pk/E��J�|iz�8�|�>Xz�^�;��c�a�_�{�BP#���!ZW�y@�7�t*��ʅ�v(�q斥���VN)��̋D1{܂��5=Y��k:��	�k��k���P��X�fbb��U)��7���e�B5�1[3���:y��I�#��sOX�ZĪ�{���Y��TL�KO}��6�upb5�D���/m!/�M��Q�w�v�@/��)�ھ�n߆]!�Uo�9�va���
S��H5���Lh�����p��R��(��/����8��hrė'��/��~�������oO�ߔ�Ęm8>ߵ:� ��P������8�=w6��m��� >(�����t�ې�/94~f�L�qE� e3����x
+ǖ2��i���!���,�;h����f;���I�a}��Կ&�<Uf���s�VX���c��.�L3��u��
ú(�'�cT~*c�ƶ26Z�-��W� ��g�^����'�d��6z��_�z��\�8 �\7�C��
�^f�scPQ�Ez��@�o���� r��? 2^�����H�UwZ8M6W���%�O*y���n�.��s	����*�����q˴���q/�uj��Ѳ����1ۋ��~^3��y)�>��6UXNI`�}7���J�Ě4��f5�Ov�eE��K,�1gg�G�y"��tw|� b�u��`�~${��Y�����c�&��ګk����/���
��Z��-*0�8W�����K���xv�SvE<��}�Q4���S�s!�OV�e0(o.i{�������Y���#c1�Z��̃�b��#:�)�R��X2�c�o��tɣ5���Uy�)��H�F
Z��5#)�tq�|��`\eq3��s��Mns��o8]��[OV���n#�F���{#���2T�����?xԪp�S���F� ��'���R�u����C� :�T�<w�{��lm���e���$G{����Û�*�/1ƾ�Mbï�RLs>�#�w\X@L�>�.42�xd?-fm�,�A�3��é��A|�Q�jv���5D4̂qx�
gH�T���n���h��F�;�j����φt�ٍ2��<ʷ�A���:痰���r�Mau��f�O��Ny,\\\�ϫ`����D�u��Ś�T���9���;"��v�f%jp���̀�i�uZ�4�'u)o�3މ&F��'�U�e].9kx��W-���ۅ���n%�<z��q�jH�{�i���3���Y>GF픘}����� &��2dC��� U��vQ���B����K����9��Hz��P|k1���~.:��,R�=B�q
R0�:�[i"�r�՗e��7�͌�t�����%m9�4�y��0�d�	�A�m��+��e؟����U��J��#�Sr/�������M�U�B��s��<�15ft�Wa�"���縷v�2��X�aT����� �z�W*��dG����ۋ��H
��א��E�ޡ�1û����2�C�Q�`8�����I�\��pZܦ�o�h?�Y��
GU
G��$���~*u��h08gvFJB�yS�����!\�v"��r|����}٧����%��f{y�+���ց�x��%b������0a	d��F�"9Z��^"OJ���xL�B��"��9�H��Ll�9�xP|5�8:p,�L��zZc8N�����S�#.$��?&'����V�-5ej�x�� �{h��@����T�Ѯ�Jc�+u�X����-����HM����8�!ɳ=�&6�#�HS1�f�hX)��?h��zM��?�jw~'bET��fB�z=h��,�F�������Sܴ4F�@X%,��ǋΙodZ�c�n"M��8߹ɧ\qGE�͒�o�$��w��M��[�OXߙT'Z��ǳ�LY�y��H��~Q�E��Tw!>���fb 8�?*o
��L'I�lO��l�����L�pX�q�D`f�/u<��2������+���>� *�����Ǚ�aZ�H ���w�0��"�� vq\n�~�^3���.��g��_��Ү��M�%EF��㶐+*lbBث���j��Wgϭ�駄W�J��:Ädo64#~̒����W}z4��������^��R� /���bL��H�)�+i�^���1|�����z���*�{���k?��ޒB)�/ ��l�_������dEſ=KN�5	��j�:�Q�l�y���/F��o�BĪįԮ��㸶�&E��3F�gBm�`�"l�1�-R?��,E��h�	ؼb:%����n�ʪ��^ӕ��[CfGea����e������I8�[uV���q�4���$^� ��6M�fxR(�|yj��28���TOME��^�Q�E�ܬi�*G؝�+-v��-��S��@����JF�jJ�'e:����eln�c�&[3�퓂 �8~�%g�0�޿D�k�+c�S�+;�	l&ׂf�� t��b�7��2��`�
�b;W�?|ɪ�2{��L��A=���u�_�3J�uU���9j|Ϙ�1�5O11�F?D4�1���'�����:j}�������_���@W4��5܎>b���l�3]&-L��Dg�y��mAluG�9���z�Y1nfuɗNG���7\�o
	RO�_��U��6W:c�e'2�?5�, �"�Ke0ЩJ�e������9[�MS���|7wg�g�����+f��ieJ=MF�c�3+#n�,�;|�N�%s�����b�Zg֭l�=��.b�?�Ty���,aj������^�	�ɸ�]2��y87�!�a6�\�B��$�I��N�z�Z���N{R��V}?�<~�����=�Ӣ��da��N�b���+n�TA\/������|���<���X��_)E���z!=�tvp�!��h���Ɓ/'�N�;�s*XW_ i����/E1ؓ��C�E"��yw�o)6+"n�+A��<�;��Ԛ�7d���j��M�p\R� t�|��u���֍�F!�����w[��MG��ŉu`��	^��\�����������@��VL�AU��2���ܯ�c�B&�*Pd�OQb���K�T�­ʦ,�MNo�"ީ'v�l��ַ���K����Ub�y���Z�$6���0�xSv������SoL�|��Y��zѤ�A��<�S6Sp���e��WbAKukq�cves���`�U��U-�� %)�<9���?��^���-����k�ZD;[��J�����}��0}���ga:��DfX郎�j��,df���n�8����ñ4وi������V���KBL������Bݯʃrf2)ȗ�]�V/F�,N�@&�&iWS-i�	z?�4������Z���F9P�/O��Q�3��g?�����:W�F<&]
�/����6�๡�5
(��&{����Y	ۜ[?h�v�h�9Q%�p4󒩤'�PXDȔ�k��ӑa��;znq� I�գwq�J���o�n��}J`^�C��|�b�B������4�J�������2��͉�Ҍ��c������])�[ՔJ�$�Jfe��^ʃ���k@b���j6İ��K�-�`�}�c4�Fa#;�^��Z�&,|�ru*x����<���ұ���ӑ���V��-AŜ	̱��T5Jv<�7O�!����iJ�V!�VbH�w}���[=�b��3���FD'k�	wpb����HZ���?L�1��W9��Dj~�Q����o��
���/'tdg�ݽ��f�<E� �F۰�E�~�&�-��8Fv��A.���bĂf2&Q�ڞ9����Qդ9􋤮i�L� �h�����2s92����l�"�p��@ ˚}���A�AQf;[dpQ�3�}b�U���k/G)�0��<�̩��%B�H��9�{s�¦_R�����Y�cM����������ɋd
����i�U��4�*B�#���tt��S~��-g���pr�a�W6���|I�Z}~LZ�8{�F�rǯi@�;�;�"=4T�~� ���h�������^3��3cH�)k�!��������ݛM��@&�B��l�����V�0�CC}	
wm�GE0��E%���Z|z�P<,H��vj�&Ͱһ1����{�����P�dɍҌl��������������G$��<!Q�K!��n��3}x�;�(�T}2R� d�)� U@6c�Bh�U}��|x�k'�Ҥ��kM�����I���qWuK��	�wH�6��J̛S�En��)4A�*f�QI�������J�Ef�g/�h8�Wl��[�.�w�%����r)eXYl8e*��G���'�|�.d��8Fa[���]zV`=����|�K�$<�.Ň]�7�*�*��ޤ��a*n��w�`go��������	w��+��~\L�q:v�O�5Ŏ�����c>���s�P���O_z7x��U���-U��>����Ϲy\?W��,x�a#�ݱ���%���Y+��;ط���h&>��dUޘ4�k/T�	8Q�]�I���䴓F��w)p�u�<QC����"�A��5d��q���7X��z6�b�2�O>L#�	}�&53�"x&�[
,��s�(�		+Q�iJ�^�K;K�Q��`W�EѺ�9bE�o�Y�԰Ǻ��*`ᔿ+�^k��e���Yi�G	�fk�x�|䬣K[�e#I�zܡ�B�.�&�Pl$�}��c2�Q�PdK����\T�b�65�����@���Tr;k����2����_?�Bo}B��9Up|���c�7�urD>����Լ�o�]���i��RiƔ�k��&�}�Qݠ]���'����oh	��^u�[����9Pd]��c��?���/]~X�Œ
OmdI�����!�����_1�55VM���"~V��rQ��A�)i�?����CS7&�v\EJ�({��^�H٦Yn؆;F�O����z�&�Ӕ0hȓ�sr�FI%�����`N����Ա{-I#�������Ń1�P�T ?㯼��q2 ��ɬ#;;AH��&��C�1ܫ�N���UqE6(^����(�˽?����xމ2�w�!�˨B�g$�z�s9i݆qEP�A�U��7S/��/{�kipY�[{���y�zb����w�6��R���eLh���v��-��vJ�!B�!�oO��MCǚP{a�a���S`/�XQ�TsK�F>�k}��NE��>�geW2�f��PR��Y�K֘�uS'{G��ߨeG��p;�@��r{X����_��O����� {J�a���-.�RGGU��Ⰹ�����`|�	X��ӻ�V��ɭS�3��^�9.K�����6�D_ߏ�Ӏa�MC(��Ti�n��Y�ʳvJK���^^^�1Yϲ�,����&Ы�%!�|������s�������@d��ˣ�^�G�����(��iRe�險\2���A�B�q�B������0�i���	�K���4_�24�2��\�´)�L��vhDuE#��G���! 2h��v�u�M��Cg��k���S�Ut�)��\�y�<�����w�c���~o^���K��?Q8W09fn���\,�=�\��)io.%7���'dpϚ?��t)�t�����cd�k�*���T4}���	��C��&��-xbiz�f{���Q\�iWP���-?LVc��ڧ�0h'��ڜ���g�����J���a`�|UY����NU#�YD�!{5��B�\��;�sc1V�N����֊Aֵ��:�����'������L�@;�BJ�ƾ>3#0"M+�z֙ܽ|@�ԊW�{���=%zO�H�]^Y�[r~���� �^�����*��J�kʢ��'�l�o e�绉�XZklf�_��.�"#Xc8���J��X�=�PpE,Ӓ ����N'�t�I�G&�W��9����x�Ω �����&9$���_vpB��塺|kc�c��c8e�Ʉ~�:j�3�������(�%�����v�-�WOǇ�kOrù-0�u���FG�M/G�g��F
̀�%�������W� ��ǆ�7Q$�۸�^��~�oV�{����|=0��^�Q�H7��3DD�p�5��C
��:�q�m��0�����`�&�4�M>�F4|sg����*�G*J L��Q�	:E���FI�|��*���K`�$�7� 7f4nANjlP����
cZ�t�ˠ�q�PO�����5Ӳ4�"Ǖ��q�J�D~}��_�1�_���t�'��L!��Ĺs�E
��-d�+���	��ː�])����x�v�T�ڐ��~$���|�5����uc�u��Ҝ�Kwy�>ݧ"|�{zth��%�n����p���b�y[!B�׹7���������/���ײ����n.�䦻MM��k�'���ut��]�;b��Ǝ?�{�1=C�ٔ�p%���P_Ao�O�ז>
���P�*��JPҜDPnݯ��m��O�5�CΦ�o��(i�m�d�)�$���A9��z����O��])�poÚ�<�M�7�y�+חuV&dl'>�GDA��&�2P"K7W�D�w!D��U�;Mhq����ʔ��I]�����)	&��òr���8�������ʭ;��) ��
������h2��$z�MD�4�_�ј�p��9���U�%w����<��n�s�M������ߗ��{=�e��YKF�,G��s����e-�����U=�T� �D!���ٵ�K�iΥR�Ź>��c 9l�����ٔ�'��ˏ-��?�}>y�Qh�r�FIB(�\v����o�leeu*�9��n�E(�c'dX[�,L���q���?��FV�q�����`��?e�{�lԜa��UBu!���:�-��v:5Ѡr>�,A�P��s_tS�~�$r>��A�C�-�d�*3h+��A�i�Pk�J��B�X�V��ʏ.��ա����mY�l��U�,��9�!���	��z������%yG���3�\U|k��&3:`֑yjr`�-��f��Vگ�����0yE��B�����{��K,!����h�2���%Sj!���gW�Ej<��P�����+�"��y'H2����Ձ� ���� ���hU�%������F�?)_��,����'?K���x�ڣwN�F�HpB��*��E�]|�'M�*_/�J��5V"�f�
bb
>��9�#��Z�����%HmcJ�����V��=ƙ�eA��2j����ɬ�A8�9n�r޼�*�	��/q��oK�e���{ZhQy,��S�Bn�o�F�_�޴�T����dQ�[|�4�%�N����[A�����␬yj̼+�+8u!�M����K�ڋ#H2��dsq��խ����$kmtrv��G=;[�7�͎$���ԑw�Tĩn���f��:��QҬ�N䵉*�8O=�����7dFRm��"�GE�7&�-I�h#ç�Q�������n3�7�D�� ���V���$�D]qX�x;;�h�3���r�!(��N@&�3S��Z���3Bq)���,~������R�+�X��`$R3{�Ar(+^q�Q��z�f��b�����Z ���e����6眖�}��ȟif���:4~����Ψq�iN�u��g��g,�k�A�̵�c���ڙ�x�X62E�j�=ԕ���U�����	  �����M�%:T,ٰ����U��
�"~K���b$&m�T���B�ӹ������������f�Wى;�_M�-Pʦf=����"��s,�#�Cӝ�20ỉv��z!K��:�{>�Ji�*��R��������h?�$��*Y���k5� �(��J6�Pc�ͩ�"wP#UQ
���gh�3����|�!{��������9d��m��:k��O�p���w��=gN��\U`i/�T/?z�8��|֏��Z��V=]"r�Y%1�g_ըj��^��~)ŉ1�=�Q�D�߄4����#�Fabj^@�����k�ɧ����ET�k�U ��.��*��G)Y{.�Ow�m�G=�*A��Pw*���nS�F6�����{.��l�)���3,��i_��:,eG9K��/� ��7#Hu�E��9�'����i�~ntM��#=��"�q1���,�������T/��7R��e�������5M�4U��T�]���2���j4�bY7�K8,bmq��
����oc李����4f[���8f#�[ݯ�m��{���&4F���~�K�N����Γt7� ��S��y���G[���e_���7j�H�� zT�����c^)ct �]8!���u�ɝ~�ӎ���G`i_7h�Y09D�|�rg8�J�=�o������b��C�G�:9�F�7!��Ƶa7z�x��9$<	���Q���YW2藙��y9��J/�n� �#�U�׻��z!C�;���>M�8 �%�`���o�7�g��0I�V���i
@sn#�j���[�n䀛��C���-R��'����K �jM�J�B��IЗ�Z@��"sҫ�Oa�u(-_lڗZK��'���Xk��-����L+3!B���eK�e������2ݗx#VR�!�RCE*ŪH�5=��7��mD��ė��[W;N��\�;	'U�A�L����2^�����%�tҀk�k��]�7�1��㝱���B���U�>?	̦��0�N��2�[����|�_ͭd0V��S[����s�<p
�Ș������r�7jL*H:^J#_�4��;nf��<d=��f�)����-m��ڋ�q�����*hZ����R�Y��JZ�1@9�PN��w~��=*79�ծ"��B��ɗck�ZdwJy��Ks�S�r��t�|�1�7�@V+@[��f�ȠЧ��i�+��S�Վ�R �t��X�c~�����7�Q�|��q�����|�~��Ýߠ$6��~[{:
���qb�нd|��b�0�/� ����t�^y�����Z#%F�dS��5�DF���ގ/]-����EYN	d�E.*ѧ��<�5dy*�.�'N}�[���-yw9X8(����K*�� N>1��݌�"#�C��Pt�%o�̃Y�ŧ*���Z�rd���<�@��Bj�&�&~t��a˗��>�׌�bf�~?ܙw���qi0^�`c\�>k+��O$�G���dX���d�\�(t�<u�V����{�i�{�r�w�) �D�����S���"殢�"�Pxq�cc�H��H���/���b��X�)�&�^�I�zq�����}!�.��J�H�I*�1GYV�v�?�
�����r�]fQ3vy�c��Tn���҄e�t:on�0{W��2����[�EN�}P���N�%���C0�F���KP	�{�3�4�3Ǒ�x�����dӸ���/�^���_��l�$b�<]�G�!pJ���^J[�)��s�)�n{j���	�J=����BBK�O�E���ǀ�D�Xl�jj���w���Xul0j~�s���5Qg�g��=���s���N���D�[��_/6���m��|�Xz�N��~-�	j���t�iw�Z��zeʘ�;c&~H�����d�{3�aʚ��rW"����i��[�q�!��D"~a�M�_�FH����82>e�Oh0��W���Y�=�o��ffJ��Q ,MLV�+6��A���am��H(Є� ������
��#0Z�^�g���QǬ�"���E���T�;�O3��,��	 P��h*�ު����]�Y�!�N���]1�����ck}��Yڞ��=�����QX��홨]3�^7s�,�Ԇ���� ��E&?��%$?i}m�st�q��!L�\���wԌ�����M��e�X[�Q�{f���91��VC��c��-���*�,�N�OQ�5��ߍ�;O�Tg�$��;*x�ݍ�����*�M�Duw։���Ul��*Tb�7�y��&��[�"7,IAT�o�{g\$�TY�cO<&(�;QP��qF��U�G�u�����+JU���r�2�4;��<�>Fo�o����<�R��$�Ʀ=*а�Қ�٪�"K�{n��h["D�Hg�x��Q*�Cø���bIS������rx]L�f�kC�ƻ�������,���1{>���ə�[��ME8W=:��O��T�����z7���4�8<�����O�m�� )xK��k�{�$A{����_Su|{�,�����x��`4u̺�;k �*D�H��.����I$�$���(]�ǖE�NC����mz#�%y��w d1vp�a����(��������C�24�+}/K�}�t����*����A^�z���g��V�<���ޏ�&���;��FsGa�%����y�:�u�#�R���S���G�_H6a���?�RYp�I�
w7��DW#ϟ�ˎ˰�����q��#��7�~v�\)'����#���������-�Wk��·2��_��v	Q1��������b�ℵyWski>��_�i�my$)��I�����z}i:��3�R��oW�rBI2���nf�G�i���0��I-��~�q�!�Od&�aenUs���1�^*^ol���$b�&����Ŗ�戳���#����[���Ĥ���1}^{w&��C_!�u�ڬ�)�m��W��	eL���7{��#><hI�3��t��B��޸5����c�S¿����ߚ���賫a��{�� �Ď�c�j�8������h�f��1�LX��a�@5���X�8���t��Tk�r_��CN���ޛ��0u^����cѩW�{�=�^i�T�@������'��B.۩�p��%�r��Gf�4s��8'�M3��������|�Rx�J�E���Kz�v��X�;ȎipL�"���*H��N9drv{�b�:�Ӳ G�S��/$b"�r�?�HzYb�m�J����*��k�e��}zʮ��I϶��@F	P�ݘ��k>�p�%� $h�i�}��r:UBͩ�}�r���������%����ZF����`�A�Vs�*��͊m�h���9AO��+ö��l�s�O�6���SmD���T,�ù��qU�k��(�!��~*���³
/KEToyIz� ���ǬK�,�c�d���d�6/���m��"���5FnqgSAه��ēiX|��/����uc�%�
o�_|5}�M����_V�Y7�������6��I~H�S�n���Zp��W�mޯ��������A�;��&b�>O���k:A$�Ek�>�(���������4���v��sE��E)>���&x� �"��D�s����l\�r�E/d�in��3�l���z�e�?)�b�39�Zi!=��KÊ8TN\+IQ�۩A�I�9�F^>mz�*����*8�]�Hè�f�^
A������q"��6dՍg��s�j�X �]��UP��Q��<d!_qU�Y���`�_��ݣ��d,�� ��Ǽ d�w�7&0�ڋj�]<�K����#q��?oN.V�h�e���̤��t݌�h����[7����T�>��rih�M����l����m����t�t���������|ٽ���Ug�4B	;ut��g~�a��
ڍμ_�zq,�Z�7�"H�Շ\ާDx/ͪ"�*l�[��-B��-�.V�0��q�Kȣ_�ϣJ��WГH���ܩ	bvHl>aޠ�+��~[ñ��<�ә���7v�2%�3y�M�D���'�����@*���V�T�J�֋N�e��qɣ�M��*�3���! s������٩���娢C���p��cr-x�M�_�X^�n��� 4�����e�ג`�ܻFt��4��M~�՞��������qL�?�?z�5�/��i� �H�V�z�9�Y�����WI����E	��e��>l)u��ڰd��ı�.���k�{̀hB]mF�K�Z���J�L�Bx�0�0-n�Nr#�Q�=�X%$^4�<[W5~�ܭ�1`��ae�nc����Yj���̋����Y]���J��C����?��ˢK�:c>�LJ:g>�lTJTK�O!�ษ��G����>5z��jo~8.aRIY�ǸgU��$7�2��{3:�>:Q�L�ٞ�3nW�U�_:�ٕ+��k���8��l?���4��pp
�Y�m�_O���$t�g�	y�/��5��,�/�LM�A􂖧ֳ�P�����A{�0Z��kWEϬ�=&� 5m���|ğz\x�� ��|�}����J!�o��>����PC��5	�M�͈ͭXV�ޫI��`�2H�y�����wQlkJ����7��p���gu2x�Y�dj����xJ�f:���9�~w�K��f�.��.��3f6�"����"�j�`��@�wjX��}����<	W��r�/�$z��׾����zU�<�#)Oi��mǒ�� ����WG��ǫ}uM�o��\��cju�׉�8�v�{��F�Ek)Ry�e=��ȑ,]߾��{*���5����Mi�,<38I6b�M�Kϲ�f$Rn|�tAU�Rf�I(�0�5��0M�X�۷2b����� ���¤����,{�s�Ll௮�f�R}��N43�8-�g�r�̶zW���q�M�*8ܶ���f�!Gv���c"4����٫M}�7qKb����T M��ӕ浢��h���4�IUoS��s��=�Cӿ���q�\�������.�s�t"|{h��C`#���xW𿩫�8Q��L��1ZE�s�}���HX�J��i�=�h�B�XA�j�[�[�=Q����q�e�����C�I���g�a�6
y^�FRQE@P�A�J���ۜGcT|���������B�|6��h�f����C��sĲa�a���֧7R�;o�Af{��	� �Ozq���6��ud�j�.l�'c�X]�Bl����ą���c͉��d�-,���i����h+�����f�D|�{}�l�:W s�V3��*�*���7>���9|�Cɩ]�^�4��M��"d~1��0���|����[ ��[X1N��~4q�jm$�Hy~iT�P�{S�Y%��a�i>~dr%>���^�ڣ��'���`x̝��k�R/�D'̬�K�u�m]m�����T�BT���!��{�c�mT_椣��ܗ�]=�bC���e-������v`��a�W�o��=5� ��>������XM��ޛ)σ�g�e��&�y���0�}D�U>�<��U<Vh�~so?,(sW~w9�2��Yoc�UqNJu�}{�q0�cKN���ۧ������}�ߓy��	9�ϵfM܏�^C[e��_u���e)e��}�g�z�*���d7	�;���-|"��9sQ�RMl�m��ʲ�������ޛv�,
���ld����ї���U�	��y,��5�+�喣��QM�4��)���W�Sm�w\��6�����R��/K����u1٢�����G�}��+6	�+��N�~1rDA[�1���r\�>�S�lG\�|�劉C�͟Ր�[�H�d�`��i��#�	�z�z�I�U:"E��%zZ�I���y�����&�'��U��Z�=,��ηw�Ƒ� �o͓�Mp\��k��Bic�|D�/�6��ӑ28�#{���y�D��͞�ӻV���=m)��m]��̵g�M������� (@׿ �U�PS��	���nGI�Ly��>J5��Z~{�-���m�8xT{���c�,/L{���� �:%��)K��!��8-cw�~��ȑ����7�������Y����a���|���\��?�_>�ݧ���yt�#6c�G0�g�F�����(�Xy�rz�_�Ż�o���7o�S'���`wYUK˥ܺ���O��/���?�cy��%p�`�\#��������Z&�,iXm����]����țߔr�9�!/��	�á%���Nl<(C}8R���H��X9�Ty��+��wo��'&ॊĽ��͖�>�W�����7���|w�qYZ�.�GJw�0���C�
����-�oF'��N�Ƒ�E�	:)�Ϟ%�^�z��2E��ć��O~�M��o>+� +e��\:rnXP?<,���9�������d�k��6ɝ�䟺-1t��f$�x�B�I'Qr�w�$hO�~�\��h�86_u�����ɳʨuk'�o��ߝ8�4���jn�O�P���T�����|N�����rn�<�2ku^�i���G'ݼNI����5��]�A���.�Ў��Ք�;N��$}`�9'�B����S�� ��o�y�\����K��IO7��<t#<H�ԋ���UoY�x�ڐځX�x{�,x�}uu��O�%�:���.��}p|���7��?���P.�?Z�aA�jH����l~�|s�V�쳯�_�*O�Υ��\C�C���#��ƍk�G?y/ב1�ڐ�������_T������/?+/^�D��m�A��Q_f�[A�W�
G+ݐ&6���2,_���,@o��l�x����?������JEFz�f
��I��ֵ�Y��c���l�ײ��Mr��3���B��_ �RϩG\����q:���MX�s�SG�����a����t��k�q�t�%�!��8P�)�C�e�0e��AmC6n����Q^e����c7�.��銎�����L!�μ٦>g�h�+�8y�o��V�,,�ԛ,�lG��A]��u`����C޺����Z�Y'p��❣��pG������ʝ2f��Ω��x�N	���dޡ�MG�7�W����!�8=����7I��hP% XW�z�2�����?о�P�ٹ(n}������#�[O��6�O T{�P+��CYmZ�@�5@4�AU�A���fͬ,NN�T}V�߁��pzO��ɶ��ȣ<hw�y�]v�8�w��-/����2e�u�xy�ƕ�8�r�X��b��I�����?��|����ŰH��K�U0>����%n*� �v�!"����/�E1��<��F�t�A���|b	�o���Vd��j�E�ġ���E�:x R�<N���h�/}�E��^g���(+̯�yTX��&����a�W��_�Lܶ��� ��^s4D���̎�0I��8H�:/gˠ2��q���ayiO���H��	s7���'�塸n�H������8���8��p�+��=-�0|�=�*hq"�u|n��L�O�wQ���?�/:�*��M�tT�^]\��F@�7�s�����@�mj��{an����[g��8~M�T.L�gMצm��Ѽo�,�}�s�:�5����u��m��ܚ��NN������Q���pr$p�}�戱 �΍�4Z,��Y����,��(��s�����r�@�T9i�k�;,���{lkN�s���Ҁ��!��*F���7�-����{�罧�*/�Gi�^�1-ϒ��8�ʡ۩/�q����o]+�������,SL�@���/~�e���� �Y[���qଢ଼X;;ԇ��9�ư����U�(��o����w��7.���#e���̭�$��o�}X~���?��ay�l���0�	�tV$!��H���M[=���S�{1!�5j&��I�IQ��i���d��Ca䵳k9�>���R�*gϜ(�s��5A�ի���pŋ�[�_.~�]y����G}^��d���'����r_���D�a�-��L�K�v�i��6��g�[o�Q~�w���^�G�p>���~�ɭ����ᇟ��]�گS�����G��7M���;��C[��g1y1���R���Ӆ�N���z��r�{�ܽ]����j��8�Ϫ�Ө�/ͶGZ5���6�Y�no.���%{Z�֎�N	�/�^n�0~d��f����<��S(ݼ�ά��qT#�����'��d=
iw�4^�4u5p9�����ӹ�������U�\:�O�u�7��fd��2z�å�������K���h��H} �d�z�)�]�!j��!��\�<�\f�|nӪ�=;5����>�3�����������KO�!�\ ��7JY_�,�Kk������)��u���o˓'�U���z��]���F3������7o���O���-����vY�����w���~_n}�My�r� b;ۺ;��9�-���\�W��Ñ}}�����[De
��nn�����N��dR��J&(Q����U�)�� �Q�!|<ʾS���?��{ߵ;o:��h���celt�g�eaq]�$mr��{q���QO����'@ ��m����F��v��[�3��n��t��MvHGyyߴNY�]�$:?7_V�W�G�KR^�� �N���!qnv��F�ڎ6�U*�� ����a��}n�>�U��uV�!��np�T�up���g?(o���j���d�H'�n�4��6���ʈ/�v�:U�v�oA�I?>.�j�O�������,�;�a	8��	7�ӯ������`� k����=����\�>G���>����١�p孌����Eu`֐�3:h�����Cy�H>�Dd��rvȗ��nv�؏�Ǉϼ�]�%�F�i��ӖP��/��}�d���-�I|Е�2��U��4A��+���L� k�Z�[���A�Ed=|6_ֶK��eÐ�����N����d���� S E.v�8{H��I���K�U�uI(2&��W��@{���.ɛ���G7�p���V���������F�[Te���
�����n/���l��iy�m`i�M��k��? �k�&��v�� ?0�<5��vԛW��A�Ar�ס���:��^���2�YL�ѫ�V�V�T�y�����\����X�m�r��y��*�:|YD.mI����C�h:��[����T�u��[�
�|Q˭������?��-4<ka��H�Cf����c35m��?[u��6��.�g�n��
��|\qnol�G�������3j��	Px:4��_걽�/L�Q,��p����g)�;�9�X��p��մ<����m扣b�����iҷ��,<�R	� ��m=�6��Iٔ���W1���2���z-ۂ��y�ԟu}����2|��m�Z�͏&��u�Ml%Ϸ6���сr�ƅ�7���c���ǎ���80����n�������� k��/#Y�4�SI�:����vo�����_����g?y�\�t������Jy�r��{�G�N��_�/>�Cе�!/𦽛N}���j��3\��v���-ꚁ!�nԝ�iYYY�t�r�R�huh��Iw�FT�cmP��]�����,�v˱����7�����?'}�LM�����[+����?��|���B8�k:f��I��OL���G���7��S�ʶ��ރC�ճN�v��Sg�;o�Q���;���sq�鲰�[���n�O��/�?��/����E���ګ,u#����!h�Sj��8��4U��Y�W�tgr� fx��)���m����]q�`���AH�S��ȾN�<K�q ��&�XݰÏ|;��H�:���T��?��;C8�c��e� ���Y]uKo�%D:������rY^^.~�� ��<G���٪𮻽�k��G�]#���s'Ӳ�9apd�N��Ñ�,��Vgǡ��av̮�����ٲ��<�D7q�.�S4k)bK��K��A���1�R~���ى� _�EhRu��~l��[�7��G�k�q�@c�]�?����:R�%�g&˛o^'�z�\�v�u�%YV�����/ˣ�O˝��ʷw����+<+�s+T�%`��`��0�����r�̩[g�������fYZ^%�#�+��/�	H���#�C�ñ��SNA�/r�2�v�~3hdx��o����\����|��t��I�K�evq�,��Ć��͍Ͳ�.��D�[D�0�WN+��\��@F��ۺFF���]/:lRV������p��:QF�G�'��������<T�`<�f�5�~@��[9��c�v`NsC
"_�@z[��Po����@�'�L�700�+_4A�
����,����@i/r��[h��x6��env%�uu"�u�"<�i�C�(����2~d,�?�.�<8����ɥŕ������"���"�^�)+��`�s�$<緧��E/8�1<�j��߃�����ANv������zY[_ˌM�zc�������t9zt"�}vv��n=-^�1Fh8��\L��w{���@p��qض���K�E���lA�̆�޼	��Κ&�v�����ʀ��@w�+�g��f�I��r��F��C��5Ȋ�D�;�}eu�,.,H��NGl�=Ny�~ڠ.���`ቮ�j��4��v�!#=����这���A���/���`�&�t�U05��_~���da�>�/�D�=D�{(C�,G�2|Ke:=���J6 'Oⲁe�{� �� *�T�B��ml-�:���:���:~ְ��?�>,Ox�[Us-H�/�$~u��O�»���U8��.�>��k�N�x枃,���<�5o�E{Z4���W���>�L�+��oX��t�Ѧi�=|���4:�2�
�uSG��{�Z�#�+���<�^�Vxęt3�N���o]mFw>�J[�8k~�Y�=/
E�7x6]��W+�W�B'#����[�A�i�	.�۟�߇KrQ{���,���W�(!�H8�2�UT�6�PD9������ ��cf����N9Ig"q[if�Z���54�"q�
������s�W���I#����-�����(�������Cx<iu�Հ�)�*���*B����D�+O�ߑ�w�|�ʤW3x��8���iCsX���P�4�[�ҎW��S��#y�R��▧>�v�Ĭa@�˹s��O�{����o��N��#����ć��*�����	A�S���-���駭u���e�C�C3�$�sgf�����O�Z9�(�|�)��,�Ͽ�]~����O�-Ϟa�q]3�6���uع`0ֲ���#f3�I��թH�8�ϟ���-�W�G��k����8E@�!38~�˫���Z��8W���H�O~�n9u�xq�;j��j�����?��|��we~^�BGt�6�{�A 4�����׽�u��e�� l��.���25ӏs�[��̔+�.��W/�S��D��#_pz_�_��w���MY�ѴC�ssk�@h�DGZ��Q�m���5T:�5�
B� �~rtGr���*��G�VÀb~~� o1��t�4vz���v6GX���C�2Xu
���n���`�N����.Q���/�G'����p�>˄����)s�s/���jt���� �W�h�#��� ��_�C�"��"غS�\�,�(;_��.�˩Q��7<�_N���h��f�e�]$�ew�5Fena�<y��z	:��:�z���/�s.س�X����K:�uM.���*���C����?�� Kd�g���mG���u4Hنޮ�"�B�S�$Nԕ+�ʻ��,o�y���iu�pi~����^���[���+��?��_B�Mڣ\� 6�w��v�"wSӓ���cy������7�:���Z_]�+��D�Pm�@��+i���1h~��n�����du���!`���-��8ҫ����� k�iv���unv�<z� ��@�:�S��F��S+�k��hT����I�M�����qq~ Fy7Lp7qd2������g�ˋϳK���nh1;;O@��3��,���"�}���P������l���#��ɩr���9R&&G��a����M;�n��KW�׎�����FG��=��%�_,�/�M_}u�<��{�>�&&�����ip�¹r���2c����kD݁R|ɻۛ�Կ�n]�g,�����J� �zj���yy.��ч�J�2M��[������K���1�Y}}N�(�K��<|�0��d�t'O�*�/_�z�ɩ����\��Z��0����,_|}�|��Cp�?�Ӄ\ԥ�f����_������m���Փ*P�r���=G�7���[_Ь�{D���k�U���5�>�s�6:~��	���R���m�Y���OX�6<��Y��ם��'
���� y�9~	�΁[;�֗�v���X�t�Df�\>�\8	�Q��ή������|L���J��3���u$�^ �Ù}�i��\tO@�Cp���u���Z̽=#^Efuu���Og� ˼����@������4��I�H����8��R������+���͖��Wa%�
q�0��uY�u7g0����?�h�@�eg����)2�L�/��z�;�[���	��&�>�m*G�v������|�	l��NL��u�����K^�գʶ�Zv-��X�+���ִ*f�k���z���v�~83�u�G�ba������Y�a8y�<��w5O�/���3��60e�7�铓S| \5�O�XO� ,F�I+�����s�n���GUZ���� ��S�SiX�U��S8Z\���uZJ�<����񩳅�|M`�ƽ4��-������[�2X��i��_pgs|@[4��Uhã����|��O#�MzUu�m�^N�ᾀ^'����W�4���Qy��8ep�U��q����}��;�٣:бUv7WH���-�ݼ���7��;QE�/��o~����D_d͖�u�>�	�=����82���Q�+�Δ��w?+?���r��H����F��p������_�}A���ide��m�����wm�(�;�� ��Gǲu�;c�:��4�!G,t���H��a�Wpf6vp´Y�w	n�g��Ht=��F�4���ղ����RN��)?�ɻ��������X#~k��3�O��u��?*�ܺO��U]\�=u�23U�ѓu޻�Y%8:1V�];[�x�|9s�h9>1����N9��� ��޿��ܾ�,Ӧ%�'8qlp�7h�|l���&��3�	�G���թ_�]=[�〟��:u�8����Z�Z�G�8�$Q�&����R�s�~�s�>u��f��u�6t�"�d�4��4�k�EP������3'���7�����q.w���x=��ݯ?~\?��s��7��[������W��+Ν۷��{�����5��Lk;���m'xk3����A������ezj��:���]����%��㲆�����1�3v˽{��a?q�#��%���d��8YN't��Ә���{u���ի2�=A^�S'��SqV��)
���U�-{��:�c�ֿ��4ȂI	�]���5N�x����6�O~�f�|�l��s���WߕO~�y���˭����%��@i�,ꡎ�!��s
b���;�4Dn�l9�:Ӗ]?��H2��Q�%���&��/&&&���r��)h1��1�i+�i�n:V��������bY�DG�~�a�޻s�|��WyK	F�t. ��Q�E�vy����;솇��g f�:�3��'��c��s��:eR���m'k>GF��F�A2p��;��on����G.�-�x?���I�_�Ug��e�X)W.�+W�]�>'	X'p3���M��?��s?���`Ն:�ie��@��&G\�Z>����/~[��yT��%�@�v��`�Tp<�G s��������*3ǎж�&��"uH�N��G��Jp��#u��Oʭ[w�w����K�G潽udٝ)^����T����q�r�t�\ں��Z<x\�����矗�d����u3��7�E-�⽝Ͳ����'��7s����/~�;t����2��R@`)����F�LyY]��T�M�x�}s�2��ʀ�[}�O�mm��� K�Nr�=�i�N��r�\�P�c�����V���*�E�N���3�R�~�p�p5�e	�0Z^4�&�st� +��uM-2j�e�m���>1=Npu��q�r��H։�2�~���w�1��ey�l䮗5����E��)@Y �[*��m\榣8����� ���O�`c���*y8�:�6�ź"����2�S�$D&�j?N�Q���o�y5Xa[G^����qa�=����ք WF�N6���.t��"��|U�S���u���s�-[��n�i<�H�<���z�=os�rlK��Dy�:kYչ��M���C������Hb�^~w8��G��P�0�FP#Dm�;دo���_\��<�Ļ����;�eO��~�����R@�Ly��-�)~�{�6alyó��"9�5��w����ysXys&M�>g��������W�@=(�
S���ؚ�|�i;6�ц�����<�f����)��4x�tU�񯅳�Wp�1���k����Ӓ+	�ԍ#���	�ű�S=���:xVۘ&�Rj�l�R}}΍��:%L��"�?q�C��sc�pQث�֝��uR�ROK�^�i��>{2��D�^��2�#���&��p$GxF�5��n}Q�c �={����ǡ��ܐN�4X�t�S8�o'嘛L���l������X��'8��<z�J7q+�1���Ѱ��t^�v�������(��v�\$x�at��;w�tzE�	t�\�ഒ�ǎqΤ'|lt�ʻp6��p��P:��(��p��m`�]� ���tt�(���@��'O���w�;8��^��8uR'F�t���f�
��,��n��48{�/^<W�~�r� ��a"[a�ІG����:�N�]�}�Գ_�	��3mǅ��h�L���텶�����L���<y����孷.�g�:L[ul�ho?��d����Sq�*�'	lq���'fm�8t��=�֥���l����� �&0u�������,�u�\�z��95�F����&��^?j����SǲN�����9`={�g'	�&���p���~��w�����.0t'9� n�ca���ˉ�G��_+�߼Z�_�@�G)k4���9G	�ƀ��qp�	�ϝ9��?��M���n�Yu��)-�3��qF^X�Cf(�����M�;2��h�9ѻ��G�Ӊ̽�M���c�WeR�j����`'OgG�Ѐ�lw�Y-���](�Xkk��^�^G	�SN;�p��t��W��J�֔� �q���d��ˁ�n��nǑG?zꇑ_�~5���@ߙit������w�l7trD���<��щ��NL�t6}�/��������岼8GP�5�rD���3����th���Q�1xG�s�� �~bpK��(��0���n~w�$�訠:�v�Sp�>���[����/�l�z����7��w޾^^�20�.�O���f�H-�=)6���pG�ƀ�������/�_oF�;�E+K������<u�����+[ä���gOf���>>s$S�G\�V�U�� ���'eeZ�"8<
��L^<��m��UxuZ�������;����]*gN��C��Vn��np�'��u�^�|���_FFz��͉����ɱ�B����8�?|R�V�����U�2��톦u�D�D:i���)��F���F���;[�����08 ���\Zn�I�LmG޴�8����au�~��6ѓ�"ehiq����5����5+4m�5Uc��w�^��v��7	[����-���������=��6;D��yt=<�����2�nDE����A|���b���ey�|�,��/Q[�@]pV�}R���*�� K��X���A.H��h�T��@���]�܊�ܖ��dR.iZ´�uH�8�£Bu��|[%�:Hk�;[�����M]%���؊Sy��*� ��i��i����!���/�<�&鸷�)�6�U�WFH�ܶ u�*{�[b'�|.F�Wم���̦Kq����Wgu��.���0��;��4]���PF�8��)�SX���I���C~��Wq��0���--�i�S�꺆�����:�)7�\k�k�*�[Z+`\\�O�癏ȧB���8�yana�5�=���O0��ѵ�}�|�
�-��Z��8��`L�&?e�Gm;ď��ʫ>7�6��Օ�:�ee;Sq�#�|Tީ���5�b���_��<����y�K���Y��ͨ���|���xv�=��6Z^�gw���9��B��\>���{^�7�>3��uyZf�mO�;� �$N@�Ӷx�μ>�L �*V%<�NS/��vv��x��|��q������	,�Oˣ'Oʃ�/��GOʋ�semy��n�l/���D�� ��Y��z���N�؍��`��淴�]?}Y��xE���mw�.��LM������-����.JE'؞��~	�A���~�o��N�q� �,�'q$IՀ-�x9�L�'���MqRş<�����1;�3ﺀ1�����\y�܎=w�s�m�f�\����,��^�b9%Qzmo�W���U�38�.4vZ�����:6ݴ�3�%��)�.��?,���]=z�)<�M����t��Q���H���`�@���[o�^*./G&�éu���)q�FǇygY���7T��������;e]��<�SK=���YK .7	Zu��&p"�(����r���֡L���u$��z���Y;3�SM�l^��C��n��q��0G<u���e'����b�x�\�[�t�~�vz���0d���魘Ƒ�g�d�|�6�#�:L�i/2�Ƨp=�|280X�V�u3��E���2�i��n����Lt�HxQ#k�W2/骜�?R������ |�C�����;5� ٩r�0�k%�_X4`rp��.m@^{܆�鹽��N �n��)� ��f�<�-ph�99�ڄ������U'�M���~�����yv���"���u�v��Y��� ;�P�3�x���##�7�YW�g_�a�?��w��u�K�+;r,��*<\���|n?.-�Ⱥ�ć���`g�5��5G�m�A��#�	�ea��j�������K�3k�w_K�ѵ�g�~��ް 4u�=__���u4V�ĽκS�9���p��θ�A2�]f��,�{vn���8ڝ��g����3�:rp��r��f��x&��#@��z8Z���!;��Ĺ*v�J塿�74t����U8*첒u���C����O�k�`w�,� ����Η'�N�>o\*�.]��?5�#ش."
�{�KFk�W�ʓ�����'ea	�h{�);[b��[�Ȩ?�]��&�V9��ں��O���
�`7`r72�?#~dX����'�g�\��M}��ߨk]W��S�~e��G�R��p�1�nhdؙp��lul|n�Qzm�G��=.��A�P4z!�4v�h��z~� �$A�$<p$�i�K����z� �ɫ k���`݀�&�[P�,������ �C#���"l�D�Nwr3�۩�*O��hR!it�t�$�:��}�̂���o:��.	���_7�����:"�d�d���%z�%�,w_d�q*����^-
Ji�%Ad�h� �@Ķcu���IL���WA��_����Q��������.I*Cg�9x�v�J���%x&Sj���
ʄ9�.mR~���Y�"ӫPU�"i*����6��zZ�U�+]Z��N.���2���	���C��)퐦M�l�N�ֆ;��8*4���/ ��#c��+t�,ߐO��ն�^ǿ�՘i\��C��Xt;O\��\�;g��&�=[�e��N`��!\�5Mp������M���<�m (�T5���Q��6m�m������G9�s� _omP��T���7�|g�\�^�2���k;�\���$%��L [K{��̬/�X���ς����U�bͩ*�jv23�OI+>�������/2�.X�{y�:��w&�ȣ�C�`9M����l]��:Y��L:��y��og��ӥA�z�J9v�Ƥ�,/�����>)/g�`�}n�P^G��S����l�C� ~���� �G���;��F]/����9��dN���38�n��ڵr���L������׍l�����Zu�l�Bq��#�. �t�#8��l��jaa6A�ƫ"N��Z��U�W���1�gΜ��mɚ%����Jy1�P�4��IтC�tM�4ȂB���ݢm�S�S��z${h��Ȧ��N��Qr��[mg�u,.��b_}u+A~	.Ap�ʩ��>�a��m����zQ�����5�i��B���wA���{Tn��i0�-�)�����)E	���N�fu���.t�I�>��%�$�8�	�^'h~������'��D|�=���1Wλ�(��(<��W6�� #���Gp~I���G9�њ-/^J�l=����:vb�\�q� ��r�5x�@��m���9���I���^ڮC�:�[�ǥ� �>pq�ZGp`h0����
��Tdb�).�\!}=��z�;dp�+�sz�pp�I�m�N�>���t dt�lw���Μ�ߎ��:�n��M�!O��;w�q�����ab� x8R�(O��Fy�١�[-������(u��������K�˵+�7���>yl�D���9�l�ܼj`��L`�x�!�P�K�t�K]?����tW�!�#+�G�l�#�gN�`]�v� ��FqN{ph	��u�+\�$���&��>��t�L_���n��TX;���M=J�2	���ssea~.0�:q���ֵ��^�x�Z���A"�_d��Y�_�7_�ZZ\n�; �f���r�����Fy9��>}�]77��֋<��]cgG̳gO��rF��������_<w�LM:UV�A|���Q�^e� ŝW��%�WE�a��0v��	6A��i�d笛��H�?s
ڟ�z��O���g� zڑ1t�ɓ'������!;�����#"<�䮬m�g��{���ۜ���C���}��8��N+�^w���𻁖AG�?��y�yܴ�|�6�mK6�'��?h\P���e�{:�G键��#ʑ�U����v|��+E?�xy�N �%�W���7�E���9�"�bث��&#��wD(T��řN<������'f�"��Nt)�P�,��<�]&Ț%Ț�H��Eػ���y2I<N#r�3�
�ڲ:+5"��� ���T$�����Xb~�X�H�-n9��B�#[��%�J�֓@Dv�-#i���;a��n%GyQ��������e�Οe
�x�6��.	3@[̛���M��)��*�8�$�P�׀0��.Μ�չ�9h�
�Uq@ִ_��ob�Kj���lOb5]œ���:�ǫ�X�x�iܩd��}�/�)�D���e۫�_:�>w�%�4X)��Q�5Μ�!(l��6Op@>ӊ�,ٛQidy`l���%�.��,o~����x�~��
� 8���u��vԀ:�>e����8�Q��Ex��<1F/D�76ʮAil���4V6Y'���A�T�T�$]u4��0�~�/��7��Q����Ļ�T�
=U ���se~�)�G���N�3 �V,q��8��H/l��4-��:M�L:�-
�rt��������leQC���欼�s����λ6��h�u�t��;�&uJk��_�TOp�y_�B�W:�(x=��ۼKe�>1�xv(퓼n�kUX��t��|��:��y�\���Qk Y�ڣ�wd=�;jIS���ܧ]45��Է4)u
�#�g&���Х��n� ����?��_[]K�hbfz��>}�\�����r�����uѽN�Fj�,/.��y9�'f�@g��]0O�=]�H	��4V{�Y���M�lLr�ғA'� K�p���0�<u����r����Y����:]oi�n��������@���:C� Ў��aR"�N�k̺@\Pŧ���<nq�'���ly��E��������������5u�������~Wv��Y��."����}q�#t#��E4 y��q���P���h}c/S�i���\~S���a^������u�گ�!��;�d�k�o��f�t�L����s�cҢ����4�`u����Y��u軼��U'e5��$�#��{��^��G����i��v�	���1���-��o<�S�cȥGG7�c�<Z}a��#�XC'i����#$Z�t?y�x1K[6(S甄�~> ]�{�AV=��4��Z�iq� ������T�/"���z�N��\kX'���骓��G	�Fy��I�'��l~4whp��8~��r$g��I�^��'2����t�ȹ�I���qd�v�(�6)��l��� p�����.%�r���x�G���<�?~�$��EN��`9���$���=�5���C�0-��z��Lm�]BOlq+���`y�ojg�zJ[�{��t���S�H���s�����FX�2Ȓ�}�.��d�Lp���|��{ʵ���&�w�g��|Z�M��6��+�!��_��G�a5���0�F���k���Q��ַ�˯��;*�1O��R��37�9�O�k`���o��o^�&g	f&2��@W���dp��"���s���2��C��{�wj�
���E7P��P�C��T7����}������3����#7���;MЩ��﮻t �_[N���R�힮�}�r�ܹξ}P�d�����	�z�)��'u�<cǰe���i�!��7 ��N\Ƿ����^�ۙ6�v}�|ۋ�t�;���C��3��t��gIQ}%�j���ӦS���G��>�H�>$��A<D��{�:#Y<�:K��� ��̧�������4�c�n>4>���#Y��tv�<p$��\Yr��6�8�&��aC��cd�e��U���k�PP L� @�2��WgK't��ε�	�Bxn��0�(�vx�o��@Fbkl+�.��uP)W�%X?�4"Qd{�YG	���3C�k� ���Õy����B���V{�`dwF�h��!H���P%yZ��o�U�TG�����[�?�O\��uF�!6ޛ$�O2���l�����)LՎb�N�)���:��xKPJ����i8.�_^\�B �,Gj�'��(f����'��4��P &�yt��ϴN��S&0�~�c����7(1�k:�uu�=�W�`P�= -�.�1��cp&���߄�t��N�S<�åbI ��f
xJ/��Q9yR�t�����������N��W�� �v
�48�)��_�u�g�y����:'ټ�.�h�t���O:
���n�x%"�
�0f4�r"s�e�i��Yws�=Ҏ(�	�.��9sZ���/4�8r4<j=Qz�%���������,�>�R�`�ě;���q��2�Gʈ��r�W�!��o5�4�x�������Nv���|מ�G~O�U�O����D����rd'�,ո�cߩS'���W�E��1�Ņ�l�|��{�>A�;�՝��z2z�&h����^�q��)w�:�4�����Y�܉
�����lT�S�n^'qڜx����.��+����o�8�iC���� ������ݻq�t~�eJ�p=�N�����lP��s�����75p�c�s��|H�`Ze�@���'g�����8��u�tie;[$?����.Q��ұ=�!�X�W��@k���ґו���]u���n{iɄL�&;�t�YXX �}D{�o��[�/����Χ:��D^�)�L�t��0��8Ig�#P:AO)�~�}�^>��&:�8����ϭx-�(>�t#7���::�=�&��S�ޮ!x��[�ն:��H�k+^'��N�|t�٫�0�q�FY�!ӑ}�Sf��ӿ���рG���8�Ϟ=ˆ:on��-�Ǚra��#;{n5�[�݁�>�	����f"U��Zy�Y��U������:������L�qt��X���:=狠���?h 7@ȿx7m�(�pr�d����oe�:�6*󀦭��~K6d���g:-���=�ò����g�l{�ԓ��yl{}�]7\����z��f�6���!�v��#G���sA5�:s�TΓ�c33Y;u���Lu=C�>��Q��󜁯�dv	�P?g�� �䱙r���L���_���%���e�`�1�w��.���/��ݝ�ҷ�`��n�k��]��6�s/_�%�#Iv�i�]��
L��'p<K�5=5#�isD���^�~��������mt����u��{�">���8�urr<v��?������6z	���V���gݸq����k���3��lr��;w�ʳ��囯o��8=yGߎI�v������6wH�|��7壏~_>�s�n���?�	<���t�)�|�b�^�VΟs[�Q�^�]��2��7@�ޤN;�?~^���#\�����	^�@U��\B�7W�8]Y_% Z$�t����ų�O����1xБIy2Kp"�a
�����1v6�_���)������������v���h�3�� 9|�U^�Y�`�琯��w�_�w�}<������~�z����kY���{����*��v�Йl�p�/�A����X]�M��R�A��������c�eX�|�X��>�#�=����+j]NG_[�����R:#��� �d�ut���Q�##��n���T����˜n7��q���0�ȟ�r.��a[�;(�~�۞I��L��{���ͩ���8iu+Z SG_pTA�H	��^B:���罍��~ ��!�d	��j��q3 ������ ���g:J ��v��^G.t��Q>�0`�B�`���P�(�^�o>�)R`�N�܅Q?��5�tǖ��e�b�A�ԅ�r��>��on�������m �D6RnN�	/�c���F{�8�2.&uT �]_)+K(e�_�д���]I����O�ŹO���-�5���:Y#}���;wً���=)�~��&_C��Й�,�3�s������/�v݆�1�: |��i�C�&�^oO?��<.huB��!x
�y��RyD8�W廑Q�=��^�00P��될D�����Ac�^ozX�ݢ���9�N	Q\�6Q�,��hx���w��r��Bow�:J.~�-*W;���AՔ��iO�������)mo�Ҧ:�����ֆS(�zH��s��
���������`�UU�ɱ��J>G1�Mċ�W������)�!t�Np�έc��<�+bpU@8<���� ��̣�i�\Y�>�O8� ;��݉ąۘ��C�l�`������3|ե*��l�*xX��|8Mb�s���e�S���;�7��
8X.;\i�S����Lۀ&�p�����5箻�K~R����xbB�e���ڔt�۶q��&�Fn�)�y��Iz��I#�o� �����ܙKC3ȑ�<7�b�ܹ��<~�>߀&���ckNw���Q^ԁ�)�^_������p913VΜ�(�O-��ҭ}ݚ��Ç���enn6S�.a�_�f����r��29s��YV04G�ܽ��|������z��c��G82O)k�`��iy���Q�!C0ƶ�������\f_�`��`V���S�#z7����S�g�?S���,���lo��O�ʓ'8�؝5�#{5����YGv�]�Wh�����H��<}��,��o��%����';��]�~��q��w_�O��Un�}�ӷ��x�P$4��~񟐥�v8��Z(�>рk���t��^C��>��<x�s�c{�ν��ዲ8�Y�_��G�^�/>��|��oʭ���|Y_A��uoO�4�@ꡱ{�'��pj'A���,�m��'�ʵʛ�\/o�}���1�A���=���S柭��?�[~�����/��/�������[���]����q�^�'O���=�{�R}| W+h����	_ �����;o��s�\9�L�a/�q��s�f���]����rK���5��ww�g�}^>������$8^�e� ��:�N9��;-��ĩ�NM�׽і�!�?t)������g�_�1�����7jI��d�m�<�.P��(B^��!��ʓ�ɡ#exl�-ݽ�Jo�Q 'GP��Ogbx|��.G����T;ҋ���#�=�v�� ����N>��Ͳ���C����vn?h��E�L��cC�`݄^�~>#X�s���E�uy�G��,/������"��<N�,�;�d;	ֱs܏/G�ж��ϒώ�^�;�F�$Y1����+eq��k�aV���=�]~q�v�u�^�#����͉�Y���W;�ķ��v�w���mxy6<z���r�Ƶr��>� 'd���w���~�I��/���ei��C���X�>y�.~N���3G@�"��_}G ��=���~��(/_�797Jg��v�\�x�����ҥ�e��A�������NW�D~ܽqay�<��,)�k���'��}��4��i�� �l��x�ƮWG�9���U'!��8]�Sl� ������ezz:#Cj8Lo���+G!�N�]X+/���ťM��Ot�[��]��yp��|�)r��=���/|���T�e�`���i�����y�����Vjx*d��?I̑u}~g_�����U�� ��?BfT��)ԭo���n�����>����=q!��r$>�����Î�t�R�=Ϊ������ f]�"v럈����������ѱ1G��gG'	���R�,���bv�z�ܑ�����[Kʴp�����KF@p���Ec��iV���pO�*\� I՚���J�4��d��;8Ju�|$0�pI ���̣�����s͍H˨��ރ�3G���z�>���8�"eMT0k��N4S(��#c�W�����c-�#�Q�:�:�ٶ�X:�~� ���I/��<�׉����{�v^���k�T�:̊����"3;r!�l����3.�T�}0�۟:�)���3L-|�C{��]�j`�_W#����:��)�rYYù6�i�`�9�k`E�M�GA�W0`�ǅ�fP��V�n�-~ċp٫k����m�x���V�aϾ��a�Gb\X�e�ŰSp�+���ǐH#G����+�>����yΎ^9�P��5^���1��ڝ8��((�/o�̠�K���*Ѧ�
D>�'��y$ȲL�GFh�����
�<��wq�!k+�I�ԡb�yz�U�b�'|.<6k+n�!?Z�=vʰ�-�ΈA?�3�����1on�!���L�*�g�k�'��yv���U�.�� Hybu �����S9��lc�k�)���:�!`>�v�+���tI�Co�"��ya���jj�	�t`�He�����m���!^q�h�c'��yJ]�YV���'�	&���^�U��ػf&��	��t�(S�_׌� ������r���rlfڠ;��V�O�>�ax����#�w]عs��̱qʱ���t�b�<+_�m�/����Ɓy���r�x�b�@l�z1��p�!���qpD{�����H9"�����
�ȣ����AB�3��h��:�gG�Aޣ��a�@��z�#�0x�fʾzB��vZ���R�Q7��3dn'r�%����&�Ǧ2j60<���?n���'��{D.��v�u��r�x\� ;�r͈�t�o�K��+j��ndcey�=�:��y�Mڱ��^V�p�:�#��u����~F���<���Z���O��2:2
_��Cv2�knv6:�5 W�^(ׯ_��;�n3��E��p g��ۯ�O�%�җ�֭;����'8h�˷8vn����'����X�B�C#Ù�!]D���r�G��'O3ri/�S#�x��l��HN�q]Z\���%�}���q�m�ìG|D����_��ch����J�Led_F��@3���u��i�vP�{��f{x�w͡Jࢎ��W��z��VOܣ��U���֎���Mc ��N񹝸鍇_�h����)��%:�;ȊvJ>v��>���~��8vHD�غ�����}�;-J��eʁ��]o��ϣ�N���9-wz- O��]������evn<��������l���4G��<l��9���ZLN�`�����Kxx�,#�Yg�<���v�����9R977\w��t8�����r���r�;A��0�t�ɟ�M ,S�ի��h��#)n����́�Rsz����ezf��|<��G�CTrJ����	�o����sx�~oyi5�iNOV�=F�ݿ��<x��`�9�L|i��-g�8��ݽ�U��\�Ȁ#I�ex�>p[��u;�6�]�g/^�{�[�=(_~}�|��7�Swb��>�0kG�� ��v �}�ӻ;	PW���-�'��B��rd[33��e�6�rj ��?��Bȏ���<u�ӧ/��~���' ����苻w�^k� ��~{Q^mgu�!�Y�Ax�w�v�[�I�gD�3�=�-����
׸�'�3�����U��wf�Y��^噲��N�f]��l�7&�jg�#i[͈�>�2[er7��y.�-y\/m��Hg��+��b�� ���v�;��L�wDkr��wuw�Y/�d�f�AV��P+�4TKg�-�H?���V�u� �+��a�#��"�"�2��bC��$*f2�ߤ�CqLo0f��H�ßm��N�'��* �a�e=�
ru�ܐ֏Of7�����:��l�p�J���5����O��84SS:>
$�?y6^,��1��t���7N�;�34��*(�Td�@������� B&P�Yp�ju�%����5�0XPa:t���i����-b	;�~��>35]���2T��3�t���WZ�=�]{���P]t�4:�;M�)N)P!�����}JŻ�O�i��}�Y�C���]$m�a[2��ѯ�s�yub{{�8�k.Y�xqu.{n|�;�_O�rt�̧��y&�8u$�)����G�s��N�w���J�/o5B�h��3�gą����#��x����@�z��?���h��4����Q��q��Q��ɑE�H�%���Z�|Y�8B�"i�K3{�L�;������=9�D��|7GZ�v{����J�jl3%?������;yh2�Tg��Q����`^��6..�����7���AJ���I8B�g&����Qd �g�0����Ѩ��!�$;?��:�ʏ���N��}�Ϊ�6�4xrJ���.^����3�9���[[{/���N�����>|���"I�_9�9�	���83��9RF���҃��Ř�-�?�د��)���g����Nu�F�N��[�d���o\�q�?�t���C�GE����s8��c�q�g�M��5�}��n����8�_���p����\���p>~���Ӯ�pݖ83�r*l:��S:�_� ��g݌��65r�ȟ2��w�E7�8M�u�ı�K����m��;���>�^�r�Үn�qA|��&p��#��<�����}��]$�܄�1v�ױ�3����G���i�_��O?��{��U��QE��|Iĩ��?ڣ�ӐWXc�	w�Z[_ɹ�f��ѯ���^�q�\�`�ܖ�k�t� o^k��#���iQ��2��1Ο�5�?v|�\�x� �|9yl$x�"0�� ����~U���v�ҧ~.`y�`܀y�̻�`)��"�j�T\��r-�]�娟<���|�4?m�i�]�p50R�`����@�6��[���%�|�ӽ��)ڦ��∀�������jK�U�cc�|��;�qg�QG��-�R�}=����!��W���=Y���Uxί�K)��M��4>�>B��Y��*Ӫ�j��d������)��ٕ� gqq[Eb�)e�ઓ��w�Y�Ux�޵L@#�2+��٩�-��Y��]�Y�T�y\��g
O8��)�l��w]�Q`L��i�C'S��F����<ڽ�	rn#/�����7�u���wuDġ��+.�1K !���a�����*�`�R����}��V��	�r@~��`�@����_̺�	�\Αu٤����t�N��U[��	�����V3�usGC��/w}T�lm�anp�h]�ϒY-�. G�F~��OV�G� ��H�C�SSv~�v�N�M�j=����/�}���l�*��!E[-�{N~҃J�06g�]G�����r��kʸ�2�L���2�t���	��=t�����/���ʝ��c��}C �?>����w�
I l��j��S����
�o۩�ª��l�J�������K�cZ}se��ٱ�����i؎jE&u@9�_�T�COy�gԅ��>�Lԑ��z8s�����((�Yc�W�E9^�� ��|�2^0�V�TO�+pҞ��Q�����55���s��CA֓03�tM�_�_7��1b����E\�����8BR7�p��(<�� ��& �;=;4���"L�`��Cen���P�=��D��%��S�!����2w%��|D\&��&���8e�L�g��SG"j6��� mA�E�N��޸�ſ~ߡ��T�{r���v�ݑqN{���}���r�̙��GF���p9R��#=�#���~;�����X��Ӏ�m>]D�r]��y�:��z��j̝8::HY#8bG˕K��{����A����Uc��O��3Ǧ����S崻���0�|m�,�l�=:�8p�밻���:\�q��I��
�@:
%�2լߞ4iS��vz�8y�Ζ�5~_���{�̑a�6:A	f��w�50�)��(��1���Y�`���p��8O�v}	�>h[t�g���z\�x���,�z^Vr8������Sm�j���3�����i���`�]'N^�Gb����?�s��l:��љ��onu;�s�u��]|���`6�18;�A�GJ�����5<B �|����w�)�G��Y�NV��<r� ���ܹ���������,2�_7���p�s����O�����Y�p���tP����a�� ����҉�a�3��hL\$.�=����,\����Aw�x�����"p�h����Dh��q��o�(#T��`v��G��8��ݱ��]載��	�;}�`t�OO�FS�K@��եm�[�ѣeei)���F��b����Yv��|׍'9��#���G=�q�C���6�(��ɵ?NC��ޓ�4�ʫ|�b�a~��i���oʧ�|��ƞ�M�=�/f�Ή��N���NI�E0{�@��{w64�p���fl�`��鬪WU�n,$/��ԃG�ٳ����S)q6�C�����t�����8mM�O#�=�,�I'8	n�R�ȋ[u���Ny��wZ�<O@W�Q��5�+�����Ͼ*_|�5��
vK�i >D=M�7jo��?�Şف�Y�6�P�S(߷r�m��w�426����ŏ������4��	{�ʙ�/��h�kM�Kg�����N��؝��w��q��gO��ɑL�q�������W�K��M�B��-�#8�Ξ��J!Om\?0��)�����?E��Do��P^�&pz
��|� Gk/]tM��m�>/d��AuM_]��������]��35=U�a;Na�N��i��?�B�� ��u�R�w;�W�[ƾ��F���⪽�w}�3�%Mns/�$����T���j1e��=�o�tt̝��(����8�R�ܩ�n�ﮙ��:����%Pvڥ�/�ծ3%��5p��Qmg#��K6HX]!@A&�_l�q�Z?�_�Ee�e���B��:It�#��vz�w��'�r�q���k���B>���T��(Ҏt~{�;��o���8��5ОD��ݾA%.SF��1n��f<��g�e�op���V���}��&N�ՏsY��\�9�n�w;�l���0�?�:˩�|_N��2�sY��t�1��.�!�7�w:����H��kv�$`2����YU���::��nv.q��S[O����äz���[�u9뷾��;�+O�:�1���b��|�:Ft�<�D ��J�j ;��qD���Ԧ�������o��W��:�)l��MP�8Ŏ�~�������)Knv$ݾ�(ڷ�SGќ"}�t�f4�BwNtO�;�ʣ����k@�)Z�G�iD��`ɷҢ��:���0��(������ď�����Q5X�����[��ik�@~I���}��d�M���K H�m h6}w�,۔%?��!�kp�Ω1C��0G��w�� >�I�G�� �c���J���{���|Q>��V��d�̮c0�Q�Ώ�9�gD���ysmƙ-[kek��`��=�z1`=B�U`m�D
�h�P�I	�i3*��6B噴 $۵sc��o�!ړm��[�Q�����r�����W��0��xߛ�� ߩYN�q��;o�V��/��������L�x��qy�bz��t��`(8:����c#]��o���0���YCbtBZ���}���}֟�[ө��F�!�!͡�V��K�S<�D5�=M���"�Ĝ9y!�#_+++�������0d�e�hA�J��S�#�(�	�(ewf������G�ǩ��@��n1��a�Q���:
*.?��c�fG�[�X)��b^�O�vaW�@uҮ�G����Q(q^�ʡt�p�����kО^-�Q��ٶ�ťe�%
o�O��K�N6� ��s��\�V��ɓ�\�y�iiw��#���L���A�/�b�f3gܶt6�pǍ+0�n�1���=���;�r��� ��4��5�^��n>8T�\j�����������0�V� x�/�bR�xs$�)~��Ѓ d�h������3O<�&`h˞�l����k���IG��N�葉�:�Ϟ>�����S����r!?A;�Ng�My\`�=M�aU�z�g�'��GY9�V�Q�"U��{��1��|-��j�+S�-S"�w=��\���7�p&b���h�Z;G��E�?����������������Η�����,���/�ln���"3���޲���q�.]}8`]�h��נGg9�x��;7ʟ�ٻ��w_ǉ�h;��A���_�~�!��#�W�^*?��;��Y.^:��bD�"��_}T>��S���u�4�p�db���s�no��i��'���o�,?�ɻ�ʕ
�^��e�կ?.���,_{�E�앧L[�"=�� ��t9�Ly��1��뛯�,���)������>����_t�4�:��n�����m�~�v�~-&��`�6�1��K�ϗ�޸��N�;����\��߿_~���ƪ����vH�����Gm�L��7����t*�=����&!)��>X5ʶ3i���L0����W��|+�:�v|<o�6����ezf��:����Y;<V�������_�����GE�]g���Ӝo�u9:dum�<�Y���/��򻏾��Gn�)[&�'��ؑ���<��E�����r�ƕ|������铘��� w���w�d�ߋ�/�{g�����ߖ�߸��b��@�	*��S��u�����@�3,E@�	8G	С�v7�XW7@cğ9{�0Mzl=஀��~�q����3��a#�R�Οk��	�Ɏl5�0l��v�2<x�ܽ:=ۇ2���	Q~��y��ԯ�GvͭSϝ�b���\�v������G���Q\���ۦi���ʱ�S��h�:z���b��	�'_"�����(�ّ��I|�!l�L�p�T9wz�̸.�s7:�uQNכ3����c��`k [�>tFA:%]�=�]r���Z\'`;�z	�7�w�n�_��W���?���r���r���r���2s���8zw�|�|�ɧ�朻ځ�Q����(��?�ya[�7�6�]W�ZƇ���~���^��6=},�ʽ{���������y�F���S3��'*��ך�<���溣k��'�զr�C���J���(֣L]~��%��}�+<��p�Q�(
����iCϜ:Z��߽[��^�t<vB�r����ǟ�����n�{W� ���I�[dg������c�L������o������r� N����vy��/����m��o?�~���י�ؚS�_�Y��{o�s����|~i=3��s?�̾��6�3K�]�q�j�.i�2��ʔ4�A�|�l��G��ř>��bG��R0�#�1���Q:��ZV9�C�b��[9�J_U����m�Q[�jL��ʢ�n�f���	��K�0���i�f0� �?��p�S�����V����Ҁt^�����cr��U+�*�O�`�3>�_N�)�.�.�q�\�f_;���|%Ț��>��ny�ן��~�my� k`{p�1Y�;B5�P�=�4�������j�� C.���`��he�;�:�A���� Dk!�!��f���,����"���(�M��L��m]��}����<���Hl,�m�-� ����C�^9A���[o������8\����kD�*7GdTNuF�2�`�0��;Ѹ�ZWy>�<C�N+p}���JH�ϠL����O���e���U8��[�Ѻy�}tn|p�t�s�c�Թ�S��OO��u��JGOG&5f3����YNm�A=	�ܙ�ު�%迒��&��]x(�ێ�JЩAY�~�s'��J� F�*(���N�rJ������y�	�Bw�Y�i�$G�K5 ����("ʑ�Pܒڹ�~�f5S���0��y� ƞq���	wRtj�J� ��UԮ'�bif`�?iq�47����4�쎆cC���F�Ky���%�18���U��0u��'W�+(/��	�"R���D
��08�1��/��^�2R��?�/*!�0���u�	Fm�m�m�eue/SA�=����������N�@ցC|&H&��<��t���sq���f������$�w�tvנ��-3SU�@*}�k�%��� �;�VEN��G|�l�(�^Tvų��T��L������#2N�tM����A�/������8��ԣå>u�4��ߔ��?-7^;Y��KO��;�Y�������k��ڪ���������9�βݱ�"MV�?A���ြS~�1�x�lt���B�{����w�����	�~F@v�+о���G8����	0^<��l�0�8c�ow�S��n�#���v�긟���r��e��qx��-�H|V��~Y>��+��Y����FZ(�N)s�����~#��v����w�� '����?/���g��;h���Ȼ!�~�Sj�PH� ggu�����S�3�N8\+o����Uh0�iN��=,���~��mt��@=��m���=��t٣������㨣W��u � ���$�F�{鈍zҩ؎�_��-���;�9:agd�@W��]���ä�kB>�=�����M����«Y�g?*�?�oDO�� ��O�,����_>��g�`	���>vڎ�Mt�;�eJ,���+��A��{oC��ֹ҇��0� m��	~���[w��A�dy����>;[2B}����]�Ӻ��~FŲ�Փ��k�M�d� 'H�!���3�0I��n��Ï�?�����o�á6��!h��o�,�c-t�A��1�� ��E����l	� ��S�9p��=P�b��:`��`Š�Q��8�NO��X+��/���R�y��SX��.�9z��d96=].�p���W��\X._~�u��7�.w���+�/GTϜ<��4'�;b��s�s��#���'i�No�{LS��Q���<�3��n8���~���)���W�$x���v���Ε��|�\�r9�B�C���Ͼ ���ܾ{7�5G�\�.�w����z��#��mxpsm�\Ɔz�_��Oʿ�?)o�u^;�~�*��/�_}�A֯�̾X��u-���(�N�;����˟��W/b��^��e�_��Ns��T��O C]���G������
�?,���ߔ~�qqM��p��>�4�&HV�A�?��7���������5��}�����D�/��myH𶵃/�맄��3�� 7Q�Z}k��ѣ�GM����Y���'ꇥ�W�˯?����?~�>�M�M�e���+W���~��wʍ붛�}�4�ٹ�lG��ǟ�_�i�����}�凅�G�-�{��l;.2�O���W�������'�l�~����ܫ6�S�m����'��J}ByN)�Y�і_� }y��4��*�՟�ttҒ%�����z�k��9�#\��w�g+<�6��tn�d�����M5f�9�A�0�a;62����r����7���玕�'��1g(�w�w��K�;_�=z^�0e�`>F"�����%���ػ���ei��3�	W�X.9y%���ۛ�Ek ��l�"��W��kEW��kK�68�6=BU�:jU{�`�����:�����\�+��P�l�@�5E��$����x9�T��m��Ӊ\{�:��#~��lә��.#~ΩZ�N�2@%�ʖՃ]���Ȓ_��8����2��P��S�4fGG�ĄS�,[V�HG,�`���5=5��X������D�u=�y�}I ���T>�e�-��9Lp���ͲW��\�>���ǩg�p����\�n;ăC�Nw�cxNtz��N�A�S�\k��&�q9�ѮI�?���V��c��� NApZ�1�=��|�u_N9����)W�L�۫l�Vw��QqZ�e;�pf��V�x��2�����g��S�����LmsZ�$�5���%��W�a�uw�����Ŭ������)�pJ$4�ݼw�H;S@�ad��#�3h��&�!r*�����̯3��'w[;BZq�z�>�<�v�S��#��
�m���<ly�Jcc�l �`�x��͝,���cGʱ���1��Ld]P֟�{�t��j~G t6	�{�qhw�2�N�<�l����Ɯ�%쁴����N/��v��MO;�zÓ���ظ��.����S`GŃ��#K޷W�<�vcCerb$�Y�Rwr�G�e.�;�����N���������A���mn`L7H����d���#:M���I���1�^Z#oW�`ݼq� �fFN#�C�{t�)����e��K�]�KyO����S�!G��~U;ug��~�Ι��(u3�E���p�\ݻ�F3��ѡ��f�����?J���ؿ�܅���1�Y��V(~�����Р�t�����ŕ���Kk8�N���U��|S"z@�Q%��9���{h���Q=z��i�X�\��>��W�x����h�<qra!�ĳ�0E��NP:�G{��k;|�ͅG7ח���:r�_.��w�z'����kר�l9s�:p:�S�u���#vR�s�[�]��R�dZ,�X������Y��������3�؛i��qR7�?���۲~����e�ږ~�F�2Wl�������U�j� �D�t�LF�zx� �`F�����{8���� 6�\�(n��Ў}�O�i��P�Mtg��O �ȑ�<Ќ�����q��p�q�)C��)��ё]eqq1m��9훇g�}�FT;�����l�;?DLN�U;��}��{���#߅��U�۸Wn����dw?n�d/,�e����l�,�Ļ8�Nv�)'�Kn���3�I;m�Y��Bv ��f��2�n� @{�U��;3�m@/��]�>;�ҹI~�,�������G�B�#�:Ե��L��k��cNv�tE)}i���Jq�GO��s}Δu�Lݚ�ϼ�#���TA�c- ǎ� �x=	�����lGo���p;�ک�N'wʷ��W�]�L�[�'�C�=x���>��)�o�\;()���|�G���<�ѩOc�!�Z�3��C��Y�Kz:����f;Cő0u�3j��'���\+��`;��[ڌ3����1�@X�N��;�a�n6�YX\��Ki�����d�wD���Э�n\-7�],'���<�/�s
�˫kn� �������l��n�-�~N��6�e~����Xz���O~�^�fY�k���Z�h���NM (�/�ā�@Vf�qo`��qt���L�3`��*�����LУ�s�)�?���<�&��-Kޖ�kPXˑ�Ų;0v��'p����Ά�֐!J�a����XR-/��B����ڱ�!�*�qF�RW�⿌�ק���������v����w���� �>
���ٲ���;�1"�H�z���\����F�4L�gD% "dg=��8kУ�����%V��zJ�R��m��1VQ�y�3���5�=���(��H� ���%��%�� n��<(|{K4~�5k50W.��W��\R�L!lug={�5:����t���u㊆X��i�:������s����{K�PY(@:����;��a��aP)��:6��m�(���^�^� ~���+������\/���:���D:�8��t����P�Ʀ:�:��g g�ie��(V�T4Re0����SOG]�[ �![�	�`o�=v���C�+�ψ�T�o�t�&4���f��t�B�@�m?iŷg�x�X믰�;�E�Y����\󥃮��:��-C�z��)픋�iÃD~��H8`8���;�C���>�s�D졜�]h��i�:��JZ���;�Սl��m0��1u���S�@�hd�
�oҁ��[32i������r�)�����·�N��n�w*�VfO�D-�d,b�t
{z����h.{�C��buP��1z������no���V��~��:�!?#ZR��nyт�cz�#�խ����!`@���08T�\��t�wz���������WN�8���Y.^:�3".�G��\���YN��Jp`À�]$�By{w5A���y��k��?~����լ�'ش�8ξ\*w��W����Y�ĺ!��K�5��A��/Aa����u8���V~O��fwt47b�T.4T��7�8�q��%>N����LJ�}��Z�L���k��х�&�:�ng�k7�d�#��:�!�������mZ,[k[�A��N`�S��s�ܸ��o���B�|�-�/�/�q�.���G�# �]`�g�����\�SJ�k'L�(���v��ʏM���o�GƯ^:[~�����^y��7�yh#��R��*�Y��2�P�^ʓO2ҫ���9
I�~�T�����<}�N`O2�Վ(��u��5�\��s%�Y��B�N=|���+S[�\�t��CZm�r���ZK���g�u��F`���1�Ti��:����t8ݼy���+�Iw
�62z[]���~�V������vp�ϟ������@2-�Fw��3��!�WWw���2����<�۰FN
�Y}����:Q�
#��������Iۜꄃ��L]oh�͓�\�`Ge*յ~
%�oA�+W�g�ʖ0K��y�I������t9s� �)�ΤqV��~��EY^Z�=��>��q����[t68T�����keYE���h�N�m���i�ڼ���v�=����/a][�J�x����4p�g�����KE3�1��wt��%t���F��-��޾#��A ʕG	�u��r&����̻z��u�\�|���HxP��3ɵ�~����` ��(vHN��G��O{�~�pWVu�r}H��#�a������zE�����~v,n�Ѿ9ڶ
lN-�g������s�UD��c����cдݍ6\��k���P��3�.^(o�������΀X����Vv*t��Y�A��hu�ٳ'��n��rD�L?�.�N���n)��7���.�b8��7ؔ��73o��"(#=����6��T/x8�Ù9��<�SG�x� )gu֍vV����+H/��H�r��z?q@j�V�fG����ȗ����� Q_�z��Y�-O_ĺZŠ/׎�Y�O��օ.�>֥�N�@
�[۬��S,��W>��p��A֩��)S�]��[�������\��ȍ/�H��Ux�8mp�,��A?��p��,�ёq��A�����9��Pd�+���)���<̓�l�{�1O3��W�i�`�pɜq�e�U��_So	av���q��S&s���FݠO#�S{�n^;_�x�Zz�p@gX�Рj���(�V�,�ke�@��Qw��w?B��e-~h"W��ھ�C�n� @���ٳ�(�4�e��1����:���[�u:-�!}?4��tl����e��i�h��7�Y^�J/�����S&��tH��5���qꔛj`vP���ҲGL��#�pJ^vs���Q#Mz0
N��4�� �;����<0t��	F�H�G��tM�o���������u�];����r�챱��6P��Kk��1�@��.�##Y(c{�tN��r�t6��`@�"��&����A4�C�8s�<Z�R�Au�^�IO�[�o��A�UʐGi����I�gڥ~�*�*����Pi�&�5�w�H�4�ԣl{��@f[�/၅�A�j�2���H�ݰ�{{�!S��k�����*�|��7y��կ����a�\G�]�3 M�L�o�����N�}wjۅ��O!�r���B{%Z�!�E^P��z�.b�SC��{q�\p���L�A>����,����N��L��M��"y��lh���c8 	�N�'�W���Ӟ#�s4��������u�ܤM
�2��Լ���)�o�sr;>��	}����Z�����o����;w����k	�t �SD��0�2�����.(���M��F��ER"��_8��0_��r��\�D��*�~���kQ��� �e�`=�ǎM���/��	B�CbE��k��
?����ӗek}�NkQ��?�6`��5�6��N:�ʋ�\>&;�dNN`_(C���A&׳�Ɲ;��=A�����	���x�P�tܻ^�[zΝ.?~��g?�Q��;;Y�E�k���zKƬZ�ʒ�i��'�� ����]��YwF�^ީ.��S�����}����;8�����iM�EZ?֫Nw����π����i�� ��hgv����s���s?D��k�ݹw�NY\ZȬ���q�j����)7U?�l��Mݫ�0�[`W��No:��2�猼�';�ɍ2ו��l����|֚Ŗ��FG�?ur��o�O�*���ÿ=*�mF!�����~ub�xV�����BG׀��~7qe��A����6�����$<h���]�|�,�ۏ�:�ct����q[c��H^y�!�*Ǧ��ف#Yv��s�Kr���V���ŋ�˔������"�I�ʑ6A�U����:�h�p�C��[�~��H���ꯋ%�BP3AY��c�:��#��"�+����� _V�/��p��8w��;'O��)o�~�ܼ~��>=��O�SN�_%�>�~���)�ʙκeS�����V�0����1x��Eϑ�S��V�+\��dԒ���<�lf��c��H>�7�eЏ����K�{,:��ю>:��i�+.�F��s��-r�Vb笇s��؉�r�����[���i�u�PtX*���A�uvO��={��m}P7B:2N�����ʎ��3��wf�[X��؁�˩ش�z|	�6PfH���5 ���>:���{�_	8@�:ϩ���Y�[�ѳ���V�í~^����Y�;�'�)���	|VLl�|Z;�� ����꠆���ڷWq��1�k��~��%�#�nt�>�?;eٲ�;�+�'�^�Vod�D[�U�T��:�u
{791Z&G�K�A���;]p� ��.Xw�r3���~��{x�H��*��AU��Y���� k#B�_	J92����)aD�2�錘�B[g�V��42C`�SC_ג4=��)��W�aMl=�-3���ϑ%�!]��{�tD�����PN�qj�M��r�]�=�~$X��Q��s�#0mq1e���1�����g!.�����>��]�g��pq����I�kV��RGAT����1�=�Ϟ��9�㎫��x�k�苣%�T� u�q����]���~k�62�fϋS\�ˈ�����\h:�)D.5ؔ�*@���:�o[%�=}:f�Rf��Ƽ�;������-Rw����\�D�&�Ǒ�l��Sq%��!r[=�u�n�Zu����5b� (5����}I��Ϟ=�~_�6l�k����Q��G���at8��Nq���=��A�SF��S�:	&^�#�a �&爻HZea��i{�Mz:"��v+Y��9�y�ګ�9�����}�2��6m����-x�28ݍN��F�T٣�#_�O�C�ʗ�u��Cڶ�L� ��k����P���ke���+����]�G蕧O	p��קO^�j������y�� � B���ى~���q���l9���hd�8��r��:9�ޤ\�VΡ=��r��'�5���*S���i�){�^�8�%Nt����z0��{_ʶ�s/_f:��@��.'��.S�N�ё�E��$���������8(�0�\HO�涛g���Ǒ9��7�pa�F4� �c�^�[B�>-�o���z���k�w�(�0�N=5(�7RD�P�3��4�9�2��K�u�P�Di\u�Պ�B��)�,NA�{,�
�(R��?�,���Ӌt��i'�1X�����T��#��xQ��^�r��F����'ș�t]��'�-N�=���S��*��:�ڦ�,�8��܉����3q>��Q:�	zh�L��m��!��2ܐ��,�f�U��H��:Dѷ޼Y���~�멓Gi�q�t\̫]����Q,�&��x�����|��k�@�;Nm4/M����>z�'q��NB۷�ػ˩:'N2稲:�ɣ�ٖY��*�4�ыt5 R��{!��^q�݅󧲉�����S@���/��2A��8Ϝ=]Β�i���|��
m�Y���8�t�ێg%��@&ww��vF5��8��FK�Wu����=	�^���|�2������Y'��� �>+���&��	�y��ϤV}��̳����ͳ��&�n�LA׹��O���4�m��,��zX=�]K�h���B$�A�O�g�W�ߝL7t3����:��V6��_d����]*����LyW�B�-xkqi)��>�t�ǎ��ב�v0;�k���{�\<�^�C�)�����|���n����˗��K�k��n���/�ӱ�	D���BQn�>�t��V?N��rF.�c{��߸Y.]:��)�-i�����)ܱ�|܂�o2z���u'�Օ���.�:������΋��k�jǠ"�F�7����C;?�{)���t�De�2n��J�K�a���k7���޺I�H��Zg����'��ofܸ���F!���@�r?�`���kW��v�(0*6���7�v�톮������G����3gNd6���<+�J����v�6B~9�ǳZ�r}f�a}�~�A|!�i��(g:�	�חKz�L�s��,�V`��%r�)�����&�h�\[/��1�o�7���їH�;�ޮ��SB�;®���Y�tX�/ub�\N��n�m��wr3}]?�n�&��'���kYs?��5kc˶���
�Z.�ûY�C.K9ul2A��a�C.�������w~��]P��?��+�e�Ez ��U����*n�q����HxO�'#O4L%�ƃ4m�`�H��.I��H&jdjëa��G������(��y�.j�
�⇸"WD�DS���YS�� ������mz$W�&h��@�J�f��d�X��k��om��T��|��&YԩZ Bk�����Ȥ��j�_wǎi����>D9*��(&�����ﴙɑ�������z�� � t�![�Ƴ��۝��r��WK��k��R����]�Z���moV7�
��Aݷ1=|1=�0�ֶ�@�{:�*�1N0B���G����m5�5����8Dm�/u���<�(����w�g�~l��Pv�ٓd;�Tm�6h����Cخb�<o_|� '���r	c���1HFG�A�e7��>
���?v��G��X�DP�p�<2�06���}ee;ӭt=��;w�/0v�WuhYଳk9*����cO��x�@H�A1;�2��*p����_}~�}��W1����1�R8rr<��Ci�֞��X�ܹw/�>x���Ġބ!���������0��6m����\u&ƫeЎm�33�R�"�����˗k��]�GN�6]�S=n���c�d��SQ|��j��� Ϟ20���R�����Q�y��7�ﴯ��&[�I���h;B�[�Aȳ9ֲ��J�}�Q��?o������%F0|:�<21�m;��0x�z����_/ڗ��)8��xt��)�i8������R����)c
�I�M;�nw��U��uV�{��&^�.�����f���WG�t�WuXwp\�1�<�f�HX�'����m�����HG94v��e�-=��s��v�]Є��,S�;�@�|�j|.Q����A�Ҡ΁Q�^�ȓk��A�Ԛ
E�#֮/�s`Z��q������o>������ ��{���\��+������,Ҿ��y���2�`���|?�����:�y��uqC�;M���ΑU.��BY�!���qF�p��Ϸ�>x�}���q$�8j��)E���ണ�?<Lv��K/L����r�����KG��<땺����F�SBG�9���L�n^� 9�c�]^�G��ŋ�
a::<l�o;]N�t$�3ײ�<:l����8�E��)�N#�������~�����pz����C�� }�j���Tlb,����Bkү#��.8"��f=M^����X��H|�A�����5��r��O>i�޼]��W����vgc#;l.ã�����k���$|5]R7�o�v$�c�:�['�u����#Lc\x��S��ϿȮ���y�b?��������Q'g�y��&�x��}}����#������׎./+�Ww��ݶ�b�-=A�A��%O�I�c�I{�����-<�14�j�Ҡ���0I�~A����F�q���:�O�D���/�h;>�rWK��~�ƅ��O����~��ÛU�ٱ�PY�M~�K��
�st�ƽp�r����)��硫�Yg���v�:"ae��:�'�1���=�r�M��b��XO;����[����/�w��'"���<��q|��M�������v���6����7�e�r���#}��{��3.^���}�Qⷛ�|jS�Qr�Y�q�*#��	ڐ:fζ�@�G����h��T��������9e�#\���'�w<�=���}�Y������ވu�������y����ѫ��z�s�P�:[��2�d�4���������4�svz�Mg�r������������ۿ�S����qd^G�����mqn�ͻ���4E���ah���33:��mc{	{s���ؾ���v��\�wMr[����o���ᡇ9?~����.!Ko\��\���a�K�v�N��W.?�Np�N����������d�nS��^��,7���ݼf
�f�rpg�Pc�K��衃&vT*��	�:�ng�V��*���u�Î=g+`s���3�L�;GG}�Û�G�`a��N�3��(�i���ґr0'N:Dg�飦w��S[)���N��9lG�Ι�8�=73G��A��XsƉ��|�i�|E���齞W�t�K��8�:[�ԗ�z�d�֚,�m�1tw�v�d��.�X�F�̫�y����XIǞ��4R��M/�C|��@E���t�NW���#F�
:�W'�9�z�~��M�e���!;	�����c��oC8�E��c�8�|A���Cu$D���5:�(�҅���wnf�~���=Ơס��_������>O/�^�Z��M��JeE�BD�{�ݡ��sp���!/�8���?�v;]w|r�������̃6o���ͩ\�޼�p��Y�۷��6�̝F�h��� 1P�I�4��)��ç9O���'qwW�Q��mn����g,^-�d��Ν�����h�>����661,���a��i�����������ּ�m�O�]�pz����#wa���2���#��#�0������?��1���)��)b{rt m�ۯ���k�=ꦱ'��-���g��K'|n�o:a��	�N��=p�T�7wM�#�NMr�k���� �@�P7{��{G؃�H@�ꁒ+�����򛻩�#���~�όJ��>���{(��rܼ�q�����1����)�,k8���W��ha<�����_�����N�S�i&/��g��߳�^_u�Nq��n�,M;Uѭ�=�	��l�j-��!Λd�u����us���8��_����[�n�E[z����x�/�WK~;
�rG=<�-�ݬ�F,8t
�K|�Ӭ���kϕ�'eT!n�J㘲V����4ݼ{pY=�n2�ܹ��yw����LQ6����i���k�֭��G�q���~Ҿ���9�m����+�Ti5b�C�#.�}����}p��#�y���Z;:n/-�d�������q$\�xX�Ϊ
��]v*�m;��J݊��⼽߾�=w�Bi�ކ��?�ȵ�4
C���;�;�%��g>�;ʹf�݁��N,w�|��5��~{��/�����^�ꍌ)o;���T��C1�1N��n6��+�8�CM��8�߹]G�q���ƨ��u��:Z���5; ]�9�~�������L�
(�e�i0��4i�܃��<}�S�:�����a�4�2�@>TY��ᣇ�6�>���G�*�U6��@��j�^zF�#��<�۵6�����I88�=0nwi��ҺK�ƽ�\h0/]ڻl��F�[s?�f�Ӟ�wg�ƶFdP�SoaV&:Z莡�iS�e>��(#ln�s�?n.���e�j:v��[no�W��.�t�ԣ��?ϝ⽶֜~����[+���uI+���x�&��9���$��z�O�-���^�dzơ�n��INQ���e�y��f�Ws�=���ܱӎa7D����{��࣏��[���#�n:ၵ�����ɍ�C�sksi���t��Ny�J�7;D��s�rzXn[��Ŗ����ǽ�ŗ_�ϐ����m�vX�|w��:U}g{����E�ׯ��8y�-i��<�r
�kjqy��E�g�ex�ы);�q}�_]��bnF�FbnV�9���Δ����]��c>f��#��ʯά��q�F����zn@���o�Cs/��Y�,��uÎl��܄���x/C�[1�ȩM���=t�:<lGÏ���A��qSN�~]����L:pt�m�v���C�Ud�s�Ğ|�ݛ8M3�X�c��e��X�ti�Mt�����q��y��q=�j� ~�o����Q��=~���}��q:�8y���u�H�9�/���OF܁��.�fMΞ?n�e���"]6�@I9=O�]Y���#޵��p�a�� ��_��q�pl��#�`٦��O �L��8`3_���HK�pইC@�_z�)�&6�(�x�F��?1asc�Zu�(�	�-�&�l�e�i���i�C���u�?����q�4�0�d��}%R�ƛ��ho�#Y��\!�bA�����Ѣ٣$�dA:E"�F�t2�W*b \/W9�7��J�E���)�Q��hY�Ya+� �2=����WH�	���(�AE�i�ۆ��<K�mdδuǩ[����0���ܺq������N�=/0<Q�7��,�j�Li̯�XA�x�#������(����Q��8N�s��N�s��5X��`�0��|���\cc�3�Huݕ�5��Uցy�pr�CE�B#H�X'A�������\F�Re��L��.W�6�s�u�<g�10k��y?z�"�8�38�`����F�������}�+�t�ě�u{<:=�n�R��S�]��tG�<������"{j,��r�7��)h�yB:�~�ݩ�:p�v�3��s?Ne�}}[J~�0�\��=��k��U����`>:�/m+�����(M�f��o��{w1�:M�E��#k�ۆ:%봏STV:;
�{wݵG��Q��N�#��m��.��V��r�bׇ��x�pK�~�ӥ����iR��=�N*�Ɲ���ә��;8�ޥ��3�������6�隞��U���TR��������Nb*E�*2{�u�2�g��3�:C/5ؠ�n��)�Ғt�<�N������=��w�N�q׶{w�dT��A�l��/�oo�ӛQ��hc�j�țwp��M�G�k�F�T�{�s�U8�2e���TQR<;]��GN|�wj�6\E�̩8uf�(,G�t�?�����_��}����[�.h�_qw�n�9��j\j8(G�{Sd:�:�
6;r��XW7A��эa0�޺y9���8:�"�.�B���B����ԑ����Zץ���Y�^��n��a��&k������]y7�P�9ʬ"Q�#ڣ/���*;�}95��g\�B9;D^����rZLj8�ӣ'�Q��)�uF�a	�(������e���[8�c<��Վv Z��K��)<��7��7�F:YB�P6��N���t�:��J3N4'{M�r:}�(���g�a���8���z��?(:O�lЮ:-�u��8F��C�}�Nij<�OwG��
���vq��Wu�F�]r��:�َQw}�q�F�� ���M�Pw�̽���>��w$��NK�W]h�ө]s��K�|���G�R���/�l_߾}�����"εK �2x�Do��N��M�Q�O��)�9#�o_�q��{'�iĻ�7;,~��lx077��b��X��<��ez��Ⱥ��8α�Y�Y�MһC��>t���ۅ�b��<������b�R9����sZ���h���Ҫ��ΐ����O|j[im���@�O�� ߿�����}�b)�!�ԋ��.���>v�b������Ѻ@pd#1�����O:���ώ4�uy�����j�i�zص;�J���Koߺ����-rs6�f76�1O���iK�).?��g7�q����q^=T޳�h3�R�w��
��:$\{��L����+ŵF�а;���u����w�_�����?n�x+t	dzxA���8gm�NO�^��C�ݤĥ	�~;k`kk�m ��ۻo�j��v�v�Rs��t`V�:�>Y�]y�����W�� ����5Qx����Y��>v�:��
�>���j����r]#�O9� 9��&��P��n�ȕ��ʶ�qtP�q4�F�,�@����F�� p�]�z'iG�Qw��F�V�n��Ծ>:ɲ�S8�H�|u������)ޙ���d~:���#e�ĭ�*����:�r���~�G8<X�8���2Ik�����8Y8�.Yѹ�vy�]X�k�2]:��f�����
�#Y�һ�
�L�/�/�|Br�ơ�� �{j$l���KE l75p~�C��F�H���1wi�4�&�:a"�Z�T��)|N�PX�]*X��im0��Ƅ�!�|Q��e8�д"А޽� D��|Ś���'����ъrws��u�׆dd��U�����W��N�؆�_�\htzb�C�N#�{�&��'�94N'#�m�:�vE�[^GAG�5��:Z.���@k���2~���8�L�#���~ �Sq�"�i�q�h{G��qdk��M,�م���.::F2���Sʑ ���77viG{��R�3ꥳ$��B=F;0ml�
#L
�,O!��=Q���y�`��w�4:K�c>�s�W�;w�#�`��q���[悧�I�t��_��O���:	:{���z�N�?D઄��#���Pg���<���:�����yV�ܹ{�}���8�Oq�\����a�(C�̤cni�:�B�Y|Hx
�M��p*	55��Q��5�S���w=u^E��=~�������HO�x�_1Xt�t�l˔�6]���Z�^:�ƃCG���FO�wN']:2�v#�:�Ҝ��ʀlr½�Cv��\>ӹҩҸ���(�Px��1mRN�˗:Ie��\�NjK!���hT�-�r�t�����N�ץy����#G�1�\c�r��6�0ng�N'C��A�Z�J����q蚒Mp*�Vd�F�# ��Ő�(P` C���C��P�.��ŵ�W����jμY������?�����n���oi����Vb��Ņl2��S�t&)����)����;C GNP��2���:U����~����,�3C͊lz��y��a���7�w�a�\Az4 �{h�ﴷ0�\ϠA�ȍ��;a�Ƀg�0�!�4���.r\ùF�t�ʘ��5�s?��K�}[������y�#��eNƫ0��u�/����_c¼lCu��*����oqGg���-fiÃdAS9��^B�<D?m�ܻ � ��3&ݍ�5�n�����ڨ3��S~^�9�����8VoaT9eKcM�=�E[�;�Y1��W7�q�ŝ��)�޺����n,�Qp�S#�����<�CV"4�S�?D���YŁ�����^�s��֝t*��Bcg����e)���f�@/ã[;�Ј�[Y�
��(�ڱe甲g9ƿ���?.e�(� �u��X�}FC�Z�� y@�|��w��V��r���8~���I3��c$�ӭ[�qv�cڗ�5���#����ӕ�,��m�G�=��=�[o��F1��sD'�M�� _��J��3�<\�C�:�3a��t��;����Z��A�8f:vJ�������h[;ڵnj�vt�]4��~�M��-���w�t-�t"�*�2�
:̮l;�!c�ӆn���q��w��.�jqz��#����<g���qiW�r}53]�ܹG�/R���Z��ř�����G���������(@��Sy�Μ�)w=^�ґy�/dm��rzG���7A�ƒ�G�a�)���N���{�r�jq�|���ǒ�L�ų��s/e8B��.׳�GC����Ƶ�����o�㮂�lIR8�$��l�ϝ!t�^�u�~�:��;]�ȲD��m���A����\z (=d�|��
�s﨔�j��&��:�������;yD'��ft�|;3�šδ�T�+�Yᮃ��H�s�����|��Z/K�N9�)���w7���Π����Ik��#\:K�pZ����a��:q��K���6�P��8���
��o���r��s��u��Ag+k�h�ӑ��.���9�I�!�	��(فK��\��a=>�уƁ��^ � ���B\R�VU�T2C� Mdi��̪iz�*�l�J�"K�2�,�����V�ˡL�%ӛN�g��~
����9��E�Yp=�0�_��é ۹�.�������p���X{�][~��u�U��C�,a��dz�,Fҋ�U�z{�j#ø2�����,N�y��k��7�8�V�d~.!�_gC�V������9���9�
�l��hcI�z���5Z���@���^�	pF��[��8v���RӵQ����_f�)��]s�O�]��E�:/n�:B��#u����$#y8*��S�_'HG���^npk�g��L+܉@.��~�o*e�;D�4Y:�~��:��uqd���e���Bv�V�H���;�����5b���Ä��qFݹG��5^N�ۤ�1����)�t�\��q��;�M|C���:��(;��5|��s4E(�c�B��k��r��!F�N��Lϗ�#4'�F(�!0�7��P���ݥ��)�8=�Ò��s)�q(~�֝���:���S�4�l��ݩ�.�u
����3�<mO�2�ˎ����Ѳw��n�S(N�&8�-�&���O�������;ZA>�w��{u�K"��it�^�P���6�A/�� ��
��������N���Tq��p�ѳ�ŗw��;�S�O�����#̝f��q��Q��0e��Ʊ͘=1�'��YIǃ�tR�B%�%t�nk/_��������������^A�	{��ڹ�y��~��d/:]���nK?��y��0�s뭌Z������k�3 ?��{����Ltq�g[)ֳ+A�f'���_9��s
�m��B�:����j��}D�������B���y3����v6X�b�#{�_ٟ���ųe� ߁����1t�"
����!8$3��*�tDj:��	gz��VnP �ȇ�̗�F� ��5�yͷ��ݺÕ6����k�4`������T9m�Fgס��8U����4,ݵ�7p,ߩp:{�?o"�j-��t��U�K�p�Mю�*�_�� :�D�k]�4q��\���k�.]Xl7n\�q~�}�Ïrp�{�Ӯ8�T�V�Sy2�}���8>��"�݇����Ϣ������ĥ8�G�ir*�:��+�{14���)�NG��dzw4F�fo~FE&ƹ�w�liU��ɧ4?-!��v�vʁ�.��Z�ߺd�1?a��K7E���<�o
>�9��*@;�7�az�]���W��7�H����(��zݥύr���<H{�����)�NS�!��D���3t�=G�����`gl#M.ζ��U�:��ZF_f�kk�I�af�����<v�$�U)��C�e�;�v��[�G'�<����p��=�U�Y�~ �����TT>�US�D\����[�3G�4N�S��:��xu��i��R��ͽ�%v�mM;<��y�J���o?����~�Ad�;�:��j��9������͛ql���5w����ȉ	�#W\3�>�w�a�(w�?{��_�`���5<��n�fu���pDG2r�����)����hV�쬆#���o��vʠS0k�/1��]��f�9��w��i�}q��tC�T'���K�8d��)����+��1��緱�ht�k��Qbτ1�L�uM�by�cEt`�?�Љ��T�ɾ'� ���u������H��ҔE�i����6y�uGkd)x#���r,_�Ȳd�e8�!:�}yƍ�G9�A��G�
n�g�����܌����r3:�x��)|�W�Ӵ���*����.���3S<S����R�r�v���C<vG�U�?(��H�I�,H�E^ޅ�z�z��z���:XqPV>�����أ��d�Y��i6b���YҨ�+�r	�^�[�V`��qBt�Pz"\,�������:�(��h�y��S $�AkoօE�]��P��x��{�_%�z��8��aT	Z�x 6:��5E�'H���	�.l̎���T%�ib�4]�6]ʆ8���E�0epklk����4���7�I�9$�(��@��8RI"\=4ϩ�ƵW�t~W��|�FM)%�v�a1N�F�]úO��� �Nن���N���s]�VgY�H@2�����et�9�:X]]�o�Q��r$�e����ߴ��\󖩭��d^�����(
���ar�$īv�����}\�g�a@�~Ϛ<�#O>+�'&꼊r2�I}��,!�,��9t�����t�4�pZyf�=�Fޝm{��t��&󊃅 /�]�ٕ��M\I�N������y�쓎�T�Қ�pQ����#>��]ȑ OAXA�=92�1<�M~t�Y>UتL" �P�䌸!{���[�&mU�Nxa;��>댊3���e���� Ϸ�~�}��١�5D���a��t��_�mw�?��Ѻ�:�RaPk��8�%�\X��.]�sF#��S;=L+?��\�����N�m���۽���\���m�����ޝG�Xt�Žm�L��s����8��rT�*7Z�/gA��wމ���ƭ���[o݈st�w�/S�P��%}�>�ͬ�����e���%��S����E��~�7?h�?n?�ɏ0�ޏ�㎦�L��S����`�s>�4��ЁU7��Јt
uu�]��giMc��/^�`�m~������ȞL�:�����)� ܁6�� h۠|u��W҆�!tҮb]����Z����l׬#�C�H�5�]G�>��85�o\OϺk� =��I����\#�zW��9�v',�P�N��|Ҹ�L���v��۴�#UN�r�g�$y�����\y���i���\�I޵u���h;U����i_��^ oo��^;G��Yo�B�� z��:��.\i�.{8��Ж[�������נչ8b���|���h�M��F������5�\��~��e��!��{��Q;*ÔA%������^�-��֐t��t�o��R��t\Gt��6�����N���A{��?�"������n�3e{9׏�<�Qq=�*tg'����7҇����Ƿ�.B>�u��2��w'�����N�u��Q�f��5����)��p��V.
�Μ�2v@9�t�䢓׶�k�u�]��Lge��#<�5Z��������;�}����ܕҩ�Ҡ#宵u����'������Ip�]�Z���Y�	�GĿ�I�|u�]���.` �/����\<t���v�ͻ;�����{헿�}�կ~����g����`:=݀�%N�S��Q������LW��8֡ȵ��ݼ~��8:�h�+��1�z����_~�~��/گ�U���i:�c�mi�����r��B��m�4���}�%N��VԻ�4�Y�������^�]�ޢ)�\\��B:���';�sy������`�&��B�:F����;8Rq�<�w��W�s�b:���{33�i%R���}��y���2�~6z�"���T��C'˴'����]y����C:YvR��`�d-�+�c�9��dm����;'g�iE�F�B��a����YVX��9�Yr$� Q�!Q|!*��J��J�?��=�e�j��|���jx�� ���b�)!���\>�.�i�f� �t!*3��Ȕ�O&�Q��y���{ �� ��a��Eۋ��	��"Wړ�o�;�m`������$Jr|�Qh0�8�����<8B�}l�m4���;�/���-ou5�s)"�mn�Ǚsq_�ӷw�����p�b c��4;d<!:>Ni�܇���8GY"�qN5�2T����[8
#���(m�r�u�M����ЁĬ�xq�C�4���Q�_.��w����+�ҋ�[a��1�®��Ut��`�v�_�U���ң0�`�\⎒�^itβƵ=�ҙ����2�1�F{�Up���W�4��/ڧ>ĝE�{��;Ey6��<���x�^���ť�iCk�s�%eG�`�����F���|h�s�m�_E��PX�cҎ4�BtDW���me|34����;��s9N�ڮ��|dOUz����QW��n�GNd
�{���s�m��ϖ��1h���/�о��x3r�݅3��I ����mwx�6?Ɵ��k�n������L�s�~D	u��)oeu��{�}����s�(�FwMҩt<S&�B�-���"� �����BGRah�JVg�u'����������W��������L�����)�,�p�@:*H]m	_�=J��2����"��G�H����y���(��K0R��;����Sc�|݆�mms�e��7�������t^G�5h��g�{�}��ۿ���������0�h�ML*o���,��20<^��r�j���#l��98"�Lu�����\�c��#?~Sy)S�稟k4."s���P�R��E�1���lu객�+k��;G�[y��?�)��;J&���8N���Җ�i`#�N��!k��y~�{8Wn���u���{�3ou��J��Ri����)�&�Yf�zuj8}�ݻ��_Hb2`Q�9:p���.���p��v�����yog��`2�
?�c�n����oj�ӽ��4��W?�K9��,������@K8W�^G�q�>�޻ܝ6z�n����_��G��P�z�U?��{:[���t��<�{����ȓ<�I)����Gݝ��`i�P�)3�)�">}6��w#��յ�1;����pF���ߎ�.�θ�TG�����.����yv8�s>��T��w�e��g]�8�ТzRݬ����6��~�  ��IDATY�c��� ��?=�a��r�:rgxuB� �t�Z�x�:rd�b��IӒm�{���֎&iL�uz�����nz�w�n����T]�����Yӎ��D�ϑ,�em1;�u�vw�b�(x�x w�v:��˗�Yí��i�:����mw���<z��N���
�&Q�;:�e϶c��� .@ѿe-88eҊ#�����7�_��7	_|�Md�2��N�̿v=���<�JY2�/�Q;���2]]�eG�6+m��49=M=��.��9�"�������%��|���� _�����i[Y�m�i���&:��@;���~{N�/���~�����>2D[Dg����P��9M��Hm#`��.m���tE�8L�s�'�t���'��\rq3_�e�-w��\to�{�kl��6A��8h�c���,%��|��'啓߂`$˱�NU�m9�M�Q6��9��劜	�`S��v��NO�\��u'k�d���dm����� ��HV�d��P�W�_vvT(S9C��p�Ɣ;�X�1�)�MZ��n��*�z��>�h0"l�ʈpӅw�]��56k���W�{�j�S�6^�)w�I���q�(G�ʃ5������:3��f�u�w������JqB_k�[p�
F��Ta⶧2�F������tFTn���W��.=ެ�q{E�=B-Fgox� �@{\�U�&N���d�[M��s���֖5mb��/�y��/l���v�sA�K =a�g��itfLc�]��G ���X�I�L|�ƈN�iN�tkx���K�c��g޻��	��J��Bu4ϯ��B�g=���\S�>-��҄v�[Fτ�ůu�iԨ�]e�����5�m�(U�8��w�IK�&)V#��^���0FIFr�	�H���/i�iI�h��Wij 8�$�t@��N���6m��*(mG��w���
F��N�8(����Pp���:�h�q`Ҹz�[�!�U9P��'��s?Eu������[7ٙĀ��n޼����5�U�KKkO�W_?jO����20��8%P�����}��R'w~�9����x�(޶���&�5�!�����
�>��7�K�k�T�v�xމ�|4DaԘ�w%��ncX�oLCXZ6����b���AI�gҨ�.�Y���c�A�mm� c��Q��;�g��9���N�����=׾����?�׿k�|�Q�vm�ҙ�.�n �\�^��ʵ&�S����S�W2��ܾs�����Hӱĳ8oҟ�F�(������N��=R΂n������`,�rJ��mG��+�T�4���Y'��#:7?���;k�4(�uA�f�1��О��q��;�`9MN#�雇�ܯ@�txq�Ёɥ�Ѐ�-7�u#ZP���]�˳����JҶf'�ul�uBң#.8�msv�cT�2j��rR��H�����\[F?k��Mֶj|���;��<�n;{;�Q��[2d�o��::i�q�g=l�p ,�e���){z�p\���8j��J�Fk�[~��K�s�«%'�=u/��t�2��g�2}��ֽOGef~����<*?��(q�g�y���*��48���g��5	lV�Y���N:�x��6�ƞ-��юz�K�����:�	!(�K����'N�sz��m4���\��j�)�����gܜ��J�q`ǎ���:_�P-�y�]�*��-B����?�����6Q]��I�ܹ�ܤɣi�͡���g�����\y�^'S�qwEG��/^�����?���V��^Ox���w�����}n�
�_�N/i�v��Uv��NQ�Ŝ9I��cK�A�=��ٲA���U����}������'Y`]�9�t_3�mަ�����T�,������G����sh��i��^H���N�����Hs��o�%�;Y����#��6�4��k�{�d�H�	r�Σ�z�o�Y�N1aV���$d������0���؉]��?��J�\�F{�t���-)qī�7�r��f𪼍[������+�)�ˋ�ƽ�Ų�\��w���;.|����I,?e�֧�#�w��b�C�Ρ�R�\�?��H����l$�su㊻vN�6���o���u��z��t�`���1LKn����dM�������e�8X��DVF�`��(�b��((0|Wx�ANU<�t��8XPL�0*�BT�YiD���FQpN=s�b�?�F�z�X����e���!��,C*��s�ů�h#!{�ϓ��ۓgoPګm� LS�BՅĮ�R8�A�qt�\����q��w8�_�􊐇x�)peC�p�6�?�U�������c�'ړGQy�����:̶�A���,��%�uAp���#~���aó���upn�\�ց�������n9Dr�>�:5aLpdݽ[�y	C�A�l7B��?�G��Q^9Xӡ�?���O�ԇ�i�/1�u �sjA�*�#X̟�,���x�֣�e�]��`��,0d���3k��Q0Mގc�S*h7 v��rz�O[�ls��A�Py��ao�mw
kR�*$G���r�xO�.�Cwn(8=H�@�Q�9���͵:V9H�ߢ©rq�hHqi���7+a�p,%��,=�1��н�>��.B����E��5*E;#��A��D���pf�]�8�]����}�Yj|���ۏ���%|�����wW���Q�Q�e*�up=[F���M��!���������sm�#X���vws�������V�C�4���'�M�bg�施�e�yX�S}ܺ�Q��Bi��n$�u�;(���F����.��J6���������e-�;]�éVʟ��i��A��ڍ��0���t�jL%���z{(�j��u�	Lي�-�-�փ��]�Pz�q�5�M��<�<�:�~:ĥʶ�����NF��ذgRm+�8�n,��ysßM�<��d�g�B�a�����h:Mp�&p��b�Z+&�Ϻe�z1��);*�#;.����~c�������v:�@���2��=Pީ��Mՙ�W2e� �+>Y���
��F�ҞE��O��X#+��ւ:J��ڧ�~��<ȃ��7����Ne{-�e3�=�yU�v��_�ɑz��Cv3�]����ރ�͝TMZ�(���t�P�#X����?t�Jv����WV��:'��w�����{�`��.y0D֪��9V���#���p7]�l;�mP�WJ� �P�v:���|'79q��/���<�õ�u���@��%3 ^��͍�v�SD#�lV��-�;���e\��
9�8v*�6�
���O_����'�U$��ږKpM���6�i~5�⮤:Y�]7-�����QrV��)�c�4�\Yos�k���l�0#뙺:K�ȱ�t�,�Dy
|o���v���v��Ed���g2�ڻ��k��R�PI���/�4s�d����|{����ܿ���3��ݐ�F,O�i*�ѐ5<>��ciE��)��hB�V{���Qd��k�32����*�9��n൷7������}��m����pD����6�΢S|]���?�u����u�կ>�lv���2�!��1��R�����8��J�Uol+�C��Uɐ�\�K��H>�V~1���đغ+z>�Ի��.OJ�w�'�~t����F�s�9��2��\0��,U��\etQ���\�W���.�R���^*�K�7ku��Ϸ�W.d��[�g�������L�v� <�DKP��Wf��c�d�y���h8kPj\�R��$�(s+��4�5Ɯ����J�`�c������[�����WB��[��{	Ab���Օ|I��l��)��C�F����8��0�|{[�%ȃ)�߸�\�����܊�ݑV���VJ6Z�_��u,l����;�.A+��� I�X��x੦g�ϙz��}⠉q�w�j��o�o}u84�M�1b[�a�L�p1]Bz��᩼k�Z�QL���F�:N�p2qU('#=�O��c�~��2�ict�i��hw��������
��wU/;��ډ����:�;p&.��Rh��C�ƔF��{�3NQG_>����w�W��FT*��<h/�]^jN�����9k�U�<B�GhC�:R�+�
K/7�:����(/@a��s�����*O�-OpM���b>�]}̳�W�>�H\� ���N:���*�ՠ�v����E��T���dM���_�׏�Jq��Ag\h��.����A
MJ������C	m/�#~�S�8ZF�(��:�E��;{@����2e$=�N�U&�V���u ��A�XDA�������oV������1_���Js;|w"�����o~�N���1�$j ��H���e `�d��D�h�ު]�wk�/�]'cQlnlęq�hͩZȥ]iH>��Ts1�el�c<�䈊����ڧ����|E]�7�m�P�9w��[o]JG��X�S�\(׹J[��oῙ��N�˚��y�k�֩������
m� M�� T6xO�3)c��Y[�X�3���)�1��ӻ�c�ݡ=_���n�n�E��)���������9;��cG�Q[~��mo�G�)?l��L��cG�����}@��m+;^�^;��i��EN[����/�O�U��T̕Mx�^Y���י�ISQ�v�ȶ��7��/3BL���8Fv����\¦!���qȉ��U�	��6ރ���Kw��n��7� ��qv�t�
۷Fx��5ň4�C	F.�����*x���y��~�j�yn�=�$_כ��v�D	��PX���8Yi��t`uih�������^�u�M��5N�K�;Ȩ�i�E���,pe�ƻ���Dl�g�s�ӫ�7�2�c]�Gpg_۽?�T>|�xN��o�d�Vsd��A�� �Bs�
�:�����;�����Yln\�����v�(F1�*}�ٖۭ{|���OiO���[�L�we�a�7�!_ԗ���o�N7ux���f;!�Sěp�L������I���3�ա�1�.��K֠Aw��gCY#��kk�� ���e�>�&&��7Zq͖#i�k�*�n�ﵭp�����ES^:9v8���_~�M���&���9�!K �f�d;-�q����u�R�
?���ʪg@n���IxK�����3���^"�?}�<nƣv�=�Sd���݃GO���olb*�/���ء��v؁��W��'���_������`�� "�Y��Σ�Lh>�Zjtp^S�pr�qu����%���C�k���e�iW�|W���g���=b���ґ�d&�F>����O2�;�Hg�A��+޴*C��qv�u�w�'y�:�4Bb3�޸�w^U���-|A~��e��ߴ����,���H��N��������
}���̍����$1"p��W*��L�dU�1�a+�eoOz׹k�� YVd�h����]F�Sj��Fd	����&����CM�1H8��#?ன
�N�4�c�ڃ���@D&����/��:
"Q�Ef����~�B��'�~�|�ka���x���^���f���h�E���H�8�D�k5��\!�G��� 8�0a�j|֙)�����z������o/Mg]%��v�KY_qL'��A7r����Zo�%�4��!3b��Q�S׵=�9UgHE�s�5�H#�SCubā�06ߌ�Z�(E	Y���¤P�S�����v�[��z(	�:�@�B��$��%AȨ�{&j{��Y�AQa����ѻ�� q��uΆ�}ViTZ�|�ѧ�nE��con�F��LFS��#h� ���ĩu&��d�� �1m�F�q�����8|�c6���|*��T�k��x���pB����1\;�i��������f*�%
ҷ�K��8�L�c;]��n02p�K'Ɍ7�� �?�N�M/��x��F�=���=q��i�����;pj8*��y�I����K��6���:��{)+�^nǔ;3���]��&gf�!�}���oo����F�J��ɢh���htժ]9=����T���z�zcuE���.c<E��i�GI*K\@���tD���U���=�GQ��2%�v��~�WG�֘�R�c@<{�a�ƅ�Cmsw ���XmO�1�]��f1�;0<��i.�8r�[8#���G����C��1���ܱ�v�6w�������9vG��!���q�T��X��ሠG ,�n:q��?o�ű��_~�C�M{�����3G5&i�!x���9�nj���V&�ɗ��9�8k����$!�߷�ǡ�����JF#���>��S�� ��
��!�k�5G_��t4@Ñw�V&�j=y�_��
�Q�:m;�8�N+�`\�k���f�9~���4���&���x��FeP��~�#�w�縻�=�:~E�NiŠ�m^��&_`$�I�S��2�Q���r�PgO�`d����?�@�/��i��is����d��%h|�f�=�m�{`:0��9�v��88%+֨�;�yΟGA V��699�nim}��eҿ$�%����,���_dm�7���A��?kK���M2�^�u�:j�V��i����GsE�y��ߕqW���=u[�?� �2\;�G�o*�ݳr��S��l����#��CGip26��3p��Q�G��q{��%�6h�����B��@W���!A����Sv�tx���~X�,��1��Zd��ȥr��TF:�O�83P���-��+w��i�Ι�/�	�=�Mtы���������8Z�����Ό�T�i'!ˇT:�};"����6wu�2�<x�����<;�����o�z�׷:?JJO*�&wv<jţX<��s��/�w��`c�mgL�;����n4Ͼ��H��;����8�:��a�����B[X�#G���pD���{�N��B�M�����(��@^P�k�Ch;�t4�_�,MZg��A�9�����:�k3���Ѷ�5��,�.�v�yv彻/ۃ�����K��n��t*��/�_�3"�\��<��A&�`I�;�a�/��l��~�>��;�z�6��LF@�4 pB�����^�[�jl\{�N,�Y8	��c�j�Gm�9]�OFqz��7\!.�������b_�OqL�ߎ��q�X�S=���ҏSٗ�[yֿ��t���i(	<H��Ծ҆��A|�e@;��T���v��e�I?��y]����-r�l���)g��΢�L���#?u��^XlW�A�o��^��j?����?~�i�5J�9�wc� �8Y@��)��tAO��[�1�p_����#{x��&C��Q��)�����\(,i�<_Ear ��\�e޹��Р���!N�U����5�-D������%x}��^%��*ã�$�	�t��HC�n��]���v�4,�϶������/�~��G���K0��yo�_��������@��&
&�*$[���
�j�VChd�@~w�N.�I��G��B�q�-�~7���kS�W�p��gq�2,[Bs��Nf��Ѥ������Uh����e���a�)�lG�}�^��Hk��5@��g�8=<רi(�6{Z�~v*�`{����E|Ȝ���t
PFz���c`��.i|�Fh8%�42d9a֝����TpR����0�SX���M���iI|r�hV�d#��|W�jP �#Q����Gyc]�V�'�)�t��mT*�
g�5������|B���㸙�����n'ktR��ʞ{����Kr-
�k^qڨ�EDd�-x�����%�5`��ҫº[#UEHQV]��iuʢL�"�^��?l�����w׀�j�#��A���!qx�.g+���j�������o����3]�mt��߷���Y/��(7�1_�
�Q�R��[EG�=x�P���ɶx~��q7�������:�R�3��7:k(,��~�����:��"_�!M=<r:"F�=�T�kw8sc��v/�^>;�F8=?���Ͷ�����(�fGL�=��; O�l�� V����H?���n����n�{�m�/abp>%��}�P�@�M��|��_��{���/ܲ�-������Z7�M�>��?0��M�R�1���q��l@����v+�Wod����t _<,�8;B/E����Os���)���fN#��j��d�螛�o���m����i����7v�D��^��|�L����(:]�-�!�6�Q	�����x9�Eg��KϷ�-��Õ����Rg�y���V���Z[IG��ϵ���j��裬C�whO�n�������m?#�F�iU�Z�9B��}��N�D�p~��s�����kW����1�-����M�_��y���;R��cD���@�9p����t��P������)�K��R ��F�˖��ŐW'b�����Z���Y�ǟ�� 7O9�#Є���]�vW&ˋ�{�p Mg�[�O�I��D�N1U��o��MG���ʫW�4��|u4�9e��hۡ�mni���-��0�ܔ�Nj^�q�gm����+�.���=J�3�槧��v�R�U'���q���W:cxp�2�Wg�=�I�Ɏ(�	��gǉUG7���<:>5��6L���k�tP�)��@�G��y� ࡥԩ6�pʠzTG��{�)�g��KN-�C�M5;?Ğ�8g(�<Dxjb��h����_s��<3����LK�v|�-m�g�8�8kn��&'�p{H�����܇q^�G<{��t�j8��[�Yp�n��>j�O��n�ho_���Q4Zۂ�<pۃ�����8�� �F{��:4�n��(����Q�4�������1�;77L���&N�붹��15�m�vNE����8::K��4�]5��yd���NmmG|�7�8ǎ;m"٨��h�j��6�)�e��FYfG��ș����Q_h[ʬ:G���]�.�<�B��K��\���'�K�����Ĵ,�klK�HP���D�@�B��ݼ'���>�h+�;x��3eR9��I�y�s��}t�4�����?|�������w��\mӣ�������'�.N�Z[ߑ�a4�Ue.�a�e�����R��X�(�ݐi��E�E�Ҫ�0F���'��;aEU�u�i��9
4��"�Sq��v�|
x�C�d�F�m�x� WP ��]w�1O3��ߥ��)cz�͢$�mI����U�\��8h�����[7ڿ������?n�{���"p����n�կ�l���������a��88��\9}o�k��{�_���S���C(c�<=.�I<�� O�����5MK��C���i������<�vY��u�d�SK4�L�=�k��t�,ǭl-Ӽj*�v@ث\��)Eg������|,<Į<2��X�)��O�q�~fڝx<�C~��ޫ�_�}6������)<��
�j�"���鑤'i�� ��+��3oFi��r��p����P٢�Tlfc�Nߡ���!�����x����Lቼ���F�cu��;��͒�)lS�y�\�%OG-�)#:&�)0��;\��%/��S���C��O����"���N"ѥI�8S�F\��rȋ5B��LEn�4B�[+=q�����(ġ����x�އ~�L�1�?�}�!"D�d�r�C�7���H�+�>�׌+8��]m7n\k������������McȮ����~��_~�~A�曇�"2{��)mt�̣�:X�/�[f�L�Y��1�F˹��rd{�������d�=���q���U�8���w
.`���_2�hT�f'FɊ���)7g�8w1���Dd�g}�d-c��x��s�w�'�U�Y� :��t+�S���<�������68|���10��t�4+�t�3���4n%�tG4"/���A �0���<!�h){\��C��1q����P�L�3�0�GF�k������c�ea�DWW��B�kѓ��Ff6,�����Èv]�X{>�0r�A:��A6+w��u�bY�2�d��3N'��?G��5��pJNЯ����&}��{5�J/b\��N�n��S�q�3*�0
vqDm�[����'�~����v�\~u�i������?~Ѿ�ηv�	�ՈM�ߡ30�#�,	���ܕK���o��b�n�`�d�����u=Y�nḹcbGp�.mNTg��&;�hku�܄<s�6�(�2!�|K��X�7�˓�[^�w��s�ǟ��=)�giP�Q����;��4x�F��� u�n���iy
���=Ng?�;N�D�ǀ��Q�se�ċ *_2"E�u���d������2���C���ϭ��r��D����{ؽ�W � �sF�=�Vt�4+O��.񥼓��s�85U[l�&t��Qm�~���Je�xToH�Дv�VZ5��ܭ�5�|vq壝��s�Q:̚v�G�NJ�4��Ax�a�(��5v2�C�9b��A�۔���Tܽ�-����s��$+��yĀΛC��Á�d�;+�Y��Ҿ��h�66t��<�s�s7����SV�a��7o��
<��P�ڽ�nfgk�x�A�=�M:������٤>v�Q�r$� ����_G���F�fue"��!hB�!����LU�ZR��;eZ�
i[9��N �X�U_���!�� D�{/��8/�6;�T�U�Y�v��,g�wډS��}Y ��>�v�g=4�7����zC���o����ʺ�x+�Dϡ�h�p��3 �)��>���V��󞥌�i�UG:k��: ��8���J�8Y�o]���'���>��V������5�����?u���<yٞ;dA�Ֆ��IdL��d`�h�iP��4v*�, ��4Lz��Cj*C��:2�U�X�!���*ÿ���a���e�I۳�W�2x8I#�]Ceޕ���$~��� ����!�y4.5$h�bAg�F��Wۏ?�^���wڅ�cmT:G[��.V�.8O����j��8���l�;�=����ƭ�g�
5���8�~j��i����f��'�F�gZ��=�s6q�+��4�#���Θ8���J�D�;����L�Ŀ=:?�4�kә�maZ��$?d�]��^�4Ng�PA�՟�,Z���AF���:1�aB���J�g':d=��<�7���9�q�,	�X�Ο��p[��L ��`�cqM:����kqf�x�O��2�>jzqS�)�f���J;릀�v.c��YE97�s6���`���)��2j*b񁸪���{S��T�����he(F|8���|0���os�)� ���n&!�nn�զR��0p�oR`�����Y���9A^���/�2�:(��nW�:,*��q�������� ���s�v& ��Sׄ.^��Ƅ��:����kW�[���29)#���0��ZGS|�ܳ���+	�5���8�����VЕ�B��ٞ�r��?tj���l�L	��d�r��1�R�)��]��ʒ����44�?7Dp�r��qrQ�Ӓެ�Hm����H���k����2�ѫ��47���i��`��Ħu��߷�u�ݥ.���U{��iv�sڞ�,s�;���w�[��9�$[i6�]��v6�pȷ����y>  |S&�k�ӗ�QGB�6�T*gXf����P~��-�^~Ua����Q`�,�׈0m�l X7�p��&�]�����<�Gz��#f�ҹɃ���v���U�Q��o�@����Fk���:�îy���1r߬���_6װ<�>�9v���[�&��6���(��<�}��v�ڕ�o9<F� ���L_tSG�A�C���q��w�v�����}�����i{��C��e9�f;;re���n���b�J���`���,�:���]-^��w��)]p=$�{�f]�O��q���\�EjkiP�i����𺆦���%�pN�Ӟ�mڜ`�_�z^����+~�������S���B��,'૛rY3��(�����r�c|��Q�x�$M,�/�)ߑ�M�Wg�ye�e(�Jw�4���KG9��/���+#Ч#�q����t�� R?�p���e��S�a����Cu�G&�a�v�(�9N];�x�
_=sS�%�@�����d��4�o�[G��ZS�蝲ȳ�=z����t^��3�ۡ�8�M�!k+��ǰò^�����UR�{*u�3e]9\/�-�>T*�{9���E��\�Fr�0ʯ������g� �%���mG�A;�]������e:����ƶR���G{iw)?��r�z��35�s�((푶/���wj,�C['q���_�Y?��2��o��Q��NW�_:���v��յ���y�.��0�7�a�j_����)m�����'��s�7��A�LS'�8"%lڝ$XN�^-;�:)�o������-�Ż��!�u�A:3U�|�\��l�gq�G���;$����j�?�4�l�,N�&7���d�	*��&�&^�i�W�s^0��j����&�6�[iȴ�_�k�`x���x�1"�+��i�i����Q���wu'=qu%�1��T긌J��|��u���nj��^��UN�F�QAnCV�2�J�.Z��yÈ�1����K&�)�tXW�>�n�2�}����o�h%H~�^1x��+�uN�5m����	�}��!g5U#�����l��¤!d�2���J9*E�ʞe��dn3�97e� Gؓ�d#fZ��1��0��J���1ҩ#p(��T�U��6��+��KϮٳ�
P��#h\S�Ni>k��G�~����H/�F3��2Lgy����rR����ď�U�	��8�[�:g|qX�o�+�ROBS��x+dTE;�Cc���4���s$t~�M�-��O�_l����+�{�����6�p��;�-\��	<OΜo�S	���	�8a���4|v�#FY�)��N��u5��u(�q�¬��h�೻������BС�P����|&�h%	i7���^
���j��w��D���CNPa���w龣A�*Ȅ:�督_#�:�F���G�-��>��B�׵�c0Y>�S�_� �S嬷k'�o��]P���֔m�@�p@�{�U�v�P�N�ECCY�k\�`�׏�㼹��� v�u�Fx7\k�6�v�����ݧ��ۏۃG�K�8�:W*ԅ>:��9t��v%҃�i`�#���:Q�_8�ϭ�5�\�0�r�=��G��y9�4�S��v�,���D�0J����'�EY�T7�p-���(��e��ٻ�A~N?��:�GG�9�`3&����� �!�Evă�������gVy>�|g Gk7xs�Yw�u����>���f1��mE�?�θ;ii\�a�A��{C�8�Q� �K�;���aP�/뷊�⎗Oh�g���{���#ȿ�m���v�����~�>��ߵ��?����v��[��L��-��Q&�T@��-��;����|;B��L�?׉�gK�9�݊��zm��m�>��IBv���v,�5��mGH�+Ym�EhL�_���s���`<�j^��
������0Oy�/���Ԁ��M�3�$�t��iΣv�M��}�E�5����Vh���ݶ�C�����S:�3K���5*P��R�@��_��60�f���2�����KY#N5�_��������W8z�"�3�C����G; °k:��zEO�Tsw;�ey�9���<^S�D!3�߶��w� ��1�l�.h��"?�!|9�-���7i�1H��<+��G�9B�Xd��8h1�!=��Y ����mn�h�d�܋���k;5�'�ϩry��|�A}C�I?9��w�}����S� h�ڭ? >�Y��.ru��v{CY�kn�a�9JY���3����ygt_ݣ�]	�h[;9��uOy��0���Tm7�����e�#��8[��U��ؖڦ8:j��KٜeG���6RxI��y/S�v�Qt�bG	�x�}+]}�4�'�vi�*9�uv�e�<חe�Y�'A�k�ص�3ρ)eHtZ|��a����#��e�V ��V��q�x�e��#�r�ܗY7�T��G��}檌�"ff��D���x�8:D��FW�v��2V$�)��1c�W��g�:*n9 �'�ͻB��.�"��2�E�����p��M���Ǣ����Z���#��iҫv�/;��%-�q�M�= 5����Dւ��+��0Yn��8y���Џ����M�#�R��@�n��D%�p'`&e�
���p�1� �G$S�0!��e�?a)��]� qH��1��4��Q���Gu�T:Fq@�������FR0i,�9��$O��6��c��F�d}t I�1��[�� 3������J�Z3$>qR�{p&�y>���4�y�������61�a��y�92lʌt��v ���}�*&�84<�������l�
�#�-��Vӓ�sm�ܹ6�x��.\j3�}�M��3�_� �ئ.��ūmz�Z����66{��L_l#S�̹k8_7���y�U�]��s�:d7��K7���on�~�na�J����&q��0F{�lp�x��([]�LG�݅͞qx���:_R�M�G�� ^��z�6���8,\}�Ҳ3ss5m�NGH�m��L�1�9C\s�G�m�b�\���
�4G�������,%Y砡���訽ts������1JQNﴧ<t�?d��8W����P��U��q,ʂV���v�������&��{��0��덚����2W�"4��&{`�u9�"J��-[ǔ�H�����3�5�a1�>����wGS1�0t�DC�t��7<e�g���De������̍�n���b��uz%z��r��Ԝ!����[w�ά�ǧS�����@^<+�kC�B���s��#�Q����n<���:P����3���Ja����$t�����%/@S�cd͐��ȝ]hgsZ��k{���ā�'���׶`$ח.^�����ڏ��ۏ��?�������I���������o���o���)���"o�>|��ݿ�(Ӥ쌰D�Ri��\��ȕ�8�Aa��]���H��,Jw��Ʋt�@磓₶/v���}�$�g�{��&J@W�֪}s��������UgC�	���ʕ�yȏ�"�,�z? �8�N�����t�\��@���`�'�@��#�[gL�؟������Pp��,�kk�ci���5���#��i���N��ء]��L���"�[7g�� o[��K�4B>�vL�Ɉ3f|���r���p$�f)���]$��ua煭g;�ME�ǥ)#���(��N f�^ҩC"����/X]�X䣉���qg�7�EysH�op!�0��<�67%Κ-;Iƨ7�~\+(OIC��YqV(۩�vf�*�t���۶�\"��#zV߸���u�3�9W:���������z�:�ݬ���P�v�=��VvӲ��919M����4�L�-�b,�Ɍ%Bě�^�٪uזϨ��~�9a@�LV�0e�i�*?i[ʊ�;�I�#�s׶ɨeF�j��4�A�c�
W:�I+l�Y;��)؄�6�^�Z#�����V�r��M�ѽ��%|�3�tl�6�ā0BY�k���i��|ɿ��w�I}����<��b�[����E�;D��Sc���R�,1��$�ݼDց��*��4]���,�����)y��'Pxʊc�=SJ(ǆ�,�b��������^����dA;p7�[�U�@͏F&?�ɪ(�,*#c��4V*#��� E���h����EBU��7�l�Q�ip���1>}F�'nFU�S�.��K�ғ��
�Q���9 ��)���N���lӖ#n��@����R�u�i�|��@�����M�;�s�� nL[g(Ya6M��=���mo���6���x�-s�OG�r�k��F��(<2�el�T�5�`^�5���G����XE$\nP��� pQ7Ɗf}�8u���"mFulW�'*Ǭ��x�c��:%���j��"߃(5���: ��5�����T��kSs�8B:V���3��ad�|�ZĶ>�Fgx��5y�*�����ؼIs�`p��8�l�z�J�ɚ��f�o��ś���[���wp��m�.��.]����8Yo�x�p�t�fp���qg���TD}�l�r����hP� 4�2� N4��%(��Rp	��a�8�<���j��!��xa��w�n��BY�.��w����:B~���J�8c:��:0:Ђ��&��ك�P���dy��T���5"����r�� @�7Z�|����R*����o��%e��`z�ɏ<�b>�^4�bԌh�+�Ӏ➘r�
|#
��h��)�ʏ����F���+�B��A��R�P�F�#���mgZ������S�-���g��UO����G��@��C���hk��F)%m�G��H�b\ 3���(+�G�l��R	N{��A��iY٭�@��[��ֲT���M{���.5�\����!gm���u�\��:�pv�_uB��`�6�z�Aj���>�c�oa,y ���	����l����퓟������}��?n����v�[��ծ��V;�r���<:�N){��a��/ۧ��?}��c�U�/58tx��_�7��	v4�{�)���6�����Z!��^�q��5�{c�B�ڜ����u�5������Lg%��j%)���`�^5?�p��y���5;7��upy1��w�m�w��vwh3G��߶��qĳSL�>ġ���_�/�����@�y�A��e�G���#�l��D@��u��[�$`ր�uVt�t����yF�p�»�?"��a�joCUg��B��d��*/w��,����6#�<V�	��r�_��m��	�[Z�ybv�!u-Րp9Ep�r����͠lp��]E�ѭ�
ʋ�s:]FҨ���ߔ'9�N����rj��9�� a�}�Վ!�ӺN�u�YW����m/e�uTVQ����]L���M�o�i{���Et�#o���i�֛6K��U߁i����� w|�́?;���c,K�O$m�3�G��9�N�r;S��]����4������Y*�/�9��K@�$KFh7���"ʂ8>$�G�uꘝZG�l0/��i�۹oA��1;n�E<� ��Z�*�}/��N�,���%BY�o�ı��#R)�Rg+�e��)�۞AV��NW�۫�N/�r�(�N�
ZF�eu���������|�wQ����i�p�0�GO���7���9,r�y��	Qd(�q�5�(�#��6B�$)��m�M�#�����.���� ���"���ie-O��9@?J`^��u�JG�!?��3�1Ӄ\0,��L9¥�1
s�\
�u��;�d�q&�cjr#r>k4\�m��^A߹�$��߬��Ɋ�&+c�T�5J$��[p*�����r�w�w����R'sg͓�-��.`Xe�pVg�/���l��0Y/b~�����Ws�j��q<SG�I�����ڷ�a@����"k�uu�`������i0����룂�a�Q�@O�q^pM��vlk-�<vq��R7~P?{j�,w�ѩ�hKӜ0�q��ʉ���4��u��X[�S�qlSaT�R�8ёtdM�0����F22%�&� י�j��H�Q�j2��P�Iӈ����*lYcBn
�M�a
d�SƝ�����wZ�B{�	�{�3C8p��q�.�'�!�h�K#�ݥ�1�@= ���0�Kf���F���4�
N�%�k�j��T��� s����ԋ:p�qנ�nm�L?CYU��7�o�T�	��]e&O;�M,��ޅ�LN�F��95�)��a^.ƞ�k�s���1z�ƕvn^r=�땞��fN�=����E��k'�!�� h�

��;/�慲�{�$��O�l�X_����\��8�x�m�dO0y�SX4�#�z��ϝ
�I񁛹(ls6M)8 �j�����g���-:C��䩜�4���J}8m-�L/|Ҁ����o�Pv��Hr�:V��.:���r:#M֬�J��r�;;�YcYv<y��m��M�8�N���̫�3�35������(�(�#�|�]�=?�W?jZUܙ$�#gq�s��
X�).  �#���`���q*C�� x��w�'?��}�8V�����sȄ�637������L�(��5;�Kv����_�/���ݽ�0���X~�Q,�����u��$�f��Ձ'��+���N�.L=���W�Z�<Wc���/�tnB)6|)�gޚq.������ղҊy���;Rj���"����5���H��Y#͔A�׌"�O�j�:^�Ȼl����eР�;!��ܪ�P��C޵�BS�Y]�#�>�Ъ��/Ӡ��P�����ҟ�2T�$����.�)���I\�γ�!3-�wf-qy6������Ͳa�]�I���L��8-�w�ˎ1+� �������^Bc'�=�V��]x#jk3;>\��� ���XI�ٔW�}:^�R,��:<I��:��W��t��O} �퐵cV�.8#M"�6�#΍z�Ed�(,W�-�ù��w	Ԧ =�R~����+� |:gC��mk�`��Q�lP���������Җ�2}^����W/�u�X3��_pJ}��⌉���o6O: .z�4�xi����z����i9����J:[�鷂�p;�T<�7����eN��r�5^����Bۄ�yUGz�c|m��Ɋ�!N�w���a���ە����:'k�rMV9Yx�F�(s�W2'����*z#�QT*�1�={�(��I)�K��~�i�D)�қG:N/���#7�YT�g���x-o��m���Q�[���zD����;	:e/HYE�4$NV�CpV����	`0��4�5��;7�ϟks�s��1�#O�x��s?>~�sE앳"�4*`��� ���(�w�s���w�{����a�ġ� c�9�Q�S�u���i��h�vL0]	�rh�(�>�~����BG����2�$�8f�U��d(�%H1{�dZ��F�#��e�嘇�����A�q�!f�����̲eh뿻��,�_F��⮧�Tګa�� �Ih&8�e� i\�"DO�f��Y��vaP�P��գ��^(	��Rt��J�N h�%MO�6k���������=�*R�eۓ�.4V�eC��m����|���kcS�9+C�j�`�����\��t*�
�a���t�~{�Ӝt�p=����2��P�I�����1�3B��^�~��'d���+��{�T
Tڬ�q�J���%���Z�L�F	x��%B7��̽�g��Jn����gk8Yoݼ���Ѻq�R�������������=x�Q{�f�쀳�g���pR�u:�j�ʃ���G�5镉*�вpB��W�}G��#I�YY�*�ޛw_z^��pk*l*r�KI���sk�����8�[D���4=��uB���_��1&�>�m�?D�U�l�������=�*e�?4 }��^�(g�%�F��s9B)����#�,�-HP�7i�L%_��E�Җ[X�Go:e9��7\���%ͩ��ku�Q~�Nz�6�� �(��\	#�mB@�?����u�*4��U(;�O��p@�R���y��-h���>�������<2jV�t�e��#��y�ѣG��o�����ѓ�Ẏ�c��R9x� xOu���ӹ�SHz��)*+���+�9%�kZ��ɯ�m��;�({�މ;U�V�ۆК"��,��BO�g����O���{��pL]k:* wY�k1�c�R/�ɗ�N��q��"�6���}(SYh@B��}ۓ���}�	��>(
���f�A����4R��t���ʑ�'�j�A �C(H&W�=_�Kˈ���	�ꔩ�;ya�޵����XF�%�V~���-�1%�WB.	:T
e t#?_v"D��`y�]F����%��}@uu���R���Ѝ�����V�6V��Q�Z{��z�@��^�*��F��n��b��[�#O�dE�w�����qm�4���zXߌv�~�{���w��ۮvlG�i-�$Oa����Ē�j� �� �-��4I��T�Z�MI�L-GC�o?��L�-TXH�H���*k[:��L'Aj��X��m@��c��%�魣�lߢW;���R��L���g���m�w��ؤ:��B9������fa#��ph��o�;p�������w3�ql��s3�ʥ�l|qaa��,G�>]j/���F�`V�����i�#�u<2G]�5�P,�A����9t�Y�Z��Ґt~�Ʈ�Ɉ�(D$CZX.e��.¬�#"N����_pmCo9�K��/��,�Z�JPD�q�`��=�q*�G��4�O@�R���&fF�9{�J3���֖�7�`=y���j4΁��2r9M��x.Rp��jK�Ρ2�+����	�!l������*���嗣q�"�Q�`�&N���]#���K��c�oӈ/Gk�B%q�bOO[�>L�{
�]ě�o|�mm����r��\*m�hQ�Ndl�C�YWf�1��Q�]��^���.�5�2(�i�ǈ'��)�tŤ2�4V��6N��N�G�'tCYE�Tec ��IkO��f`a�N@��_(��]UrU�����%dN�>xЉә5MM1PP��.�O�����\`q��؄S�\���A-ӳviNwRr��T�/���􃚦�P���oP��PT�Z@�o<�S�@E�w�����x�5,Q����S�kpX���t�і�"�[��j�w>�\����_�{�Cy\:�@Uf��;8p4��t7ΫW.��޺ڮ]����I}��U��ot��?�.a�4Oۢ��0	�e�/@� �!����ށ>�C��d�|�@�E`=�7�䝪S��A�g���"�X*o	 �h^����~,mC0�8|�Yp9V�M��S�)�^��'WJ#�u���]>C��>���xȸ�2-�ąu�9�bd3�0`�K�� ;z݃3=֔?����v�3����M3���t�����A�N�i)ڪ)T���Ѭ�A]rN��z�_)f�DŠ&�t&v�Q؏�#��7pXe��z�LCm?7夗�#a$T�euʵ��(��K�Ϸw߻��}�]�K�!p(h�<8��(S�n�����_�_�����W���'/���Vx�vń��x�ړ*vV�'����U'�#g�z� 8 Y�qʐ+^(C���B�=��B���߉O�$��J�p�]���Ⱎs���[~�1����X�M��OO�:R������K0�!�Z#�p�FI�+��|�7��7⵫\�邼+�����x�Dީ��-Oޥ�^OX6_�%�M��x��2)-�t�{��e����?�����Q�7^ֺ�-��I�|�y�n�h��^�3��,i���ᨩgU*?s�x�L�O:O��a��1UKuz[#z����; ��d%����b^=�h����I�_�tik���t�R��O�`�����¢��韻��(e��Yq7�C+/m#Q ���u�M�,�[�u�P�������Uy7d�(2�Amۧ��0 |B舌��w�p��i��'ӑ,R��]�Pu�u/�L<Xk��JGU9�I�X�X	���4%��Ɨ�+�r��ڬ����s��E�S��2�8r�w��oӞu��N�
�y���|�5u �8��e����uq�]���������O�����|�=z���X~��Z�'��T$w+v��q#��OO��Rk`����e�6-��(���U
�Y�AE6 r����)��s�B���9�;{��p�������Ձ�a� �h�I2c��vN�-N9��ޢ؎P$�0bN|�^{(�����F�7���o��W�TG��qz���L�ə�,�}�z��|�Җ_��WK�mӃ9-G�B�D��0�!�.�*" �j�3���H�@#n��=���z���2Ycs���YC��IһH�d�����߭Q{F˔0���v����g[)@B���Wz9���K�%J��͑%���^a��qT`��JB��1A9��Z����n�'�e0�|T��G���/E�	�a����3Y"D�'�q;RJK$��7����$9,��v~�rF9��h�
��|�����x�TNb����-e��*X<�8ܲ5�d���(ut��6�|�&q'2��%t���t�#2u��*��>4�q\�9r+tYa��Cyq�d�̩G0�WX��[���l4`;��u��12���"޲IzH��`z!���עk�G�����%�0���0�!�\�_h��2��T�Q��=�!0�ٛ��+�mqA�s���҆�)���� D�M�� ��i�+:Y7���W/��i���8v۫W��ɓ�����m}]���D�7�8�6��۰�M�a��u�n���?�ո/C�銶~�YwݠSO�g�V��9wm�BuC9�^<�.�G�T�ʊ'� L�*�V�7q,�!�#���_�:�&_�W�t���*�;q0�󍴤w���%�N�,��kh�X5�T��"$�8Kx������ΐ����Gk)l�4.���ʋ�*O�V' ��(Yd�2�gg��`T�l�)Z���Q�!��5�tZȽ~�T1��'m�_�����Y�%���SiY$ B߉A;:*l��}D69��&+~��qڜ@�����\�ts�A��|p�z�sz�Ƈ�jU	�:hk��ٓ����ڗ_�m�?ooޠ��g���/a��c#�4�җ#����GܑU���ŭ�' ���vR.R25T��G�Ʃ�G�m�,�,KZ��8�&a�@	���� NB��UI��W��6����ܤ;�	n�,o��A�و	���J���>J^#ǎ�����^�@y:�J��[�9�C��C��Jw���8,�%��Q��
?�	���;����˼�x"ҞwjCZ��Zg����P��1�q<$+�T��i��r��J\?j1�&I���T�*�G��bѨ�v�lǦ�����,#���Bo�q�cQ mP��.`���H����$J�>��.���&#ś���N�]����H}��:����LW�j�x�4kx{~���r���qv� ?�����dpʉl�M�c�v��L?%#��U��V���m��go���k*fk��G���
��,6e)��i�C��/���Y$��C�C�z��G��{�M?ĵ6��vT0���%-�� �HGY�����6�eh�ٱg���ƳV�X��2��f��TD�$����G���A�M2S�V](K�Yv-����6;}u̴=���K-ĳ��s�o����V-Lc�K�_=�hY�hw���d���lW�ϵ��ܬ�M�l�����d���r��K+9�-~�,s�c"뚬�.�| �hL�RH�᭕i��u=q�H��*�R(\�bЙ�WFbh��H�w��R��*�h|�]���RJ@�M>`q���=��-òd,Uc�<�Rb9亅��:��s�m��B[X<�ff'��������ޖp�޼�h[0�þي#<�8�Sg@�*�S�A�g��K ���Qp���_ن��֥�1dX��@fc��
��ե�<�������<�0����#&��bM�6_F߫��Q�/��N�s��+�H*���ey�;�E�Ʊ���G������C�]?HE����f���a�Ѕ��mm�|�*��4�2��j�B�0^�.���)��k�,��&��w�g�*��xG2UJړ�0�H�R8N�1�)��<�_�u��%ؠ4�8�Ўla3b�ҁ?�(�߉��,w�+\�����ԣ�����Fީ�}ߏj��Ճ�s�<�K^����E�q*�o�M=d$3<�� &ꬔZ!�������o����{(�7#�A���E#"�}�.]��n^����t�Qp��;9��#�O_��-Q���d��`��ˉ�-�6ڢ����.���|��O_�%�W�xw�s��X���_ '|}��n���i$~�91��U��a�>m
IߩsWƷbR�z�]I�G.
j�N.~w�}��d�E�^�pT/#7�i�	��O�<ŝ<�=����t����S���?�t۲:��2jW�A�pW�H#u��,�h�[C8R{����"x���v������Ӝ��G��:Y��K�D���˼���2<��zNdO�w��{��N]{%���?��^&鯼?�P�LH9��L�1�PW_�i��� ���>/�h��w���Y�'߫��c}"�m|��!F���@l��'�j���M���'�������m���ꥡ��)�I_���9�	_"��Ӵ�޸���V=v&3�B�\ң�b�i��	����J����BQǌx�tz��_:�ŝDX�P�K�}m-���?�KSG��J�L�C#/T ��#]�S��幜�,qLG�UF����?�TW� ��:��B�u�\��7�K-�w]�\�����K��t��zu�}ą�X�=�+ǁzr��e]��D���L�^��V����ԃ�Ʒ؞ST� /�ov�Nm��|:g�q��9mJZ+L�}�)MB6�Ԗ8Ih�h"�I�3��6_��h��g�fdr`5y���ԟW�i]�DWh�����)�d���ۦ�G�&��v���vnn�MO���:'k'k�=x�"�70�0�4�ͥw�D��o����(e�>�'���L+�JwLP�+R�h�ʿ��r$�H����q$P�CD"��!B�SDQƧ�a
A�EH�[h{�G\�ӭ�əB�ar�j����v���v��嶸���������ߖ������ب���9}/�� &��W:\މ N;c�g��L�G?�r ��t�jO��x�֩���Wu7M�PF)	��D"f�g"&��sa��K�Й&^L�3a�����wa(b�9w��.�doc1���Yu�}�����sZ�6�6��ev呱ij
k	���i=�N�,#�#EC�|��/i04D�]Ѐ�v�_�u�1rI���;aߗK}�qz	~�qQ����S@���o�9��p�����y���w�6N�A�	?�+�UPnU|B?�_�+{-���6�?P�H6'wۨ�
���&0�{�_��V��t�v���t���yW�~�QU���~�N���~��^9X ��+o��=o�׻W������l V�'m�|9��Ю_�֮]u�q�{@�.�����ы���R���r�cX��O��ʶ�g�-�M�"nDj[U�����ÙD�:[�our�.��W_�Y��V�ϻ����u!���.�?m�>�����;���w�����*��W啇��-#y�ϥ���o}�/��Iw<GV�L�BfwYH���ʷ�K9Pϼ�x���-;^ik�mc�#8W;�7���v�����W�	w����S�Ud�EW���~�q���uߞ�
�<��@^q�
fy r����}Wg�ϛ.}�Ζʓ�|���;��L���-}�.h�eotϑ%���t]��+��� gz�aj[�GO���z���f�L�\9ɍ���	�(>qx����~���Rl*n*G�)w�F'�ɿBp�Ѣ��] #b�N��x�Ӑ�.ܔ��m-e����*[ӣ����8
�%IF/
F D���2����������*�N: �K��-���*�(o?�>/�dT� @}g��J�0��j:��� l��W�B����~��/4a�<GO��c�v�W�.6OmV���1�rz]o��F��Ĉ��CtrpM����I�6t2Z�3廿�}`���]9�G����'��6��M~��ە�x�F�=�/v%߬���C�=��6Y�G}�?G��\�t��#l�%6��2;\��]2�Q��{�e &��G��n]mɓ�'j�>�z�����&��ՉP������RO�9�sr]�'��b��)������������?���~w�=G� RrNV�Bk'�r�>�)"��l�X<���*oV�-��a�"���I��T�+�;���� hH�7�Pm͟�h�P��b�:�J��s�,7����ps_}�J�y���{(���&W��t�ݮ�����ƍ��mn��8Fdk++{���f{��S�w�cn��V�u��(2~� �8ʀ�-~�B��Ν犹���)Rv�z9ZNG	���O	y�Gv�t|%�"B�`��ѱ!3���}�Gzl��7���x�'ܶ��k�]F�lS�� ��*������o�a��Mh"mL���~��� ��t4�4�eH[+��S'��t�:�ҍ�Ꝭԥ�<ҟt��8Fķ��A���C��m��G�|�J�mval��@a0[�rSt�;z:�n�Nn0Iw�;��`�V�Q	;�/�aϟ�6m���D� �#D�=�4@#��^S�l{�N'.Txĕm��LH/+���^���e�����C����8Z�:`Y��Gע;�M�Qb� ����Ѥ�j�(@�X��B��gw����V������pi�ePTXX����ڮ]���
N���ڳ��C��'�[Y�&�!�q��"G�/5�l��mű��KOjx����/��ҿ�:��)Z��N~wW��+��q���������������.�����:}��U�z>=���]�x4�z���U׾g���ܥ�٫w�J��,	|.���]�.M>v���%W�H�;3t�6��q�<r`+<�F->i�o�m_|�M���w��O_���u��F]��*ݬ��:y0����K8*�)l�I_|P��&���$$?����/���{�8z�ջ�2aW��)���x�Z���μ��(�V>�o=�6S£KK>'�~ۿ�,R�I��G�g�O\JRw�F��0~sD���]`�\��Rv��;�R��v$�-H�˹t�)� �瑹'�IMZG|�6�C�cur��)]�W��o�	:X:"�玶�EО�"��Bi#D��V燏�]�E��"�������r�d�\K�R�>�9iX�����1�:��|��,~��l&��wFX�z^�L}���	�R�k?�ۅ��X����"��j�i��G^#�Cؑ�J�_�"|�o�Y͆ɴ8p�=�S�Fi�\�8��ZRO+���B��Ց��q��S8V��ζ���������aum��c��QN�e[Nl+�m8��Z�!|q��"��^l��A������y����K�f½
(G�%8o�{�ލ��]��w�:�qS0�m�]!P�0�5��i�R�����{�z�&���y���k����^�i/2K}�}D�t�fە����m~�F��d����O�q��<[�)�'_H]�޳��j��+A���fǢQ$������<F�����C5Lo�����2�^�=-06��"s�`���B [u��r$wb����6��ɩ�6>9���>5=�fg����|���o��smr�mm=;Ag�M"�%�ܹ����ﶷn��.\��&�f��ӈ�q�v��7;mu���a6��g �9@�8����rG6(*Ϧq>���8q��?�]�+m����ޅlr��LIԈ�'��6��������n���s'�u:�Jd��TQ�.n��O)�d��swa�(8�~,;	��&op�ru�e��u�|�	���	���VA�T�,�B�m�n �a[��O�q����5;P�tb�:J��Y���r���3'>�EA0���ӑ3N-�Eh
k��t�T�(��/.e�r�,#�"p�H]��ɩ�6��}ҝ��׎�ɇ<�$u�ų�KAP��I�
w�V|���0�?�����ͨ(�]A���}�F�Yq��s�JX�7���"|,<�`C&A`��u4:P�O
�w3��� ��!-��߶��J��U�v��"��!_�s�,SL,�5�Bp�?ST�`��;���g�=�Ib��;l�ss��˄Km~v.�\_�k/^�i���O�.�0�E��"x���(	��P�	PG�a�Y�I�P�"���e�?��L��.u�����
�3i�H���ȳ��/~'Z�4ٟ�������������!pte�U���_��(
�V�dy����!9y��}�#�����w�O,uX( 2�7��&�Q�"��w���c^.ү���?����N��M���<n��=l�p��?_jo^�9��̕[�}=���^�%?���ӫ�����J���ь�����;B����V����e��\ͷ�H���������,�b��#���9�+����ްw���;j�A�_���Q�J����`�������]c�������!B��uԔs{�k]�pd�K��৪���㷢OY���d��0��=��,4h�g�QBm
��e6�Y3\���'ـ��Cm6iZX�.Q��D���Nxć��(u�Qp���sǎP�z|Ϩ3{��Z��aj��>�Q �م���'N`�Ʈ�S��������?�{u��I� ܨk��W�A��z��,���Ԧ�^�o���1��̹�
��`��`M�fj
�;֍r�_�7�s���:HD�I�6�e�w������� ��Ӯ�G��o����)���������2���u&��	�>N��n��~'d�k�8���D�w �x0�M�m2���n�q&&=pz;e?m�>��R�����u8�q`���=�SXB�!<q�N���L�s�嘹y��t�{�>/Z\&��#vl�p�=�4��%�Ha������x;��u��Nօv'kj?�F�������q�&�-�=_��,������F���d�JD��Gz�2-�ŋ,�M�9�(�	��$N����<�RJAI^J 	���������j�� 2��Sf��F��(�ff��9�N-.���N���m�in~�͟[h���:Sh��-�=�gxl
�E(��0��L[�x��s�v���63�������8���okk(�㶋�:8�)�	�c�d5Q������N��OM϶��9�IZ������b���}NZvt��8�:.�	B!���݃�L��������8]�Ӗ���3�ޔ���f(�CJ�Ɋ�D��A��Gl�=q]�!oG꺀(L�{��IK��n"B݆5�en�O$(޻B�f8�(�FC�Y�sd&�&wS/�8I]�CbcD���;�R��)mH���`�vq4O�%3�{�Ό�N��p+ǁ\`@�QC6CPЦ��:�<T9�>�s5�}zh�|�T0�Gz`Ҷ���r���NO�DH�!�8om"l�~�a	=���sv����l�l�#~R���*��BJ���m^��J�PF����ֆ/�GR�ِ^P1S� J�~�ptH�(�J���9�ӓ���]4��Y���H��+��i���S�V�X��烂2�Y��0�ӻ����u�M�;G���w�s���W����͛5��U\�(ʂ�:8|���W�޺Ĉc��D˷������S���_��c[;��D]�Y2v[>��������֖Q�	���]�|��z�?����-���s!���	-��7�u��O��W�ϻ�P����YGs�7+y��S�&}��r��њt�;?�F~V��"��ҳ�`�~������ S�9��N1����H���A6�}�;�Ca�o��W ���|�07��s�t��������������N���/�����Ս-���ޕ�pY���=��m$��i��3�.I�}��4�Ī��2�}��ʰ�^b�L�z��*v+�|����5����弐�2��$�p)��Q�4e6�Uv�k|{/�ɀ!L^nFq��k�,F?�L'�	ɧ�)���s�W���'v`-��C�d�x�@ָ~
̑9�8�L�����a�o�tAR����!it|t���x��޳1���}��R�:����E a�Mc���u�
҈a_G�F�C\{l��p5~đ�S���q�ϲ	t|ߩ�@�Nց��ɰ��Kg���v~贏iwi/�7w3Ύ�2 8�ѹ9l8�z�[�k��1� ~hP�xl:�#\S:-�v%�eX?G�t�БV��#7Ea�}�ٖ�#���:����=�N�H{���g� x0���t%l:f�G[�";�'�Mz���Y˙��ah|�y�M�*l�3أ�"|�?�!6�B��Yu�x���Yl}�*yU>��!�LF={��4S9�<�d�������-��W���ɱ����5�un�'��d��O׿�d��k�j�Z1�A�O�`�٣��hq���p��#!��R(�J�d=�<L��ƌ@P��F�'��թ����,Mc�� ���n򽌽�?�IF���L;~G�r�~�j�z�z�x�b;�B[<��[8�����/t���"�4L6>�����fg���9�^n��\�"Ԩ:�1�k?�����֖#=����\�\��Ն�]�t�����
�868Z���Ӕ�TB,G�H���5��g.��YZ8�����0O�W��M��#hNM��Ӧ�B�h39�<�t��}�s��4Gh�9��N�́s�ع�I�11?`�����.����>'��"�8NZN8�<�]�K���z*pu�,o��wʡ�ƺt�����Oş|:05t\�t�2�ceZ&ww��=���9p��HVũ�D~S��o�n�
�$eFA�@���WH� �'�a�8:��/@��.�E�:��8Q:��|�O��t�63G<�Q����8�(�,Nw�=��J�'�Ipk��q�-I�1�TٽN���N�aʬ��tDYg�'��FE2���|T,1<�e斆��Cd��3Z�y&�Y,��ƌ���{z��s���,�~�T%:�&��!�B�>��;�~0�q�4+kՕ�%B�6��]m������a[]�hKK�s�4��Z��yT�^��o�ו�����_��/��G�����ϔq���w�����ͤ$o�����������*p}�ݷ�����A����j{�G�Կ�:��F����������2�����s����5��ݑ<k]��5N�\���T�͈AC"�ķ�t�W0x�,��(��B���9$��r�W=��W�e��	<u���9��e]g����[�6M��c�&�`)'%�gI���[~{9�S6/R�	���v!�pB���<2��R�Iq�4�p��i�Cӻ8����h�lF�A�y�zi7	�i����iҙ/y҆17Up��7���alGwf$i��?�3��+w�Ʃ�|�8���%}�:�����':2:8\�*m-��� w/��\ƣױ%�&v1��1_m��~�w��IW���W��H��v�irL��cU�&��Rt�~&��Ym�����H�b������6�Mg�B�qrtb&p2l7�r*���2
B<�G}�O~�@�8��o'���x�p��a�L��i��3�S�l���2�E:AV�F)���2�e
\���!��sj�N!����l�$>p�J�������L�$�f<��v�l'��T#YP0��tb�w���g ��td���/t4E���q6���gI_�hZT�Tj�؞�4Z;��u�2.iͶ�C�K���oM!�^���~����8��t�-?�wNXd���{�;)켈�5?�.]<׮^֧�j��N�#Y;�&��R{�9Y��fH ��E��NH�2�0���E�|c+l"sX㓴
'�ʤ�ƲN���=iz���Ù]B����~��b��:̊����67V�h	.75�9��/\8߮^��n�\ݼy�]�~�]��*k�F��/.����T�I�:6G����( ;J�x�5^1���75��F���l��4��7;��ti7��T�f��X�5�a�A���:+::[Н�S���q��稏=��n���::I���Lc�]��<<iGD�_G��q�t�D��)�:K}�ɛδI��ټ\��G�k��,�� smv�\�����`%=�4�YG��8X8K�:?8�2�qu�FeB� �(it�t�t�gg�QN���R�� ^�̓���B<���9�(@pr�(jP8����йM�u�N����yʛ�����
���(幻fbZ�S's�43N=�l�#���2�Ϧӑҁ;��ӯ�EX�y�rsP5�ר�Oĥi�;�A�f1�����x*N �Qx�AF�'�:��#m�{k�˗�^�,�p�Q��^3���ִ9n:Kq,��9��V�N��H8�d@�a�ę
/W��Q5������R��N!CQ���4�R�
K�y
���4������Wd�7� �u�m���{�r�T�s��9h�)���t�6�+8Y/��۫W��I�.UZ�����ga��+X�΄�W��.�Uu���\���:y:S�Y����[��E��O�5��W�3��-�}G�5�y��O^���2��<�����ŋ���c~v������ ��L��M�6�G���E7I��e?��[���<,Z��>����Z��s�x�pU��di��O�d ��̻�%��3������^�,w��O�L����+-��q�K��
���?���:I���%��BU)�vF��eL��di�	O���g9�U�gZ쑠,�K4;��|���ܽ�>���w��+�md�=�� 1@ο+'��ձ�n������X_�.4�����A5�����h^	�K�
���%1���kMV9Yq&��F�:f"QcVz��F�#;�J%��p2m����q��+��5�k'`g<�r;F-C��ߖȔ7J�3@|�HۘƵSq
���N�l<�	�gd#�&�������5�����3t*���n��Pi����x�#i�gT�:�9g[�����ҩtdJ/�[8,����8�|j�(Ԏ�!pTJ�ߑ27��=��҂�Mk��'����#z�I�q�n}����x�#p��M�
:�>;��i��=�h��r�t����"a��WGة���J���	g� ���W#c�z���s
޸[�1hA�����*���c�x�l���,K��mt�ě�M�M�^�H,�9I��,��_KGPj�,ˑ��Pqt̼�_^i[���R�����.x�¹v%[���:Y?-'�s���l/_�����;G+�Z����d��5�V,���1W/Y��!2�]�ʈ�#�湳��8���)�+������$� ��08Xk�:��+d(�٩��/_�ɺڮ]������<�&^����TE�N;�8��u��%P��]CPG���@� 1b5��]X|{muu��Vp�����F���&�N�Ɏn����ye��9:S�1�{�݅�w9\q�t�X52�񎣠�ᠾ� ǘǮ��4�n�+�t,���6�9�����ұ?��M�{=�_��C�T��]9%��o���EȤ�8Y�Ε��L�&#�c�<�'
���:F�)���,�F�g:d��ϨO��rz�F�K��dbFx
��|�t�tVm��B�������o�(��e�a��
�n���5��cFY:F��
�6�R�K4܉?n1a�L�xNspz9X�O� �?�`��ř�����)�<R�9���f5�g�k���{�)]�Su�`e��3/�=B���	0��C�(3�Su�����h��=j��S�#Φ�1����,��c���Ĺ0:cʊ2U21 x�Q�;ڥQ� f�3�)C��5�ӌ�=��W>���@ ֹz����t:a.\��.�OC�m{g��^Yi/^.�e�,�����W8�YX@���$��5N���N�=y���m&��R�]��X׷�Q���ǃr�G�ay��B��V���	��Gߟ��s�b������� ��/���믆�۷ޝ^��l����h��V�.�s}I2�$���W]��:@C|�����aӎ�G��)߼L�����Li<A]�x!l3M��;����Eɱ�W��&W��r ��,�S� ~�{ϷI�%�Z� 0��Kַh�X�o>'p1�y&V�"�*���|�����Թ��/5�Xρ�#��)w$�fZ:Y~�{_�I�yC����e�5��K���3���$/��W�!�ȣֱ�.�§c@�;S������E��^�Hd�r�:r���cෳlGJN�&��>u�hT�h��q �~�B��z<�!!F��6Hl-G��D�VXm.G�zGA'I[ ���rYXsV���|�O���`��/;as(1N���8QF.��n��N�˒t5�c�:�QgN'�Fv<#�o�;����f׀�����Љ�:��gm�NڲG��r0z�����[�����w.������Y[[{Y�)�I-l�ܠ3e����)��gշ��)��)��Ӵ��A��	��5x���l [������Lp�f]c���N��n}���j��e�D阙Fg�N�����p���l���֤9���;�0��_�"t��[���;��ͭM�'���M|K�:X��y�/�f�*e,cǩ�З����V�M��m?9>�uX�.̷˗����ck�=��Z���0b;@r�,2�h㟽z���K�n S�[TO&�֡H �"+Ï����v���[ u�<J��01�9���,ojr��������yh$����N�ŋj*�B/�+�K���9c��1��8{�0�1F�>�m��e�P�Q����ﶷv!��&��]ls�t�A�C�nt��@ڬK�,�`�x������U�Ҙª�����tq�$��/%�;\~�G��0�3����N�7M�}��8�t��L+S��>�'�C�eg��nH��{a�iU���Y�q �'��	�.��M�G|����#�ԍޕ�1l:ʎ����DZ��	с('�~[#{3�7q/&��8A�Y
��ʠ�I��l���m*GI����Wkq�S��:4Ҷ�'�t����%��uY����1+��7����̳y(����M\;�΅ө���k�qLqfu4ŝ#���-g^Z�P6�b|�uT�0 u.�@�ԡ�q{����X!~5ȷ���Y)���!U���O
C��&B�����#��z��M�T"��{a 	y��ژ�!ς._�Cc=��P�1"X����=�5G����D�\���W��I�o���W���8Y�Ȃ�٪p�?a�N�Gx��zv��2����?��_uY�z�N��>�d������"��~�������?N.3������XI{p����\n}�u��v6�*���U���N���6��A@sb'jů�+A��>�EĞG��*�c9^]F4�t[y@v�0��g���/Q�FڞǢ�����y}�Ѱ�L�U(?�OzI}�F��?�����w�6���)����Gq����o�&b�gRԽ��#>N�A|�=��<w�E�ir���"�	֯�'���lxD�|E�L��ߏ�x�u�V�ӦA��DV�(�i�_�J�<�M�����'��'~zcR^6��׎n���HݕR�Ǔ�?�6v�%�#�רU�g�����˔Hℎ A�t�r,�O���lg�D�[G�%�v��l���M�c2n�Z�`b?�����9?�`�1�SP�m$҉S��ֳ�S]�y�;�[ ;2�]��Ѡ�8s�*�u04�]�-f��^�i[�#:\�<�d� boRVL~�S��3��\#:�B�����-�@���\�F�82\:=����08-N|Z��`�/N�|�]�E���Np��8:L�"����8{%pW�ĩ�>�n���i����>��ě��fN9�������ea�g��:Zw�e�k���;uvc3�,�UmAy�Í/�[�qř�Y뺍�S�V�y���Jl��K�����-N��޶�8���"�������K,����+�$�:���ebl�-�M���e�yG���V���-�����������������Ͷ�EV�N��0%r�,�;or~c�L��v���&����Y��I�V����vr齃!6*���!F�E�kkk.<��� �� ���Fn�8����wb(ö�0r�������	m����W��[o���z�F�Ο��x�0���;�� �	"���P{�B�o6ګ�[���N[��qrX_b#]�"D$���W]�r�b��+Xb��p�D,Y"�OG�V��䡄R1�'����%���\�7�RA����	'ϊ�b��<h�o��	z�6.�%f�G �ޔ�ۗW��c�TH�����u4T
�r�<�m+�w�	h�����]�h��F@��o�������-�3"}أ1
�;��t�;[a|�I|���m
{�2wH;��UJ)HI�0�� �-V�������p��T��]�Au8(pܙ������(�l�����o�QBT%�������@bv�1����e*�]y��w�΄ݝ����¥��a�Ys@��?x�Kԗ���)�_��ml��>������TVO�㝽Z���߱�T��v�ه����R��E��l������`t��U� +vv��8���nZ)6
�Z��� *ߤ52 �iOy�ɢ�ܺ�~�Ïڏ~�q{����8�=}�>�����_��}��ȍ�Ȯ�N�{�˶�y����u��9��;�������(9qN�뻿����r]��V��3�UNKQn�0W}�.�fj�I��W����'���$�?��zW��/_=k������������)0!��7�|��H�>E�W������s/_rK�£�~�v���i�>���1���i���%��T���t�'��̂uW�����e����ֻ:!N�����r���<N�<���w�z����4]:��W�b���^�(��H]���9�� �V��.z@==��p}� N�@ɦ�öEf��K����U��.`��^����NO*�sF�i f���s�,�v���o�xe�F�~�\ڲ��,\��9r9 d����r�4^��x���9
]�zZ��;�AG������t���v�V���ף:c	:��/` �ΓӳFF�����iW�q�i��[R��:Ru��EM@���ȋ6G��d�{�􎛼�~#(�Iꪾ��v�,H"3Rt,�p97����8��v-���;��"�[�ko�A���~�o��I��3G�m�
�h�_b_Qo���d��?Gu��?�h�#��;ڰ:��:Y�I�c?y�^BzQ����Z7Y�m������K:��2//�`6/Gvt�8���|3�H�X�� "
>��X��'�'���)u,m7F�oq�Cf|���#ެ�N��$&��i��,,hR��N=�c�8�Ni�DH���e�8s����ڃ�$��"��O��H�Nq܂N��N~![�r��>�|���l�������+���~���ݷ/������Wvq��q�~�e������{8Y[m�u��8#��
���t�F��{'k+���aͽ�������"�W�D�{±!���c��N�J�a�.����֎Χ��wp�<�cg{#�j�,�rKH����;q�t�\��n���Ef��9��W�Ǵ?�a{�1�ެl�`m�e��zu��m:K�TG��UU�Bˤ'�y��3�oa��8Y%�R2Os��B >9/��D5v^{_�`�F������Asr����|��I����T�H�/	R&�	SB� e`ۭ7z�d
�y�(�;�i��.��h�h=�q�¸��v�N��޻����`PП::��q�p�)=��TxQ
���&m�X򔎃N��}�I��3��Э�{��[�W��X�r���I�!�B�afi�:X�Lo ��*sp��ҸҼϲI�
H=�9�02�p����7��)���C�t�0�����";T>�[�" _\�JxU:��'��o�uI����9��2��}HQ,���W,𿇓e=�$-'��Eh��
v�^?=0�4�n����Sai���"�<�6U��'���t�~z�ɿ�o�tc ء% ��c��i��~��8X���λ�BOۻ����������i��r�Mzy �څT�RҖ��g}��suxP)u ��+�\E�ً���r�v���R�~��r+`���ʖ�[���s�M���og��5�_'����wu�޿.�.�30��[?���/]�D�땺�_W����9?��`\KNGh�ה���^��u�J|��4OZÿ���c�Mˀ'rƺ̷�B�Ǔv"B�U�rR�3W�^�ힺ�?L�����l�+�Y|�-���E�[0J�,�)���ϼҠ3R�(W�� {��"8�=8D�j_�8�ɦq@�Ț8(�+�Xl#�m~;VH���NeW�^�K�"����wn��ov `���k��xgtŶV�9�K���o�U�k�츣0p�ѯ��4I38�~�uKDJ�q Ե����>i�Iwzvs$��]t��ͽFGgѽ��q�� �z���	�_�S�G��:�B}gEu �F W�Ӯ�u��`u�Z:h;m�thp�n����4��k;ќ�&.��):lꦚ�_�둸���:
83jE~h#LQp.�X��DI�s�caY��.v���$2J}�~Aeő��u��� �C�=]�Z4��x//zI/:Mq�K�!�M�ҷ��mUv�q����O|/� I�r*~����!��K. �0�bW�p��:��~���?������lR��g��O�[W���t#�*x��.�ԑ��i���6���c���U4kR1XS�O|�e�2��"��r�Ӿ��Z#���]:hy��� �g~z���c����z��+��|�d�#Y��������,R��K� D��v�˹i��(V�p���[5�EL��1�jF:�1`jƔ1bt�`�+����Kd�dI02��j��E�-�nﶍ�M`�Ah@h��嚫�7n`��n�}�]��ZX8b0�a�0$U�9�I�@3;��[�d�ƹZ��z�F'k/#Y�q�hd��,"�KiejK�鈊�z�hm<�2M�6���t:�?��_!�3!�W�,<�����q��E�>�c�K�|.�5�)gyfkܔ��� 5)�Τ�ʨAPB��:��A�4��P^~?	�q���z�΋�<��pJ� �+�PF�k���թ����^U}l#q[�>���ZCH>0\�Ҩ�����N��6�H`C0�>�f���!�]=��e*@�3��x6��U���ૄf�����ҥq�Vx�:R�)n���2�^:_�BQ�m���N(�Xg�G��=����|T���m�d~�\��)�2��AY�R 3���&��N��I!Vgs�'>�?�.�����NX��_܀۠��l	LɎX o��c��u�?w�Ukmm�u���h���ضf(��ly�6y���Z�������?��ߴ����{}�nܘU,!�s��/�����'N֗QȖ�;YE��TT���(�hԒ���>�OE������:�O_5���]�\'����*�<z��5�/#F���{E��<�>������ī�/W�_ʨ7���,�Ig��]x2O��S�N 9�Yw
�+2$;�L���>��w'��"K�zJ7⦧52�{��^yWɨ��L:g �h�|W���������c��H>�\U��\�O��E��=��w��qY0'�3W����������}ܓ��+xȿ?��}���(�34�A����8z �=95Ҧ��TSΖn9�A=�Gwa�{�'"��8⎰�����n�9�k}}����D:�T2Ü�p$@(��D׳����nkm3�L�"���e�ĳC��l_�@eM:����ma�lm����ѯ�2*���7<�A� O�>����y5B������ �?�͌&��i�`���i'���:t7���M�ӄ�އ�:���MQ� ���:�:Y�������i��i�����1�����ͪ��x����X:?vV��o$���9��U^�_�:뙤g`�|$Й5M*b�|�*��c�ɻ�&���(����d�6nl��唳�ly���~��v�m�D,�x�Ë��8�Q�V�cg��b'*.�[I����1��8=����G�<F �څ�YٓW��Ӝ��(����iGi{;�Ň����6O��)�1�.�������⏴�C`�q�l���|�e}���&�q�s�So���8<�ɒ�h���vnf��wv$�+���p�.'�����j�Y�d�����E�5�j$K�%��ɉ6;5��a�]���uG�`���.H���VE�,��C^�#d��E*刂A�3�`�V�Ew�Zi�B֡�+a66���se/�B��\���~��L�t�r��s���0D$18�$�y�f�dml��k�&���s�����ES��%�{��!�E"<҃*���5B)XeŐ�v�BBq0���g�0C��==#f�u7a�}+�@�Q�����E`0�uH�;��%1�0���7���)�%yJ�����J�m�6�2���wE����5�D���
g~�8^�s�ƴfYeh�������߫�M�H�7a���-G�]w��� ;�Lk�fY˴�RJ_�TZ:Y�!2�c�R���1��������YN��-�dn�&�{`$U,�t��[	1�4�3�&�g��F|�Xt@m�G�
7�92I:*�[ȴ߃7���6k�� � .q.N�i#�5�8�N��S�㻽l
oG2k$KX?���v��!+��AF���W����Wq�<������6�S)q��8
w�H�]�-x?|������_�'������v��80�d�o���~������?k�}��ԓ�����u�hq�BۍRux�H�i�ψ�eu?��K���K|$�p�2����ۙ�s����^ف�L��o{8�.�VC'y-M��o��? ��}�G�M����~��_�����(ͥs|��o�r�}��nE���w�����?�
V�v�U�W��M֐��h_�"������;'��* ,�T>�3��� #�qq�J>\)���UWj���|L��g}�<���+zDx���l\�}6m_�����;����s_�,eq���8J�@���Ni�s��s���s<� �jV�S�6����㔲�	�ӌ�!��v:��l������勶���l��a�J����I78B�Ձ�c��T�_/�i/�-��W��_v
���y��\��C'n����V��L�E��"ln��m7`���qR7��1�	��C`ݩMzSv�d�%������M';��l�����z!nY>M����	+�˥L&��_Tc�;�H{�F�p����d!��d�`g��#2��RQg���H&[��Oh�:+�]���@�9S�k�v��cV2����{���
�������p�#�YnxEg��g�7�e �� x���;�ގ�9d�e�(K>	�l����_K�}�W%�Y��a�ݫB�����ʔ��}�;C�����Ȝ����|uz9ܵq�m��/�'i�*0���r�Rwx�2t�b�P~��f�n�*�N�m��N��&�����E\����������U����c�Ni��x�H�G�$!����Cg���I�ɺ�'G�u�F�é�8Y�H֏~�n���w�{�\m�q���h��g8Y������9Y8�d�@���r4�邳�18�^�5"������w�;�� ��?[���P$XIrt�M�F'(�3��7<�AiCQ��8X~r��D;��&��FS�Ϸ˗/# /�������Nu��I�@]��ߛGmy}�-�`--o��7��N���A�Ƹ�,�^��"��D�NUO�>۸q���t�-����5�֟����6��+���g/��?F�Y�w.�K\&�3��q&#I���-�����S>�*��;�Jf�>�W_�N����T�ˬ!��̷C�*1'#F
"i��n��4�MP*h���{mSe���QʳV���l�e=%.���3�el��Fxq�CԽ3O�O8�F�}\�^����VZ1�W���'K{X\%��Jk��k$�Z�@�rtW!V�OXvZ.x���P~%+D�C!�I����������Q�
Sh����FgH�A})G�Lg�IK�d�&Ȼ�De�;q	�i�/q�p���N��*����/�E�d	_z�'�K�@���/`��h�+oڶ#Z�#_{:\�'���!�(�L��A� 88Ba�M�ζ}��/��O�?��ݸy�-.N4wu��;�ﴟ��_������}��ϐS��])e�QAm]�(LA��"��[�u�w�R��������#�r�J�.��s���(���k|���t���OS��q��W���O[�����5͒�<���*3#�(]]պ! v9�743�p��▸���<�!Dhݥ�RgD��b������]ݍ����������ݏ�7��;q�_=��2���~3���Q_�WW�sq�]�Qu���2pO���wB����l���YP��~�󫺦��)��	7�!cq;�,�/���E�`�������o����eL�w�Q�7�������p½����2�Zi	#J�3��&}6܉߹��%'�񳶼<��޻��{�A{���q_����w|�|k��ze����xO2|�7�̐{O�>o�~���^Bۓ�㊗���]2{>3��b}�����=z��=��I[�
�v������א[W0�<����U����W�FQT�ƈq��z���'�vbpi 9޺J�����	�� �|We�����<��|��+߫�c�7���׀W�V��	�K RR�Q�j�-���<���M�kR�]���='U���Ġ�c���r��Um�m|LG�zt>&ǒ��E�Bf-��c�!O��Ex'�yI�K��I����\4b��U�*�j�<��ɢI���1�j~Y�q�L���IZ@��b�b]/�ъ�IP:��O�Ў�ѧ̜K��i|��<|NX~�E~������.����l����d|1�Ĵ�
 ��1�p����5�\�����_Wm+'VkK+Q � �O�P�F�yZ�}E����W�	d�K� o�o��F��Ը�9���H<ʓ�ʟ�I\�<����+Yn��w��/F����W��Y?�%F��^�ه��ȂK4�v����s/���X�=�����Iˤbede��������MmO���uu���)�5?;߮�\m7��hw�ʡ~��͞/P����2��4� _����^�<���=mkY�1����
��{YY�"����m�F*�0od/�G:��q������o�@������x�yh�2�������m�������_�^�y��ɧGL�v0fR�V���TLÓO��J�!;o-�����Q�߾Hڦ����Ψ
�l'���|p?i�� �W33�8��0B�i��5��p�t��_ջS��l�ȇvx/�}������]�G���*��-��O�T�`^���<�ĩ�4 ��6�_j��r?9���tO�a�������"@sQ2t˖Hh���Y��*P���t�j膠�Y&i����rIZuI\���c:!UO#vSo�2��@�A}�W�W}�.���e<��і����[X�G{mwo���x�^bd�z��v�721s���:AF��PT7v�<D́�m�Dj�ȓ|�������}���i��V����@�I����O?o����M����_�����%� ��V)����d�N�!K����]�Ԙ��pn<�[�o=˟���<��0���}q�)����<���L��eMUά.��UA����4D�����{�L3r��tU��wE�x��n/՝ڕ^>���6��=��%����Ҽ^�LHt��y�P�2��G��{9��x9�?ʟ�);�T��H�*�*K���!}�wb����el|�U�����te,�����(���K{�����e>��C�M��Axۗ������>|���[�O��������;��G.��M��ɬbmmm�+!�)�t�K�3W�rH��2N����	�mc�1�o!����3g�3"sl=�#������'km�٫��s ����L�%_�˚|�$|#_D�;9��R�[/��dgok71������ϡC��ܼ'	��\��<0ƈ�.$���t��%W����O�����������W/S��d F��t;d�����Jh�C(�����9��$b�V'��UTcL�8&�~�S/:���z&���@޾�%+�!ŭxƷ<�gW��WJ�	�85�M�g(#r��sx"[SPȚ�q��<ˣNRq�2�Y�\��mbd�F�H�L?m����N��u"��Z�վl(x�\~"+~�Z�bS��WҪ�7h�_}���k&�4�B��W�q�����7���5�������'�y��ƥ?Y�/�I,g���F����c�4p�z�:����4��u�I�gW|	�W�I|-%x �Mhf-�Rm��C�P%���f����� �4��-�]Е�;YɊ��ޝ��/�N�=�h�忕��J�+9;f�Uﲠ*�&ۂ�{݋Le�}��v0Y�YT��t�#�\�uP�H�c`QI���QqU�ܮ#��qu�j�vu)3G��tr��=��s��km���v��ͬb�]��t${B!����T�Y�����/e�}�v����;i�[�ڳ���ًm�������w�v����	&�@��D�Q7Kl蒙8�g�=�ap�����X�G�J��a�T�I�}�!��e�49�L<\�5�q�G��tD�'�ߐ^��+�"C�W�_��WUx�g�g|��%�����UI-��"�åN%t��4��$�#��*�@�̐�#��6�ǆ����"�.�s:
EtH;�u�MYtr�d�#�Z��TFVfv𹠁�x����|�x����T�c��_5�Y}	�Ĭ��NW�jP��b}bѧ��ԥ�u���s�bh﬑4I��+�%�hϡ�Y�8Jx�.�O�5�����)!Fz�b|��?�]�+ڍ��g�&�9�v�ӂQA�ns���5u���E���Wk�۫�(-�2�񵿿#�-���Cg?��U�z�5ѽ��9K����{�?��?j�G?l�A�}�Z;:8�b�٧�����m�W�~���@O���ț�<2��%�X/˰M�X�4�7^N�A�/q�tpv| �����ѳ�Eɯ{p�wQ��T���1��]鬻Wڳy�W����|*�t����ﻜ���^�3?�+��C�q��}C�M߈�;������5�+%��,��Ļ)�|T��91T���|�t�(C�a�"U��+^�4�e��K.���0�K�s���e��^^%T2�m���
�"��G�7�֪�W�7�B��������Wշ��i��t�/��V�$J"��˙�g��m��_������?o޾���G4�Q'��&��A[�J�'tS��,�0���t��;��nW�
rќ9!���	�r�mc��!O���1�N}�B�z���gyW�h���4=�A6�a�!�kմ�Ólt�t�����⣱55]u�.�]���a�wv���Y�9�#������?��k?��_���M't��e�^@#tB�;��'����0�Ȥ%u�Y0�bʬ�Y����ģ}ڎ1\�����sd�1���c�u��<�B����mg�i{̑F�-�E��D��1F+Y��
� �5���}U�5�5Vcl@�q�iȝ�k�8:)����Ǿf�$X�Rz|mu�P��
>蹎+�?'ҁ_�*m;�wëҁ�8�[�>A��j����i.��s��<{_sa����m���� Y�!���ꤣqjh2��.$ue҉W��I�,��9V�G�R�k1���IO�j;Ki]��R��-~v^��:�����v���{��q.�K����/��?��N9�g��[��#2�|�
/����w�j%+F�����<��������/�v��'/�W��ahl��*i�Ӑ��0Y@b�R�8	���o��C�{P7�	qU����Yџ9)d|�ʏ�����q?��S��wn���[�{���}��;�[��>�ֻ��w�g���w�;wn��ׯ���n/PeLa�����QBI�4��+�!�u�z�����x����=%�zg5�+u�6C�ӽ�4�����!� �PA�*�;)}�:�R����MX)��Cx��W���0����ØF�/_X&��K��ƫ߃-�G� �����Q%K�r��Pa�g!_������t��O��G3�yU�����k�'�8U�*_?�^��K'��;�*�Q�Mk����~�u�ί \aSP�ֱ!G��o�|D�%F��e�[ ̈��M[s��&nܥEh?�'��*�V>	�Mv�E�:n](�Ⱥ)�|J0)8�牓YR]�\m=9&y%�x�S�:�9@��\�J�@�W`��6�3D��̇U0�Eޅ@��c�5��a���ll�y!�0'h�ҿ߿�[G���TNܾs��j�q�z[YZ� �`���z{������㶾��2 �T[yeV�cX�Y8a�Ryr��G�QJI�|�����$�����m��<�x��@�O���>V^�Nɗ�K��3N��x�/!	�_Ҙ_�S����?�D�?8F��@\_{��a(�/�����Q�����M�_��G�Pϩ?��_yg�z(���r�2y�'��y���.uHxh�m�<��q�'��x����D9#^�}��Y�w�_��͐�(<y����a�^���ĭߘ��Fq��O�$��DL俔E6��֭���w>l������-O�#�Ep!��+G�LN���.��u�ᬻ2M�m~��(�*�u�v��L=�&e�V��e�!߸�#��ojYvy�v��(]ď�����x E�� �4㔒i;�r���l̻�N����t:'�<\*���v
�k=g�.�;[3�_�c�5:=�	<ɩѰ���M�³����
��^�j-��1�`,�wcmww$�c4��.W4�\yY�:JC�\'��F�8�vI�]'��Fo�m��R|�������U;߻�qEN�;\�� ����b�\-y�5u
9(��w�݂�F�9ilL��r�q�rL㊘bx������w����N9`���r$�4�rʤeQ7��ԍ�u�s��w�m?���Ic}lGZzH�����n}�.�C�7m݊/ms�F�����¤�8��pX�|��8և2|�p�:���j�ir�>yI�zo[���4�ݙfۺ�b�UW����u�Q/�~���O9�/��S����V�kEY=*:4�r�Lg<�DO�'OV�!:�J	Tu<i����kK���;Yׯ-�w�`�Y�;����<F�^�,�H�'V�����A��bd�����*������!,g۝�UxH0�$`�����;k�WW�?l��~��oc�o�jo�u�ݺ��nbX]��Hz=�'r��f��1,/%H�9f�P�h�(r���ֶ1����.�L��PA�VA�Q8�`�4��|2���qEٖI9u/FM�){�G]7@���Z����3H̢�x�>�{y�Q�0�)�擠�]<�4���/eT�p����{'��-O���7�R�)I���\v��E����xh�{u ��Uq.⍞�/�!]� ��V|�:��Z	��Vz�j���GA��i�ǐw�?FV�5,��x�"l	��Sr��a��eX��2��)��%+G�uN�B�q��S�J{~Z��@�Ocbdh�W�y���3�
@cgH#���G����������)#aeP�R�G��4qu��5�����B��v�uw��	����NV��Cl�SG��r�.����|>��ʗ��3���nR�`��
��V�s�v�ze�h^���ٓ�1��^�#^������e+��{�A��;��/�=Wn���-��rN����} #�#w�%r�g������� x��K y�M��H��*M�SqM#tŸ+ǉ�!� W��F���E����ט�ϖ]Ͽ����~%ɐ��i�J�CP��&\�F�^�N�T=q�W݄y'Q�׻�|y�sO'�p7,���'ωT8X^��iY�1�Wȏ��E�4sx�
1�*G�<e�=����2R����	Ý���e����ʏ�'%*��4���z�W�A�	��ſ�j8��5�WWW��o�oo�{?�)�y"_&��~����̓���V{�t��x����ll����w����g�t&��Fv�����\[��?�!\kk;�9�_��cg])M ��cgg�|�{�^���W�ڦ��ٍ,+9�e�rW�a�!�	�Th��X)Gwv�I�A���C^��E��n^9<:�<��TY����J�OT�X��%jm�4x�-����z��^�$�yxV�:"��Aޮ<� GIVao��ʘR�s�w\P�D�D)�1��2��-���>K���}�?��2O�/��iʆ�k/�Q�˹�C�0�� XY^�k\�4~4V4Ǝ=�4(��o��9��y��v��0�@����t� �[��Q��1��Ӟ�8���z����R��c&�֝_WV�c�O7��K�p�s'�)�����[��>t��S��U�Q�d&F��j`yҸ�jd?�@�NY��{)ǌ=Heiy�͓Σ��)am���Hd�I>�Nɳc����^� ڐ�F���Gy����1=�_^X��Ww�D�0ˊ��!\���5����b�N�������#{C�,�������έ�v��*�b	=�]|�mV�v����ۗ����/7�|(���ƃ$�d����;Y�q�Q�Z6T�@$9��K�Uf[Y^�����a�{wo�?���ۏ��X��g����a���9�0pF�.3TT�:{0aZ��$N;�q׀Ou�C!j]���ZV�4�d1���!�w��\�'/�[q��)O�[g;��[CTG�G� �c�S����5��4�?�[|-'� �w��cz�p'�[���w�/e� @��C@���L4v�ÿ�O)U>8���9��OA�mD@�sDL>����+ƏqC�x�jL# y��(Ӫ��2d*�ʭ:�~��^�*V�)�� ���v����g^��t�U�{��V
��۸���Àl��U�dCe�V�e\�������KnP��M&U��#ys7�ܝ����؍�ػ���XlWfu׀\���0�R����[["���G~W��Ú�(c���=�>E+��3*?��|A9�9�Y���hh�W1��T)x�v��8�&ʁ�*BٙC�P��B#k������嬧��`�En��-b�������v���(W�'�P`^<ў<~���Pc�R�}�Y5�͔[�;_֝,Ӓ���]l�ۗ�^Mϕa�{�<WX��{¸���=��6�����E��Jݽ�W�
�mC�9J7*�4�?� 
��q�,�2�[U���<��� ������M��;A�x��R�����8���d��5���1<��.��m�
�՝�o��/m�_������FhH��ͤ�p�r;�9�
Y�?q*�?�X��i#��!�j
��޾<��r� 9ee��;��A�[��G�k<�މgy)S�!N���R�6�Ĩ�j�=��Qi�$l�:�8~�f����7r��2�����X��`���9jO1�>��Q��/>k�}�u{�����������z�ϭo�hk�^�g�^���z�>����'�}�����ڗ_>���=z�<�fkSCk����_���Ϟ�'O������ٳ���^��͍Md�ʭ�7#�5����^W=�S��앁����Ã������2����^alitml���W�\�iܒ��Q ff]ٺM�[ՙ�s��c��׏�K�����h!r]���f��M]��"d8��6��_����W�4�����U7Oi����%��� �%y�/�x���?�vn�s�)�/lv�Uy7i��	�9ܫC�RW�����plr�Q��S%o��k��Htߜg�7f5��3?��ު�o��=\�:i�Ջ�����K��!�i,[��0�GF�_����d�~}D9��L�Y�2�܂��I\��]�>�r�6u|���B߷�r�$z�Ɩ�R��Ls��d���e��V#˴���;~J����;�:��H�y��P�_�����X.]��Nℶ��-�'Q��9��pW�����.��Hy�t�Ke�}Ŷ��%��@}�2��C+�Ϲ����*���F�;�dad}�x��E{�����0�FV���Y�Y�ϋ�:�Q��	�v�|[`��q���uP�.O�����$�X�[��l���n������߽�F�֔����4G����B`=Ɍ���
�G�.��]M:� �8:;�i2�>*Rc��]�+'�9<Byڛ@x"<������3�
O�U���h������\섴+"��|�P8�[���!D�F�s�g(i�n�KƦ%��������@�m��n懟��I��:��)��8� �RV��2�7�G�o��s�Mɯ=�����zr�퐞܋~p�
��*��ա��l��~�yY��2�3��b�_�����A2����M_t�'~����i:�����0��8h�ҁ�@|ɜ2��v&E���C���^�vk������;�T��j�p��q��o������xN��*�a(_!�wB�҆`�\]i��Y��Z�<C� �	������e(i�YF�ǵ7nH��gW��<k�1��]�2[OA-n�(�[�m{s�B�߁�8�[�<�\��p�M����%W��#�SI/1�j@��m����-28n7Vo�w���y�~�qc%�:]q�7��W������mo;�mꄉ���~4j��*u��C��+��G{���	q�?(�m '��#%�T0,԰�w��0�Df��KG0��q���t�%oq�t�^@��Y\�ɟ�oz�q� �{X�TDŉ8��2�*�2��o�$Rӊ[�ax��e��a@?�+�8�����x�X�� {q���쯾�} 	�䥟���7��(����[���r�x��땺�ֻ�j�z&�$�� �����&����ÓvH�	��<[�	��ݽ-K��]�w�Է�\P�(_Ȟ0����L�p/^*<;��
��o�В�Q6q�'������ ?U�֚<3�<�6ܸ҆�[���y��y;�:yZ۱�s\��;�n��&ڭ�7�[<UP%
=�����Ρ.�a�_�������_���������@O^<m�~�E{��	�ǋ���ω��}�ۧ���}�����o���y��ן������ˇ�ۓ�/0�0|��1��Dz��F�����_���Fq^�od�� e53�����Q��m���v�.ak{#����g���%�"�^>k�k�1�^��Wo[�o������Ӷ�j�mo�@C/W[.g����Xo�x�/��\�#�5&��Epal�I.]�F��n����#ߙ���g}o��;5.#�F��Of_p���!��8Ȗ/�荦Q�ʇ~`���xy�H�A�b-o�9��qbrj6cEm�7�f<�q��g�5�y߇r�f�be��c:[!=��������;k�:F���=u0���"�y��d�M_ ��ʻ4�d!��A���"3E9���K�"�8i�GOH�������ƾY�kh��i���.��9��D���`�NM��h�juzzc�'e���L�,�D�pU㏱�~�~m��]$�g9~��#���M0�u��E㹍�S2�YYŢw�7��U�T����x�LVM��y�':��OŜ�<�G�]/w�V鬾����A`��e��F-��0i�_c���&��ą�f5���^�]p��S����z�լ��(0|� ��2S3C�Q�˚�R�L�AB�2�� �0g�@J�zqB�VhŚ����O�z����b{�wۏ�����E�Y%�_q.P���2Au%k�C�Ջ~���.�E�l�PW�e\�!~�!#U�����y����������?ka�~�n�"�ÅqSg<��w ��P���.�]���']�XאW��p^�,;�J&#�=��U��m���:���k�=~U���߈��7������<�s��(i�k��VC-�~�J܆���W��zy����x*&��!J]<�?�rY�W+�(w��a����4����p���#�;�\Ϻ`�[eq�����
�V����ҿ�t��le�_�B(ˌ�mT����#�_7���{ō���s�ʙnzt�?��й��{'t����p'z����,��ve%q�#�q�x���wv�/�oݼ���{�<h75�fQ�^���i��8�#�*�dhC�L<�>�L���>�q�.��^ 'F�`P�r�N<ʡ9���f�d ̶n��m^�����7�4�n�X���q{xǳ�S�/��G�
S��N钏�1^p�����ݯᕰ���\�)<�{�������W��� e�0�wAϫ��3��;�/��,��_�k��'�rz`����|��q��ɟz���'�������c�r���P�2�܊�t�mT������/'���Ey���K;���ɷ�b���O�3�U�{H��w��d�}�	��4��n�.���e���z�/��0�q�����K㨨)�I��*���󽶰4��y�A���[�(~w*}�ͪ��W헿�U����I��O�>��a[��A�66���/���u�jO�b� ϟ�
���v����@����L*�"�+�\ǐz���=��y�V�<����۵ʴ��+�v�'F��`�a�=�]k/��	�1����m0��Cd+B���vѹ^���g/���O�w=z��ƻ�zi�C��ho�������ÇϠ����!Q���r,mj���*�U�5z1|T�1J4Z��euVX����
��!w=�)?�����ۃ�O<+�p��<Tȳ�C�9V��k��?0Xܕ ~⤲�������5WK@NB���a�sJ�c�u��X��c��{��;{���1J�	�m��C���Խ5�\��s��t�}M��t�.�'���1>��	@�ں������p+�+j⢿�R�]⧟��F�!<!���7�̓z��:~E7hM��Z$^83��F�}�6Հ�6�l��,d�֒�ݥ�ON���T��4\���~�_�;��lW䬏C���ǻ�'�Vh'^�e:�Ґ-�`��'�c�eD^�PLf���+YV�.��57��~�Ȣ�w#+BV��c��4��PX�,�)B0�xPxb�F��M��]u�'��Rܻ�����������Ƈ&T4���E�������]� �xUP`���v�o'��e��`��?�r�U���Ӷ�O���YnA:�C��y��g�_`'W�*��Y��Ζb޺A�V�p�������0P�7?��3�c�q�������e�{�q\z>E��a�|]������� >��oo�%�Pf�����,y�����~���%W2��_�7���C�^˪��c�/�ƞ�0)�W�u~C�߄�~T����U�� �Ѣp�/Hw�e���'?;Jy��+���-}8w�
:�nK����G�U\rRV�xuw�Hz&n���l��@;�O�֭%Nf�P��	B"�H�6�ƛ��3���n���;�!
�̔QO��e{�3V\�]�,�o��^[�������<~T�(5�&#
!*���}��;G3�����2K�(����^�E�3w�VuA?�/局��7@�'>�4w�E9�_��Ʊ\��&2�*�v�o�n�^
u7	{3��sl����	�?
���S�~Q�]5�_�3| �(�H�^�7@��%8����įǫ�V��_�c3��{/����ߟ{Z��5�</𫴖��z=Ӯ$�tI8c5~�'�DNH+�Qp׎�e��H�B�灦�ᬽ��0lh;��Jq�Y�,'�Z�8���o�W�%�钦ʬršʼL���ʸ�K��w�cy��mB>1,�2Ї����o�]v;���m͊�~\��9�)�ݼq�}�����nݼ�|�Gy�;�ʄO?�������Oۧ�~��^퐟z
2Ɗ��'o�N���~{���6^iTyJ�
�J�I��:<tU����࿋��m�� 2��&Ot#'��6%�y
l�xn)���0��0�4�և큺7���<O>�n��b[{���n��K�:�%�u��t]Y�4�+9 ���hd��`�m�/�zھ~��: ��UK���
�@��3�vX����a�ȡ�w�p����I��~*��t�f[F�;.��vA�!�'N�*ݮ�LQ�<�N��2��u�_>�AnYSQ�ϔ�_���KV[�C5���0��r����y�u7�1�mz-u��WL9e��h�a�c�u��r a�,����p%��oV��S'��.'��k�:�]�8�1����C��I�	�,��ԇ4�"�,xi�DNpI3�d��IC���(@��[��mz8��_Z���P��-~��2OY߬rI7�1Lz�&��`��Q�Y����[��EF5��8-U�� ��QV����w���kW���4�b�N#K��Ε��"V�è.��Ȃ�6���T�8D����e�_>�{YƩ����kO�q�re����{���N������tTm;��=L�������_�Ͽ�����eQg��" |q�.�GŻ���Q�7�~*��e�4&���Sg%k0�|'+F��FV�@>1^dT��[���g������"`��kC�YH���08�������i.�Q��m��Ǖ�����+��p%��w���܉ťc�0\<�C�~>�{՝��+L���P�>��wv��Ex�{x�']ś�`A�a������o��8���	~�ȕ:�\����ׄ[��őQ%�ܑ<�'���j��{�T�(.�
O�Y�
/�N�@�w�o�5�ъT��|�/��9���3(�V Zg�=��=ۡ�81�)���rDAkt�����B����+T�6�z����}�=�˃;�S}s�z�w�n�{�v�z�
CM�lm����/>�?y���*�Q4�a���X�7aP�����pH��� Π��2�(���g�Ҩ�B9(��∃�.�������y�������86z�,�K~�\�_?�E�&�!ݨܡ�Q���ᩛa�`(��%] >� ��Pw�P�N�*�ұhyq7O�6~ѷB7.
��É��������i��_iG�Է�-Џ��Ƈ�����W�Ye�\����
~����!5���hjˑOI��:���dU^�w���U@��<��{�I�P�n�<��b[�_�f�m"���e��<z>�7��`d�s�e�㩃i���E�j�*�"�*���}�N\�?�B��>ϳ�<�C/���o��}�c��Q����Q�;���``��O�o~�yV��Bxyڏ�N#;&��B5����^F����������n��xn����Csu�w�]��*�,d�S��  }�6��H�=�Vc�լ��Wygk{g;+]~˕5���=�X��ܵ��OFt#o?�瑇�����U��kW�#�U��Y_=|���c8"Y��2���z:Ѯw��w]�B|1A�U,��hx
��-���!-IA��{C��Z����my�~p�r\qq�)��$�7�-�Yī�~p�=\�/�V抏�K[W�40<�]y���o����(�wls{�+Y"�QF��%^)P���w�,�G��GM�bB�p�qa}�C��] n���i4� ����3q�
�|d��&�6yĐ�,��?i`�5�{QÇ��.1`�o��j9��V�\���د�mW�n�3~V���5�(M�K~,�1^#�:�s.��L#�6�*��i^V�1�B&}l+�P;-�	_��+Yn�s�Z�ze!�}�#���:U �H����ٺ�5�|NI�ό��� ��UR�CX�Ȣ��\/8B���˷�{J�[���}�-��М,s��gL�<y�>�����������j_~�={6��`|��of6I �.I�u��(���!���튌J9edM�]�,��U��<*V��<Y֊�C9�f���l���	�7t��ϝ�I���d�5�Ѝ��~)9~>����i�M<�zY������W�	�+&L������rW�8����7����"��+gw{�v,$�ѿ���[��ׁ��Ɋ�w=�!H^Ic{z�=@�7��> �7m�����n��{p���#���ɃW�
v��w����߅qGn0���1�ː�LK�Qe%�(��T��q^Ja�[�������C��_|*�X���
uߑȬ�
��I�ap�'�2g9�-d{�q|w�`�Y`����jd��������3�W�,�[�o7�
n���͏?m�~�E���/�IYGp� �2�A��y7@�&xf�Ϫ�u@Q�hȠ�2XAd�B�FAT%�Jn,(}��G�cǔS
/����x�����q�6◟Je.H�QX�JBV���8��Z���U��)o(;�*_�J�F�CX�Yˢ�=?�#�p��A�u(EY%�L���@��E�ɣ�'��nƏq�<.�U����-�H�!��+~#@hu��r`ަM����T�����*�^|%�<@z��#_V�eԐ��	3��Kꐲ��h���6�-��<E��K!�5��7+�i߁W�r8�Ⱥ�;�-_��]A�ū?��/�pk8Y�E��[����x�_�q�FZ��]�tT�T��(e�/�߾y�}�ч�?�^���![0�!uw����O��ۿm���g�%k(çmfvd�,�R%�3�����
�m%�*��*���s�#\-�Y~��G���RWkiU �l�4��y���۾��!�42�p#?կ4�\�:al��)g�c�/Ç���Sg��uYX\��\�!+�A��!�d��y�߭��ny�qa_�#���
�J���+���^��mg�*� ������E�y �D��nd�(��k"���mz�I_|�ĸ.�b]q��B�K���O˸zC�|���|�9�i����g��S��~��.�e���V]�ϲL㮱'�q���A0~�s�5]�K�֮捶Ʃw]\��A;ܦ��Y)��YX��o9����(S��F��|�ye���\}Lz�,��9�t�-��?�[��v���á����)<3�3а��r4̲:���Up4��G�?Wm}�V�NҞ^)����Z>���,�������oyN_:!O��O2��-ٛq�==q���TBCɗ+=e����PD �"�����E��G5�q�ۃ��ڃ��촳6T>�G~�j�}����g?�e���)֯1��α�.m���ʾg��+1�ff���r:���B�"2hp;x���z����0�0�v}ޓwN۞K�'�d9# D|`z�n=i,�))�l���6I��0�q�oCat���v'k�_��.7���&�4����&	��Ly$l�cZ�
�q�sq���~�<~
W�kx.����Υ_)��U?܀����N� �d\�<*�� ��-�o𫛼0�
��k��9��b�s,`��G����̊~���n�xW��x"���$M�����CY�l����E����W�ɆX>�8:p���q����3�_��j���9~�+rGc��,�4!�|��Y*�#s�	u�^�_t7�39q��򿳁n=1�����Ӊ�Y�o�l����J֍�"��V��o>m?���2����v�:?<g�/���=
�����N
v�V
M�K�Xo�U�R�c���`B�˙\pH�K���T&u���l�wӊ�F�yY,�?����qp�K>q�3�@W`G8�O)�*#<�?���!�a*�t�@X��C���T��I�O��p�B����˲̻�bl�t	�%�T*EE� R�tSO�φ�Yz��P�A��k��|(�r_��07^����5wT� -��`��#��k4�;��JQ=~�3��/���^>�<��XA�DW��v	N���E��]�(a��|�E�WҐOڝK^ ��{��o�%�����w������Q��3~R�O0��a�:���G��J�����o}о��o�w߽Ѱ�"��y���~��_������W_>Ɏ����D��o��{p.)�n_���q����.��t����Q�Oe'�aVӕ�Cr5@�?#%3c�+y�]�L9��r5rܱd�Z1Y�_,9�P�dRn���l���)Ʀ�%�����T��R�FX�T�K�G�M=�>�C!F���J�RF��o��|j����ab�
e4��0�DI�>�5(��b*�i�h�3e�ꓭ����.�i�T��W!/C�~��`@�c�P��BD��Șa��+}��S!���ķ<��	"�������7�D��`��j�ᶉ��A?R78�zd�g(G��)b�;wSe<��4����<��. �<R2xR�:ɸ�ƴ����ʗ��R�j�����W��4�w]1�R����{�W��J�;�y�H���73�Qg��Uh�B����]0�b`ݺy��,ϵ٩3h��O������D/�WB@��1i��Q�XC���s)nw{�my���N��T�q���@`�h�Z�n�}������}������?�i�����j��}@�ö���m��t��勡�f9�a���ȗ��j��y6��d'���
.`���'#��z�=b4���gv�ߢ�`\���B3'��+ �_��!�x>���ciF��ag<����8���ÿ�_� ��?�_�/�{*����4��µ������ mHO|�}���bL���������i��:��.�@���nٯ�@���"��߼���CM�����Kj$�o�_���`*И)�w��|:�C�����6a5�E8�n�g� ��qR��סfX����)[����c'W�ұp*AY3r�IX����<5щ��L)���2���	&���V{��)�ã������Eɟj��2��/�W��A����V0�!��^������ώ^��<I�g�"W��Q��K�瑿nú���y��cy&�P���@�$��
�����E��_���g�P��l+�����RO�X!O�j��S*G����4`����[���(���m���ӛWI�� �7�B˶�b��A��_�����m�1vB�p'q�c�)w�*�O9;��;`��Hu(0��eK���-��?zp�XG<�+^��y��!�
҉m7������v#$�l��*s�#�JW�b�Oެg���V�8��{_�e�8��3iN�QJ=�9U�_N�b�xr`d)��I��(�,�[��������mw�@�Q࡭x׬����{�i� ������B�ʊ��A|���0>�\:S6)��gG<��Qj�[ .nR�[�u��枣�a�	y����E��������=������}�>�*k�0p� ˱��e�c�;�fف�!eNl)����U+ܾ�S�'���~��rRI��LyD<��4�V@V�i;����򳽤w���-�z�>n_3��b��QV)e�i�A�k���H*�U~�f�:��g�K\�e�m�EM�`t�o���y�L�o�kHfB�62]݃_��ɸ2V�刟�%�����ʘ+dY��iX����4�����mF��m����iqL��h|�"�����9)�8	i+�$�}۶2Mm���q��7��6��¶�q(]�3�{=gLI]�@��da�w������
T��0i����`���#�ȯ�Kq���wU.��Yϰ_UpP(��A�����x�w��n�[,�Y���{;��)�ӯ~������c���ݾ~�4��x\t-i�>	��y�݆�Q2C�F��A
�k�����0����Hdp���\}#G��@Q"���tw n5v~�uóa����|�=�S�r�uO8=����@�����C���=y��(���,+����:�J���Ɵ�ŏ[������~c��+���p�#~ԯ?C���!q�6l�����#� ����_���,���h�:i�D!��U���';�eɣ�V��hb�G�o��p�C/�S���T�QH^8����xϝ��F�v �I�a��a�f�����W�g:*���D�H^*$�6C�TF�[�K᪼�*���(��I��vP8˻\~fo���Tx�U4'��wU�mБ;�=#��r�O��EV	N�u�mׅ�̬w��� �<����Peih���)o)�|W�2@�v��(�#�{�C��o��`�8�k۷+�~���@ߛ����tG�#M�)��G>�f��2x�|h�N?�3��I�#�R��wx��j��^XAȁ9�!�������s�CT�R܀𷼯�2 �>�{��������wC���ʫ�g�٧]?��ת\�~�o���	��t7�x��Fd1��w�ű�E��6��!?�W�H=č2�.ı�ܺWw�xHÿ���M�W�$u�H����x =��P�N��YC�{�t���i]u1�ф�p��>(|V�ڙџq�&*���=^\cj7����Ϥ���~�U��}�����r(�ȓ�rj۠@��%�`��FV�m�����㝏�N!���.�.�\y緔��jkWFU¤�z���_����(�$��6�Ru�Ih@\g��H�F�J�h%I�J�j�?�)n�Rxx�ޞn��0�|�k{3�ª�+3�E�`��G:��Jo//�/����]Y��Y����Fc�g�O�_e�-c�о*������v"�+=� �c�X��O�˪�f%��J�+��I��r��
��<k]��u�t�����o=,�r����oVץ�-��	��#�+�랺�e��x�Ox��M1�e��s$�3j���X��}�2���zeR�8j��Dg��t^�g������(��>ۅ��xNyC��D�N(#+�Q���i��d�bp	>��|*b�)��ʒ~�i��'���J_����������<�W����8���^b�*I�^�ђ*��� ��А6�BR$D�I_�-�g����A̗�]�����>�"'
*�jﶧ�x���u�C�i�`����	Yf:Wfe��ް4N^`������"|�
�gx�H�"2�<�a�� v{�(ށX�/��Q���]<_�>�<��]�_�=n`yVa7I�!����$nq�9q������9~�`�o�K�y�U�Hx=�7�P^��6^=��}���p{�C��ۡ�/�^�o��¸; *i���q��5J�L����q��n���	�\e*<�s/|�e�0^�$�5�Eac����Q�5��u������2�+�ߊsQ�G]Q;C�L]�P���v?C+�Y?_7r-�xT�Ό?�j������@����^ځ�2έ#n�3�
�_���uU~?�t�^(��*��B���/��� ���Dd~�E1�n���o���t=��G�,���\��A<�K^@�w%5�s�p ���1|��x6����X���FH����uL���մ����R����i���3weF=�q�?x��U_W.�6��a�J�-��lx�Ӈ�W^�/H|��0����Xw��yh�B���q�(Р�m��_��t(�����������P~/x(�<ݘ��Exg<.�q�|Q\C�4/���~2�7A� �ne<���3�f�U�ݽ_�6�̀��^�q('�&��9E����ƨ]4�t�������]�B�K��?{�<Eج�;naM�/�"�T?2Y� ����U�Uy�.��)ĐRUw��ĝSɀ�Kb�p�1f\0�=����3��Eee\]�AzYG�Jd��<��σ}Fz�?�F>�E�����+�K�K��ի�����T��e�U��D�����(yW��mUvb�H
���V-�^#A�{��H`v ���$t%
�1Q���m�0~�������b1��*׭�4�@�1�G��Jj|����Ęv��G����,hbz�.+d�iP�t�M��2�ġ�UV7�>�w��F��S�[F��i,�����2���.k,Q���8�����э�B�Ѝ���WtAq^3��7�)n�gT�^�N ��!��lהC@�0Jk��o�R���]P�7��2^�t�؍���W�:X��i�ϴD7�42��S<�g��~�G�=6���kpz�s�(s�ҧG��"NU8�2?��*���C��r�Z[�~�ݸy�]�v5�VN���2����]mdFļG[x�<٤��<�&�A�X��/�{�8ذ�9R��;VH-"P$�̦��a=��^���� ���2Q��EX���~�<����zť�Q��*�夬<w �C�
��zU�TH�8�c<م�
_�� #�a���A0�����=.=m���Q���o�L�m��p�����5^���ʤDi��q�z�g�P��'�<��8�00�Nr�e��G�[q��C`࿦ �>@o���ِ!��+�S6�զ)�3�#���V��|�t��-̿�����X���W��c oC��]ś(:u���x2�)�ܦ���?4�uw�:F��f_�}� �<�����Lz/�Q��;3N�$�lPb�3�b��Eq�����u��E�q?�%�}I��Q�K}㐦�2�
P-��*+���Q�4��*�B@}ˈ��ď����ţ�<������;��2��_�DT91�'q%�t�=i�Ώ�˷dH$�E�ŏ�����Cq�%�F�&�0��Jy���^�>@x0|H�Ľh�қ0�M��s�L��8\� t1�<n�w)�ک�VmCS>�m/-*��'M�w�Lc��z���5!q����Ǡ%M_5Ը��SVOH_q*^K_�^p��UWjT�zY�NC'�Y��.�b�Q~�x�k��ݱQKy���=<C��L��7ş�	�d蠡�q����ж�OIS�1d�6��߇r��ߣt�|S���!��\J�� m�	��!�}~N���٩����*����&�&i?���ET�]��͏�:�$T�,#�&:l�n��,�҇��h~���1��������4���Q_��������lW�x����R���=� ��������5�T�A����5�Hk�glP�#�K<b\�ۡ�ƨ1Ь�@\��s�H�ܶ�Jr)���n��6��?���# ^�U�l�L������"����Yp��R�锃�=��`}���c,��x�U�`�7H,◡P�b�F�1����PN�W���û�5:�{����T�keZc��g9���9p,��[�@�"�[[w��}�~b\�L&t����>��rBۨ/����kJoi,ӗ D�Q���4��>�wE�vH=��1�Q��Wٖc|Ւ������~�W�̈́��i� ��C����������~��ѓ���#�ȋ��t֎N����PVve��d���MA|���A�1���Hr@��:+�=�����J�}�n{�w�;�ծߺ��Bt H���c�m��{����t��ӣ�{��&1�.�P�)�&�����|e�]Y��VW��+W���)�����D2�1xP�v�� w'�����m�v��;�$'�B�y�eV@�L\
��mَmd: X7�#Xy�˪��̳���4�� T��8��
�Э��d�L!)���ٗD��y)�a����h�'��;-F��#l�nP�0�����:v���Τ�7����� q�o��T��C�'�2�)�I*2~�Kc$�}�y;�'EB�N��ɒ,�����y\�:�$�2 '��� �նUN�H[q�uȻE2�S揿n���[�¼�g�j�/���<�'�'@�.< �p���9 -�S)H�Q��[����+��C��i�p�\��~��1��w�Y��œ���� �{	�!�D�e��Q�p�o��D	�{����G��z��$]��-2�ͤ���(&�(&�';�s�0��f۵UO�Z�w[��=8��4��pg��+F�g�;[mo{��o���?mW�.��߽��z�v�s�f��*��N�Z�����x����zF>� "c2H�B�&4�%�����.C?g�'��ʢ��[��'
��2?��3f<dn�/����P{ګ4�M���+���r:m��S92�u)E����ͣҩ,Ap��3��RD]�n��������Q��;�+w� �A�<�.FiL��l?�N�1��W��-<;�X��Pn�^�
����D%��_�g��%��k�0@����}Α[ʟ׀��2��]�J��8�Ed�b��%k�r����� i(���>eW�QAR�H]�w�`��t$�fs�mqa� P8���N�����e%t��(�i��^e�E���6�K�x�����4Wnꚝ�ns�m~v�r���x��/y��Ƭ��>#�i�� �YѴ�{�I���7�
?P����G]/--��Y��&t�->�僸K[��[�oӤ9@�2Q�T2�ce:E�T�La��:�$}@am���(/A�/ˋ�ݷ�{��bd�@{Ǉャ������'���M�C��T)�{�����K���N;;���P ��?�;�f��@n]B�]B�O�.�����h�sڏ~fw�����`<�̤�1=0h�t�(��ϕ��vtL|�=���k~,8ߌ��|��P�2�>�,r{���B�y{�]�q�-�O��Z�maa��ܦg<r����\oݞ<}�]H~#�x{���w\&���[����������i��dڍ��.�'�=��iWy�ռ�=���\����~nz]�\���<�/#CgO�O��(�����We1�Cߓ�=9��ʻ��?�#�q�H�϶K������N|æ�unf�-b�Ϡ���3  ��IDAT�q_e�%��2h�B�����R9n�:�a}��m��hЩ+�'���9<N��k��y��P[QG����<wK+���;Y1EO��6�ƙy�.��'��x��	�n|��������-�ϕ��`7��Ҡ}�G�z�2���B�Gn����ē|53?�x>f������4���KK�q�Y�2��^ʗ�O��s����?/DH��r�]�ɪ��0ҁy�k�՜'+7����.F����[���H�yc�ݻs���um	??(��]���`m�0G�4PV��Sa���ݪ�3g+9����� @࿕�+Ynv5�pr�;�ę���v�ޝ��G������{�sP��0�LN��������_�Y����q��w>̑���N�bZ0�,�8jCY�<�?ò�|�B^�-���w��"MO_�yP�qM�s|+,�Hx]\���v��\��ϲ@��`�YN����cll?;!m���Y��,�
4��S����(
��&���ێ�@���@P�趣��K���7
�]��?4E���(�����ch�=�i��x��q]\>w?��7/��q� G]C<��<���]"7\�ak]�/�t�ڤFo��ē�1��s�����x�ܯݩ�^�s�u#�5�7�xiU/��l�xV^@�R���ތ���sA�#r� Y�7p�g��� �1��*�g�^�q��q�F�!��k>��gF�4?�Ю\q��J�I��h.�E3ڒV��V8���a�!��G���V����x���4y_b�H�2n<��R�̬"KM��"������@p�n������ZÊ�Ư��#pI�ƽ����Z�\��iK�D�(G�K�~!@�)��p&����Y%t�a��K�yQ_�� e ���8��0�@�O�~���3-!B!|��a�=��̆w�N%�� ����g/q(w ^u&6�@�f� ����δjX�0���Vwx\�v��Ӛ�,�h�KN�GET����
m��V��0b��X���ʞ0�"B\�2��#I@i�F}��t3u��[�\�PY�Y'��*��])1��㼻T�;m:�N��Mu�8 ?�D�, ����*pƯq��Ē��D���T��Oդ����@�B���Y� L�P�h|^A���z=Fh␏�2P~!Z �'u�p:ø9<��b�ܺu���ރ��o���Bi�Җ���,J.����L��2XYĸ1e��S���|[]]jׯ/��W���Ut-�U̝Du�j2�5h�s�K�K��>'p0z�Wf�Ln����u)�*;UfC��P�w\�R?����k�eg��%<%�U�K��.*�2a%�Tn���8�n����,�'��*�~�#c��q�Ƀ1��i2	CE�m���?|�����	����1��
Z?���v�X�Fr�$����pf��(�.��~��n����9����˖'m2�(OS���ƔA�� n���N��QF�-�QN@�>�]�����ʑ����ʁ�����}SU�����l�20J��������?o?�Ƴ>�U�+�m�7�6~ǣƝ�w��f�P�}O�[�+_M��3��P�8Z]���ϧ��;�&=�'��<Ǯ�U�N泸�Ԗ�V�� ���"��d�j"|2)�A��0�4'����a�\�3��p�M�ׯ�o�B�7z.
�p��y:/�u�T�ryy9�b)�L q�F��/c�޽s��M��G�m�����t<;��[~������o�տh��_�O��~�'���FȬ��d�� �T
�ǲx���b���G܉R��^�P�o����hܳ����H^��X�K��{/�ֽ'��F�H��y�2�+ �j�U!�P�:@�q�K��,���R�+N
)A�ي�Ui�nIq;Dm{8wv��̭Κ%���s�D�y�0ˌ���8(L�c̩p����M�A(�<G0F#�x6E5�-5�\���ý�ҍ�8C^���?_\����_�Yh�	�2�`�����npT@90����������=K=�$�
���27��;Fa֣��w����C6����s��e^�G	���0��l���G�8 )k,'�d
���$�&J�w��,,"��=� ��[��(;�U�f���E��k�V�y��Ix���ʼJ�e_*��R�ʫ �z8�T����+�~��41fHW�L1��M�!]藤+�Y�G�Q�\A?�#���ף�\��UA����>`x7��x4{X�sO�(7[U���:$�:8]'a
wN[S�@�+�x��6�c��%��Ih�����5IV�ݯ�ĕ��� �~(�r,v�5�D�+W��+�� ���G��֠*?G*q$�<�{h�K�n/�
� .�����<6CK��І΄[���脷��<RR��|����W�k�N��*j�;����2��v������b��NӠ:|�������p�J�R1�w���xE�:�8�gZeEt��.�(K��B�:�]45����-K���4���<��T�gQ�<�.��@���k�`�����ۜvF������:��t�Z��q⊟�PY��W�O��#�b;?����kW�ۇ>@��~������?l�������SS�s�c��.ϴW��u���T�2�][���ޝ����7��n�w޺��t�=�w��X]lKeSS����:a̢|��4���﮸ц��=ӓ$
���<��;'��K��mV*���})�N���Т-�E�3Q�i3'�mw{A�'e3�s�i&����wm5����9d�m�
��`!��Qf�6>��2�)���+\��O��y<M�����g��θA��-g���W��"�S�ކw8?��eW}�퇔I��4t Wc'/a>;��?��C���Ly
�1a�H?񊜥�.��6U�|��il�-橡�$@�|��g�A�7�>(o��gC�)��2?r>�W�C�h���t"�ch��ꎎ��+��e���E}�H�z��_s%���I�r���|�Xo��g�O��W�Uh$^�u�2�2@�)g���?��y�i~v��LAVe�c�^�l'�J� �	��܈l5B^�"��9����:�y�����~V�a5J��hx�O�Qp�̔���̥v��|{��n������o?h�n]G���ׯ���{!����~��ٟ������q�������x�2���Uȴ�u*O�)�V�7��89]�{�ɴ"�R��F��<*^�ѯ�j�����4�uq���W)��,��+H	/�G�d
Kh���
	:"���5��U�;C~��/�ǸV�
�
 G'.W�M�!*p$l�� ~ĩ�� �G���G���@�2��5�� ;�JiDk �z��6*�L�-s b1d�N����A�
�C�j㸌���� ���ϳ���ʻ�t{K;��^M:zLGN�����rTy�6���c�iӁ�^�Q��[����܍k^�E}�>��	7�e�{��`�8�@�+:}���P�[���1���2=�k�������}(�]P+'|&P�N�g_X&}��V&�22W��$2�M7H�u֡,�J��J��?u�jĉ, ��3d��(�n�c,�i���g{(ل�5�8Hdp�,�o��r�/>B����b�Lv�VE��B{q1Oh��N�wܦP\|�5ʵBg<τ�4�w+��T^}��2���4m0�}���@��L�hL2@f��AU�и� P�U����\��F�J7�s (�c(����-z�>�Og�ὸ���c��o�q�f�7����Δ�����z�$2�7CSH��ݍ�����j�����m�-�~�r����4�iLґ�x�A)�����Af�i[�I.mzBe�6ƨ(��<�C(�*����MS��u?��9�����bEE�=cm�.!�p��q{��{�`K��`p�P)El����������}?h�;F�����"�Q��k��ǚ���
�&��0�b=�r���N;E��@יk�}���>n�����/�ş������V��e���󶂑u}e��^�ow����.p��b{p{����z��������wn%��V�u��EvW�ܺ��sk�'��yt&?�<���J�
�
z�˥�2ձBw�ڟ�j��}_�]ey�$���R��0H�b{���񥁜v�Y�I�����,�m[)k��A�Эy�l�01=�{yډ�Y�TZ#�$�B����z���(�� � �\�/�d���{�0h�6�PVM�sngw��F����[e�@���2�}2�ֺ�8)�kB�~���I �/+����@�V1P��q&�tꅴ�y��r��k�Q֗�4Q�Kk�<�N;n���d)��K���/y 5T}��R�@�H�(�XZ��A���#��rK?�-��<ƗG�#�xKG��+���w��������1 yByPc�<H^~���Se� 'cl.��|Vڒ�2��)A6:W�60I�`PW�JPVXœ�
٪d�S�T$B��!�����L�?����M�"Y[Z�jw��i�������?j?�������q��ݷ۽۷6W[�ڲ,~#�ڕ,v��1���.��A���@]3���U�Ġ�d]�Wx�_�j$�V<~T�n��-:���WKHØO��p����%R�;w�ª���3E�!fB�_p�h�&����&ԧ�R&�B#ʽ�G�E�ޅ������f;َ�7�W�h�U;|6�!a��WH��Ml*���!VF[\Y˳+a��W��4�bf�+=�C�D�γF�q;ȷE����UO��&}@w�ϴ���6��?F������ߘ�6�e���%
z< U��x������Fm<@@��RA�Q�e����Qޥ'�<ﵢI>��":��o�&^���0��4�6���ob�2��U����ꊼ�Ц�g��kW�P�ꄣ2���;��g��
A��<;;{m������>��3�gݢ0�n�Bž_Je+�R��� ����n���h���@	��(y:(9���u0�p[G7�X�$�Deo^5�]����@&��J���/�}5k4������@ݍo~��`�Ui�c���э�
�b@�VH|��sfZ�٦u;ω�`9rf������e��U���tšVu+{YU��>�� ��%�!�?��0n��(�A@�W�kd�F�7�
����Z�x7�
u�4�)r/:W�8̓m��y(�~����|�{�r���V��|y��?0U��%�gNW�־B>H"�)�L|�Jk:?�@7���i_��m	_M���誼(Wr��+�j'Q��р���ދ.�t��!�Ц:*�Qc`Y.������|C�K9*]�}о�X�>m�m�7��}�:�R��-�h흽����β��t�4�i���꜆����^�u�E����q��	���4��ɶ@-�������Go���w����������^k7�εWg���s��������ݕ���k����=X�J�+���+�[�
���T����S��)F�9�tqg���Smee�]Yqk�ʤ�
���m�KҴg&�ԛW�J�ڷTHm�(���[�W��? �mઇ+����k�%�Vq�p�E��郂<7�!�(W���2J�B&mD�j��#g���5L��ޫ?� ��f[wq� PM��/�:��|'�#���ԁ����&3�!��i��
t[�����1G�Ɖ�� o�}���{���(�3�͈���v\"\�P߱"��_�o�1m�ŹƲr�8�C��٧�� ��Y�ƭ���y��X~�V��:�б>d�;��ڄ�����`_�֕�	����C����C�B5y�M�l
y����US�c=�h��_�AP[����3������È��v,��5N��K�ۿ�?�r{��=z��>~�^�m����cZ4�jp	�r�/��3 ���𤳩�Ұ&	3H�!+�{2D�$�LS�xvܖ��ڽ{�ۃ���X�2뗞a�2�3.Smyi�ݻ{�=x��v��Ͷ��k<� �zp_��x
@A�C� )�\���O�&1��Ɩ�shmck�m��P�A�˄�m|��/3�4�n���ī;�$�cW�����y$�б:�0�d�;�LL��)�J=#������҇.@�i5@}�*/_�ve�ʐξ ���7��7����N1�N�I�bt�.8>tU��_@N�:&��<�|�%����1W��ϗ����+��0�;WIG*��"���҉<����ݒg��b��t���Q�L�pۨ�� �Nd���^C.y(w\���W����������e�Viu��Bܽo���g�9L�P�o�a�C�`��!����p�:�U��[N�����QwT���=j�?p)<-;���L��
��WJ�l�AQp{��THDOH�(����L�����`�3��N��p���\��nܸ�����*t52<!��/?~Ҟ>}��g���Yf�{�ʋ���d���ٶ�@Օ�}Wܞ�TG҂/��]�~�)'�p�PC�Aa���I��<�����(t;�Ut<m�Z�s �w���G1��R�X����;J�^�$큟�t�t��z۾dx�]��6�t��֖�r�x��B�"
���*9*e�5�:���=*�����q�w2���O��RDj�� ��àH��kye�5�����K�!>�;]"�����O�H����m�{m������8�)���~&�]����[5~-��p5�`?26��2SM�����S�3�]'9b:iJ�$m��������6�@��
{̶�p�ñU>�,q�w�kW4��7��W�)8|rB��.����Lx��R���sǃ�K#3����Gf��ku�ʙ�[�=-���q'X"��c��0����{M�o^owo��p�_ԟ���ŋ���Ͽl_?z�^�mP׃�!��F嶲ZR�`�`T-�]B^y��,F�|�ze	��\YY����[���[\�nK��K�C�8��L��'����Ƈm{k���|�vw^��1x��([~���n�,,R.�W�+mC�J�	e��-,̵���lt��zYt@'�l���������񃺮����漢=�-�?�>i�Bw��K��L�z-�G�����yd�ۀm*oۧ��2g�����1���@>M����U��P�+K�kҹ�&��6e�G�Ss� 3����Sn�ݙ �;��$�<l���LuQy�t�Iy���
��ݝ衙|#�<�1)����U�26�����-q�#Ǔ�&;*ne��4����u�Ú�(+㇄�~O��xnP�c���?��9n�x5� {���LL�HY27�|��-��1`Y]��_ʌ� ]�~j�;���1�-�|������t�l���� n��Ǿ�7+3��yY'��Σ>�K|m�u|�.�4��t�F���%����e�[���~ _�wY�||���*�ɝ�v��5��}�8##�F֓��K�,02�D��N�'Ȁ�ʎ����Ȣ�Tr�w5 ���p���b-��)|�l�*���F֝��[��¬J�
��׎D��~���hW�^C�]	c8����5_O(�qN%�%F�C����΀#� cq�mn�m����#�0|�F���"�$���LDGɏ{)�@Fq��
�<���;c-����F��F��q�Q4���/�ع2K'�9S��jx�m;}PLkŭ��1�b@Z?gl5|4X5z4�4��1�0���]:�|���A5�u�K�j�8��3:dm7��:)*�*�/�ЭYd����satI�ڦf=l{�g'����uVŏ�����JMy蟎��0�D�<������~r����⪰�ϼ�Or���|F�"|�0��8[�<[�ʡ�W��^���8�q�����C���a�G�����7EVo����!W��鑡U����������I_���@����6w�Ei���J�<,:+�3Bsai�]�ve�*��B�p�S�}���=zҞ=�{���N�Ё�!��^PQJ��yp^��gKx��AdDd�"R�A�t^[��n>�6��ug�@�0d��29�Eg�,�A�8�R��42T�Ke ���r�c�90�0q�R	�^	$ˎ�L�,��;3}ĥ*���A?��?3��[VY�@�P	�Ǔ��Kx�v5�
����O���(�Ӿ�C�w�� r�� c��a�*r�d��S�1��L܀m��q �~%�*�Ȫ��V5w9E^��Ա䠆	r>}��(2�v���� ѐ����x\�F�)�I�m=�'���M9�PJ�mO�b@~��Xc�J��ƨ�V	q�W��<��<��x������.��A�.a(�6���7=�V&W8�h_�j_Ǹ(U�Q%�pr��\��l�������f�j2T�:&�o�;u��9O�=A8�vG��H��$��g�j�{����W���[�&�!�rE���g�ۧ�}޾��a[[[����W���4�y��%�XjW�ϹՌ�|O�C^©�^>���v6����H[�����@���#�b�i��x��9y�1�8c�����6�����s��������UM����3��6�.�^��ж�4<�bei���*i�~ڧ�]@�����.��}�ѩ�<���y�d��[0����ۈ�Sx��	'e��T2�m�f'�qr��~��|#o����_������K��q��q�R#K��<xg��NNB����G�Ƌ)e\yq���]��t�U��P�F���Dq�d�tUOU6z��<�	��}S������ɑ��Sh��Ĝ�Ǿ b�G�����=�����d���&)�ԗ��z5���A�Q����Ǿl��n���3��:dK����1�����/cΚ��t����@c�P?_�в�	�s��Yzd�	eX��xkdv�1�m�B2�9n)�B7��uޡTf�(�c���l>����>ȇ�~�ұ�F)�Q7�[X�|d�����&O�}�*6��~V�__Y����s"�N,Y�����
�*&ΜefցC�'Pĵilx�Lh�)M��"��X����ݿ�ܿ� ��� ���R1���y"Tb��נ��J		�¬�c@�/<��I���4
����5'1���.�󶏑yr�����_�pt@f�C~Cg���z��������2uhz�c\\C��=Й�Ԋ���4�o��=@�����'��p��FF�ͅ�3q>G�{���aUR5�4�#��Z�"M����:��ed�7e*��e�j֠�l�R���� )\ʝ%��+�j%��u �`\�1gS��eV(b�K��q��������h�J�x#�W�����(<V_Կ��2��V�ĳ<y�?t0L?�^��>'�(����^��vqU�����xT/��|�o ���"r��s�r�_,g�u��YaJ!��?�P�r3��Ҳ{�<X��b��Uۿ�.ΔϢH,�\�g |q��R`sk�=y�$3�*S�� b��~�@ڈީ5m�8���dE*鐥�D��W���]���B��T�Vu��M~4i-0}+��������?�����m�ব�`Eʱ\i� UuH1�'xQ����HY�ATH����^��C|��6F(pI�[~�����N�<8�f�7�+3�l��@Ի�%g�XC����#��-�)e���J�Ȑ`0�]�G㍀���x�M~�9��p�1
�N�r�������Oê���F��8���w��2A�F��L�wk`�k�dּ�Ld�0�?�x8F�X�w�;#OɡQ�����QO���������cª�:�����
�}E�T��r��D�IY1n���|G���	��6`,� .u�����$m^`���z�X�{�MB��9d�ؕ�{�o���}�����v}�J[^�ԲI���%��/~��Y��7�W�\�>4#�������{��u��?�����JR�ǄKh���g?���Ǔ/��qs��|{��.���v��d�p�Zeq�mmmf�I�e��W�kw�>hwn��X�F�K���5��Q��������A������b��A�I7H=�g���M�$��W_kd�@a�t#K��2�oJu���K�)��6���n'��<�w�جr�m��PYV��� y�s�Q�����H���Q��<������f� i�)�u��o���)m)����X��� ���ȃ��>T��Q�Ϥ��_�)�e�~*Ic���%/ٯ}'0�>������kߓ/DS?�|s�2�ׁ�SpO�^56@s���e	��@Qd&@5�����QV��B���$�_ŧ��7/��cI��1g��d\��1ѱGy�X&^14���m;��yJ;e�qS^�is�@�C�O�)S��ɁK������#���R��r���Z�j���ua�v#K��km��b���r*뛍,���T�]L<�[);RN�!�3�~� ִ���� Ⳉ�<$�Jρ߾B����k�Xw�}��y�����X��*)0m���L&
�):�9��b����\�  ��x��,��o-q�>�b���1i5�v�Q�����q�;��E���n�������1�m����R��I��p��ֆ�#���e� X���
��(��Z���}{ C]ɗ�m�1P�z���U���aE��8�VP��Ej`�UQR��'h\�������"#�ΥT�K�+��qEx��Y�Zөį�Xn'�v�
+Ғ/u�Z���w�k�H�m���i�s̋ �n�9�N���d�����O��"Ou�/�jϊM;fV��zx]:g��W�ÿ�0��t�O���+@����4���P�>��|.��o<r3M��T`��{��ǟq+d�G���W�|���)���/��B�ih��H�0?�������X�K���O"��I�A�\�Ү_�������g(_~�U{����"��c�
�X���� ��6e�O�.��h��
�H:���}=�ǐ�e9p8�Pc�ۤ-��t�Kx_��L3up�_�+�z��r[�J�����������d@�u7\������als�����'�E[�� �J�/}�� ��;!�?e L�E]ޘ��OAɨ�!%stT�ρޡ���%e��1'wq��t��Myy�3��g�>kA�i����H$�'V<~�I�ϝ/l7P���d;^�L��B_'H׍X/����������O��Q�D�W:��(���o�5n��Aisp�)c�,�芞��M���v++R����	�u�Ji�D�:	��W�\�p�º��(Ϛ� K��E�`9U�Aϰ� m��@W�UWX��ރ{��ￃ����^] иkȁ���'�������#����v����͜�^^Z�*�������~����377ޕ��țY�k�x���{]Y^�a��d~[ȃ����[�ٌ�ȳC��],��Q��WU��]��F��g�i7�;�O}>j�n�#��}9tp��X��vt*�[�U�Y���@Y�����H�g��z�ս����˵�`��= 䨓��u�U~��$�}��J�jb�ЎG�in��d�G��diV����D�lSE��h�dB�q��S�����x�D��WV8���S<!���(f{��$L����,_K>T���r�	�������pV�;'YD�0i`���oY��93�x�b4���ykwFe�1Z��՗�ku,�.�p3~в�X N�E�+Y@>��?ZO�T&ێ��|��m�hPE��.1z���J�e���,����?~���*'@{D'��a�6Gތ��/�,�s+,���2e�)#�,74�_�+$�.�!�r�������3�G��w����n����6��;��ͬd�q�1�<� !��h*�<���$�{Y'P�ƢBVֆ����V���^�w��߻�f!�8v��Ν�%ꬊʏ�)s�1�~K�l"o� ��Wɧ齙�	b��*7$R�g뜲��F��c�u�pq%+F�LV�&a�� 1��`���*O1��a�yy��j�6d")�#n�q�1N��DJf�3��QT(3���j�"3�s�����T4�Tn���U#c�)o�}+�,��=����!�P�ՠ:"/�J�[�8�G���U�Z��x�P����KAS��LZ���}��
�l3HgA�IʐY���sz��*
���Qkȧ���
���C|�URü�ߐb���\��{i|���s݇�
#����^�����A4ٕw��#E͐T���櫔��+i�5�s����5��#Z=�]?݉Uφw���yF�O����r�~����O�RV�s@%s����d�ھ �/��H���?h~���v��-��T���j_}��}���ɓ'mwg'ʰ�z�zq�/9��?�:�����6�u.�6�o��<+m噴�S��:گSH�9�GA����=�S�ǀO_��l��AV�m��}ξ)��7�_y�����_��o����r2������*H�u🠍�_���pט��(�8@����G>$_yF��D���,w�/���.<�2����xt�$��~��L��/e ��Z�7�Xv��=2��$)y.^�I}(/i(�1l�˥d����<HS
�tw��_��^�`��Hq�B����W���=������D �U|���eͳ��2ȃ�U�j�K}2 5F�� r\vr��t"w�F�@��L]d���ގ�V�B����A��|�#i�|���t�)hxif�� c�+�d���z���1��c�LC𸭭��_��7�����Wm���++����++�{�����������C��v�w����Yׯ����z���v���r��?w��+�Ȥk�O;ދ��턾D���L�W���%'�����u�=2rv&�W��n�����ow���u9�����`yO��l/�Ȼ8��լpYY���e��I��-T�G���ўB��O������r��'W���}�ns�T����逰��D�j<�V�Qv��ĝ�&������Ǩ��!���I{�+��79U����+}��E�W��Rח��w��<פA�S��'��?��3�c?M��Q�?����˕/�r�$9�GVj�������]�*"w�Ӆ\O��Y��1�� (,�H�������㬬����a���Ե��i�C����1r�1���,/�Gxԅ�&���xJ�2n��Q��{h*���X1�] ��1�CW�p[���H>���ץmv�>`�v�^c�#�.G%��t�Ed�;:hjss�J{���|�N�k�;��.�������흣��Y?�b�	f>uFAև�e�W	q���8�����S�$+rVJ�������U�6n��I�^Y^����K���X�~�ܙ9����tas \�P>��xw�S
�60�b�-.��g��o\�����ɴH�(� L"'1��0���Ξ{1ݓ)1�lx�B%,u�ì�W�$����;{bW��;�$6|r[�0�ĭ�cv�3���D���l�N7	}S�e(zH���2Gڑp1�pj;��0��`�sW���� ��s�����D�����6]oǇ��`��r?9�"�2ܣ���К���fݺ	21f:�Y��H3�`q��v���v4iU�=���P�Xy9p�By@}����0y���+�~��;�_�q���ߏ�$�^_��S�C��(��:��:���S��]�pq��*��m~O�Jq�h.s���M�ׯ^n~�y��C�@Ņ���>��B,��mMX	�j�\����D�:���'��.����tHY���N������s�7~V�r����q�뾩��ɻ���{yJ��6�"m �a��ig��y8��*V}��}�r�	��c���F�1
Z��4t&8J�F�uō�(;��w�y;@������}������?k/�>i'�#��\�w�K��w�S�H
l*.���'<����ʺ3�Y�.
���Жp�*2���`�ʥq��>�J���Τ���/��"����~�ɒl&NʊQ���ݙ���i|e`&W��8RN�)/;���7�(E�Mo�X��9mJJ�i��Ų��h0.�?!Ql�@�U���m=�n�h+)����Iޝ�������&-��se��*0�rB�X���qf����	?mS�%��EB��	�@^�&�K��v��&��]�1�	��&���jY71q@z�3V�n�5�jZ�L�t@�(G��9%�2���ϑʓ�� ����t�Ę~��~z}������a��,+%T �;;�!���2m��|�!t�B�C;�۲�]
���6>��G�w�$a���U�I��+٢_�3�CK�'��=	�J�>=T��Gx)��Gmk�,߳v,�dx��m//_�(n�S��~d|��7����1��$�v��J{��{��w9��D{�lm�/>������h/_<C��n�G�3�c�+Y��o����kmg�e{�������oR�y>r�6��>lw��k�</�η���ve�*p�]_���v�i�-���r�B�@����y�9)�ι��Jzj�,z��͑�����FO���v�3夓S6F��b����t�곴�����w�˱@�y@�lmﵗ/�����=tJx5}Y��`�'�������muD�	�S�R�G�TP#����g��6�mow���xZ�6a�{�No��'��+������=Y�rc�-a�������㘾�d�[���4��lm�c��*��M���d?������~����5���x�:�?mc#K�R�+2j�>��z'e�Kv ���)�A��N�r�r�{��VLpCW;B�;��-�Ii�i������`����T����7���ދ\T�?��B��_yFD���j�FϬ�F��}ж#N�R7#~OG�����x��������u�[����!��(�G���Y<p��p`�g���zM��6���n���
&�	8��y�߉����F/p�vnY�6��3E�L�k��t��<��޸�ܹ�n]�B3Ӗ�+�ۿ���s�=yY+Yk�d9��Q5�Ҽ4�ʼ3�S �� ��@�m$�����WihEH��0V%�R�L>%�`* �\�
�q�z�(�?������]�r���΀�(�����0_TS�z'���5;Ge���U!��3xN�����#��/���X�����rx ��^���a��+�↑�+w�:ϦOb�윹�g>����Md����<�}��1�5O������})�v��ȭ~�����Sʈ���w�J���� ���4��TrUvK��%�ڮ��� �"!��&�C�U�;d��a��5�	�ze�*i͓6��sEKR���u��?Ǐ��"NJ!�jkT�@P½R���]�9i@���>"d��>J�^Bŏ�(�O��-��Fg��/m*��j�ޔ��z&�W92+��0��_��NY1�盗~񽈖k<��tu�W��SK�Tl�j���=V���\���qh�oi`;+?4l�OO��̗���wY�K匲!���s�l��G:��,���|IWYt���v���v��md�t�Dz��i{��q{��y��ޡ��(��a`���P�Pge�u�Q>βe��2Df�ٗ,HXJ!~��ۙӒ�%oS�y#Q�yGxU��?�B��Q���c0� ���t�g�k�G~-C������W�%�*����z��˼/ʕ�KzT��׻�G����ZyƂ�����= İ�F�e#ws$1���5S/rB�H|R�>Tֹs��C��X����m����V��356̻Oƈq�"�e_Z:Ԫ����c����Zk$R>yQ��l�l��JK��7�l��BZ���O1`�9�t��ɿL?�*'5���l����A�z��1���{)�LxQdm�q��$�q�/K�&����=����K񘔫��qB�0}N��n����#]m7���r���\x��;o�ko?���{;�>��~�����o>k��k���ξ��6�j�[�<�b�is}�=y�E{���F���)�7o�h�z� s�\��,�U�zg&�E</,, ����C�|gT~Ӹ�0���Qd�fE���=͋o��]B�?m[[���ګ����~*�0������ƶN������g�[ ��й���d��*��������0<�JwGM�}+�^켪mm7'��d��;�Fs|�5,T�/]''�1�N�<m�8�k"��q��B|W��by��R�}c�ݹ��n�o^[Y�X��44&,����q#�6�w���vsu9��\�T�+n�D���҇Pm���O���zʺ}��95r�ts�P�IW����{����VW���zͶ�K�zi<�s�|�i��dg9�n]kwnS�������,Xxn��!bg��w�g���2��b���L��>���.��~W��-����.g{k�i[�Z�'��SA�.�([+���%�'�}ܩ��ǘ�>i�x^�˾,�^w?���D�Βn��̖ٴ12��!�_��_9c��S�cc,�f���U'0���0ˁXޕ��a� @⿣xi��!�{�iwϐ0��՘N��O�������^,O�𵽣�n���w�l��o~�~������q�9�#xRK)��a5	Cζ���62{�t"�8lGζ�4�U2�f�N�b8a$!P��3Oɋ� �i72�����ŏ�;w��J���@C9�Agui���V��f�G�K�{�gc�p�����S?\|����Q8�0/P�0a��{Wۻ����x~���������n�g����.�ב/^��<��Pp) �*���)�S�_p�9�(?b�0���˩I@�w��}�)�卌m@�ʘ���p����A�	&A`�1� ���������=�O�*3�t��H�<��x�E�*����?�Cc^�N�ė��\Oj���K�fhrg&�Ze�Q���Au��W���+���2J]'"ט�]�ȳyF�` � �t��n@�(ovv��\�I�0���O!߅Q��e��y{�NXݡN\�'@$8ú����K2D��Wв�B�:����[u���[~�`*e��q�uh��i��"ޕ�<�S<x��cI����&��.q}�R�κ�2,q
��x#Q'Ő.y���D-Ή	g��Q���z�l��,--��W�(!^��g�<]�
���3��r>�*�G��::���|���w������}����{9��˯�h�𓟴����~��Wk�m�Ke=uW�������O��c»m'y�z)��a�*��i3ג_��/T&q�pE)�^�7}�2TD/�����C~�c��y��!#�-\C�r���6���NWWHc���U��0�U8�qٟ�
.��FEZh�� L�c���yJM?�p�WYԽ�.�U%'r~�]P�+�W�'}������?�l*�-ct �?�P7j_҂0���>I �D݄�"̅�����ҝ�����#_��M������9���։[JMpJ�
�:Dzy�J��O;�S�`Q~T��H��d��n�u�)���e���*(O��ݬc���r���u%`�1���z�� �L��/�4V��eDW:�ob���.�K����l2�ɷw��As	�F���a9�pW���:B�G���\��Z9����jN��:��h^�@�n?�އ������������3���o��h�����k��?���~�����I[x���c���P�W�[����n�8�̓N�1D�a�����G�|��9p�my94���n�V�b(=4J�۫W�׿�E��O��}��ox~E��P�K�eKgA��|�'�Y��I�D9��'��ݶ�j+c���9������֦F
2�Ѹs���{�m�WSm�6X^Yls3���U�w�mcX=~���g�l��ͧ�%��B��s�s��@�e�>����t�V��<=�b�^�}��Tp�+O�{��tѳ�"��,G7NN�s�����X� �z�j��],�x�pw�a$�o�����Z���\Z���ܺ�j�1x5h�S��1�y������ï��W���1�w��\���s��z[���(���|Wn�����g��㇤[G�_h�Vo�[��}�|�8�W�w����������	_;F-��..b,��{�����ʮ��/_���=��~2/L/�?���$:�n����wy3�����,�Q����B�ԥl�>�ޟc�1³ˁL��Tn�(b>�W��#���}�����N
Զ��]�����<�����z�I&kh���vD�K2	^�ϻ��x�����]���gg'��l��K�W�%ON��	�&0��u��c����PN@l��7^��y�޺w�}�[�������w����|�����F�I�=�s"�{���-�XK6*�r@�o`��#�NbGp�(/�wv�׽��!Dt	Ud]�{���v�}����O�G��ܿ��9׎`d���6~�fC˙�w�y�ݽw�N=�U���-�Ţ�k�2�3��5;E�1P�q���"�����s��I�JC���/Oۗ���|��!_0�`���(+g��2�kFV����I/*zb���'�`d���0��1�p�)s�p&�x�
]�>��`nU�~� ��")�80�=+�S�2��d�����pf��q�e�"��>[m`�K��Ga��)�r4<*�D�)�/O͓W�,���I�ԋ�"-ӗbp�F�s��(hd��P�QE� .�M|�P�?J ��1�>
?�Ihc��Y���2��\�ns�'�$�r#뺛kfo����I�R��Uq����Md��e����>�h��s����~I�U"E� 4��5���H&ÿvUz�C��k�o�ׯ�n��m���e����8͘��z�2^n��m_�>��x�0N.À�j�_��к_��ꇨ]y=8�C�n=�B#���o�x\�3Z������O����28�_�쐾�>z���s�V���ؾ��o}��u/B���G(2����o�������|�]Bo����]EF��lr�q{����"���(Eg��o��gi�;*S���\(j����]�
-UʕWǙQ����g]i��$�h0�v'���2���}��I0}�0�y��`�/w�@���B����Њ�83�?���SoO��W�c�HC�n����}��g�L�����U�!<�xňJ]5n��4F��3���E<��|3��D�����T�7#�g������W�pA#�D����h䚸Ǜ�*.�<�F^J~�W�h��]:#~d�Dr\� ����b�S�x��iX1�����/�C4T�A�Π�y�"��Ye�����*� 3u@�A7����{n�Zێ�#�Z�s+�����G�g�Q�(����*�"�,��_K�4c��
s}'kn%��=�0��9��H�O kO���J�D�.������?�����uw�-�"ѥ���Y�����_������?˄pY���w�\ź��\�@F-���Ab����~V��y������}�ݶ��~s�OC8~y�HR��5����v��'�l��������?o/^>O��n��&-�s*���U�X�.c������~NV���{yp�����v{��J�6t�X\Xj׮^k7o��!e7n���y�sug�����P���k�?�U��O��=}��|��1�C��# m=����C�2>k�--]��}O�~qJ[xꤻo��:���$F�B{�>8ݽ�睊gh���~�{	�������?�������O�Ͼ�
��m�t_��5o���k����<mA�~���tY�|��}��g�������y�����[o���n����C�T��?�����z{������b�=�oWڝ�o��߾O���[i�X�d�[aw���ƴ�(��]�p5QC��{��Ή��`�s����|O���pW)7w���拶����#�0����>JS�_�;x��B�B�h��-u���.s,E?$���ㄆ���|]��W��.V��e��߶'�����D���Š"/��s�����nI�����d�O���S�]�t}�7ߨ�V髯�K�=xh$�O}�һ_�a�]��q���
h{�qB�h,z8ߎ��ol�͵W�����Wۃ�7����ut��K_�ӗ{��_=Zo��'�j�������i q�lYub��ΥX������a0�{jO0��m0�O4�4���X��?�ײ�e��0
��۫�~�����o޾���!�˗/��~�֩�F�����>����[��R)'������+&_Rm���Ѱ�3�Ч�e rb�U��Ȃo۳g�1���Z#k3+Y��1Ď4��F�и���4������-���?g��(�m}�kF�a��4H�y�n�dj(�˙�ʬ8�P`MMNWz˷N]R���Vg�]�ʉ}�g�Q����x�`��(�T�TRTO��SHp��r%���,Ѫ�b�8�7��oe�CK��.���C�*����T�|�*�5s ��j���8T�T��T�qi�m$��@	�̮�g5�ecv%����7.1�L:�39K�
�%���DIh��W�R����G�hx�Ս,�1.�%&����Zm���+��� -�$��Ȫgi@�
��Y�w��������!���z%�"���s��Gy.q��$���7v�<+>Ѭ����r��� �d�A;��f������+��D{����:W���Ŷ�&�
���V{��������Gs�2���1Ԝ1�F����;���O�����(�c,k���׿j��w?i���?i�~�Pw��Y*�ֹ !a�ϙs%�<;������I��g�\�J"�;(9�p�ď��*mk�4=A��G\�s��E��.�e�QV�� ;C\[c�e�4.�Բ/�$�ߛ)��O�G=]y�OG�V��ϣ;�p/۷�<wF�>j:��x�Sbq]�E�w���w������|[�(w�C��>�s��@�R�����E�����
�WX�މ$d�3�a} ������W�����>�I6� ?e�:�ZMZQ/iAX� ��`���G��S��n'�������.y�α�$��ip-��k��I+���|q\��<�!d�������񎣴�]wa���j���;,�jÉ'9�wp���4
�+*t�~F���n/���E9���Di��KK+(�K�J*o����%����WQM��n�0�2
����%k�#�A��-�O�z��i�����``�������p�-�3B����FF�/~񫶉���*�
~>x��vuy��A��������2?H�rM%�%�N��[����]�q��,�'
m��^ڷ�^��=��W����߶_���Q>�#�B�o���.��Yhhi�^�(��^l��W;����9I;N�|�g%k}m��܆��퉷0��adݺy�͓�"y]��C귪�5�;b�Q��cd����������'�����a��C�^�4�vw�0&��hs��r{ە���y��Pgmw���b{��Co����n�����w�ի��e~3n_��Vi�{`˄i`9Gs��4_�>;>k_?����=O��zm����N��-ͪ�P�ۧj$}��Ü���h�jd=x�v�y�
���6G|5�CXvcs�=z�t_�k/h��hd=h�n_W�1i���eY�-u�m�j7���mK���Ճ���X�j�ƃ���o�m�d�� ��W;��K�f��C��o����:�rӇݪZ;�G\ Ah��;�Q���w����xG�k�{J�+o�.��o��ڂ��9��Q�WV��CY�l�ߕ:�7L<4��1X��x��l��|�zm`[c94�n�v˹�,sL���J{��媔[\�h�	��Ex:k���\��9>hd敁���Y+��53�3��f&�����������ͭ������գ������j΢��\5h�d�}R)O	�|g�ܦ��*����D�IQ�����*��!�Bbc���g��[7ڇｓ��Qb~򓟴���7�k:��b/'�p��C�G�?��O��˨
2�vc�X�-e(L�0{�j�"�0��t ��c��}�YJ���E)MRj^51����U�3x�WOH
<�Ѕ!<��(�i�!~�wض��o��޺m1�U�Qꮺ�<�#�������tV�1�|Y����3E\S*�մ�^F�]�虚�|�p�U�qa�9�fip�֠c�7�;���hkD�335�/� "t�RR	��V��[/��/�a:��❲�6�@o�F?����8-�v�%^��ܒ��J�*���w���-��,�f�u�Ío�J�=JӀ�k��x�$�>�b�/nuY|��_��Xu���+���C�Q>w?A�����G��:�rFa��/���:^����g��V�1@�9f��3H2_8���Ŷ�6�W�X����E�8K]���#��ð���#����{��m�'xݽ{9t�-38Lc�� �]�W�󽋵�н=�gh�d�΃�U^: 8C��y�|�h���\$�ٲa�Ⱦz���d���\i8�XNf�8U`���/�uĻ�4��߬q�5���b�18H�dI&1�(��*���A���a�$q�P9jj��K�"]���N��q@�eJ��z7�ܙ�&1�&Q� #�RV9\@uƋ)�ʝz�w�J�=��2�����=��*���Ϟ��;�S��sB��2�>��׻��Sdi@eϲU���� -� ;�z��
9�,��-�����ĵ�)'����MA녆N
�E_��,����RB�	�9V�%�����L��}4e��?��Ƽ5f|a��%��h_\\��=(҃��:}B%��ݪ�6*�bģd����i��/-��!ur}����h�>u����)�N��W>S���a�����;��o��O�.�	�.�+��
F�����;o��D�8I~_u�O~�i�����,�O�X����Z��N{���o㥢��^u#g��!V1f�h.C�� �}l 9�$?y�=��a{��N�(yw��K��N+n�x$�
���J�	2m���c�m!�WM1�)�C�[%We܉r���G^ZX��i�ˮ�ۥ�I�v.Wz�5Bf1�r�>��]7s����h@�n���1����p�M���}� >;9���F_|�~���i�۷?z��M��N��kW7V��^�񵲌މ�8#/A�,�VN���$OK�u�zމ{�-�����߇���a-P_y��n	�֙�߹}�=�w�ݿw�ݾu��)Wh[)�D����zOIC��j��i��.YzW�4S�[�g�Q����֣��a9�����N]��Q���fi��/e���"<�@�\����Iׯ���n�{�&��j�ﺧ�6�&4�	���U�*1�(oc�ާ�܁��{��	��ܺ���]�~�4sY]5��E����*������3NI/�=��j���HcN���y�nÕ�+9���w��ɟ�b����;�(�F�U�o����uL��)34��zs��u〣[`oQ����z��ѵ���)����bV5�=��[�R�����HN -���_0���_nl����X�X���H���R�ڙ��Qt��k�,��_����BJ�F��3L!������s����86�G}ؾ����8?{����7��4*4Z�n�qV8��
�a��ܻ=����=\R�^U2�{�P�d��>�������ɂ�X��F��W�u&R�C���_�J��N����
�"�x�1���܃)�р���`桷w/�*DUa�[FDuª�4.DW,)*�+? �Q%���;W�_�`�&�/�������
C�V�H$3zD�4
�̌_}���X
[?N84����D J�TE|ů�;A��{*v*�*lj����.T.F�P{b�]����@�҉� �D����>���H�e�)P�<����3��1�
�z�\�a���P���k�Y(>�^��s�өH��T��wEC��_����5��M�ףp]����<$�y^+��������x=:]F�n���JB)��ʣqo;5W]�H8Q1@�%��W�n�,���
��mhd��ao�~��^)P�ߗg|_#�e�U���;1��0P��)8����E`���l�qu>�4 m)�=��"�b��#�s��U4�i.�B����2|Th4h�M�D�j��N�d�g����3ۨ���M��k�LYNu��?�\��V�9]k*%g�U�T�j7�L��mh{IW�YN�
]4��K�[�a�Eۮi��7y����u��"�TN��<�{�N��b��wܗ.`�`i�` i]�`L@In�3<�@��G���5�3䛧�M0p3��O�8:�^j������r��!���xZ�y �'�(��P1/c��b�i����	�M4i#_��=����g�Ѩ���\��U�
8���$�G�h/�Sމʏ+�f\��������m*��+���|�o�q�O��"a�%qF��1@y��Ã�F1�ڜ+L�nY#dPy�/X?W&�B�$�����z����X�y'c8x:y�V����ƂJ��,�:�Sm1�?Puw%XC�J��fz�Y�%d�"�p��!u�����S�t�c��(�|qu���o�ə���_����mw� �Ⱦ�jˤ)4R&�D���D��?Wٔ)���P&?$68۔ѩ�,}H��W����g�ۋ�O�2a\��u'b���R6��O��mW6������;T~[*�Aw���C�3J;����
��=���+es�mCH#kEx	%ܼ�9��=z��}��a��������'�OP��o~4����������4FpV6�My�?�u�WP�?x����}��}�+�u��u�C��� E�)<t�	y'9$�݉�Unppk�"u���E�:�_�Nœ�3�S�$�ʡqv��h��U���Ne�LR����[/P�}G�:��5$��SN���M�^#��fJ7ˡ�MU��rt@'s�n����\u��2ل�����JeĨǑ�}�NG{{<�:`9�x~&�����bj��6FP9�H�����ZH�x���H9n�w�^��Чy'���� fh��9�>��/[����j�U�+ԅ�Z�Lk��]��Y�f{ ^O�g�&�|�����4K�l�<HFC�+Q��˹��y���]5��������2����c�DN2N`��0n�A�ҝ�������^3gC��̥P(���@�����5#*�Ȥ����w�i��裼�����t�X�X�2�BԴ*9O�=��>
<�mo#��$9���h$9{�d������z�:���H�Q�� �������U�(��W�}d��[�0���}�S�������=�cf����,s��K�����*��[����"xz��_៽�+0+����v�Ɲ��8(�"D�]�0;�3
�`��kyi�N�G�a�E�nے�� t;��ˬ�Θ2�qG�F��GO��/����#f�0'b�%�ih��Q�>����ݴ�q��[�=�ӭb4�F���*�]q��b(�|!u5"κ�s��r�. ��?I������2v�R�U�8x��E~��!���)����$�.�~���c<������>�C�r�]����w��Ah2J+?���"!�R�Q����W�� ���� ���,���(�B��2�+�88f��lf�+ӡb�ÿ����8���U�v�ȁ������r����g��n��+O�u��s�_��^Ż��U�l��3�'�:\v[R&@��]a�I�T_��ۖ?n\��'-TB�p���u�Jc���q�JHe��;U��p�'��<�c�QRC�m[ӗO	SaNx�����0}���~��3���m�����O�Q[�9nW�����v��t�wc�ݿ��޺��޺�Zh�o̵���ڽ�(�7�r�]�i��N��W.��gmyE\�=f�=B�R�40un��{Ļ��|y��#�|��p��e���A�Y肛����	�4�!��er�DW���	MOh��q����o
i��z[m�!��َ%�3�`����Ћک�@�;�a٠�GK���R��*������$J����-�*��c����t�ʱ��p�
��ODY��cF����[�"B�����sp���3�3�rYl�X�FdaNr�q~'jv]GF�oX�+-�*k�q�b[8Tt�Y=``��Z{��q%�X���2�讉aqd`&yS�����+�|?���EN�������F�Ky�l���ہ�u��>n'�"C�+���;i�t���y7�|"k"�
���;9�ε��lgۓ�5���%4��	�d�\R��}�Y�]%uӉxZc]��_�4=��:rJ~ ��;��
@��l珲����g>����l��
�W��=|7NCPz�dEhC�����h'M��;刋|�����2��Ut�Ep7Q�3<��[_q<� �]��lS��c���·	օ$��̓�\@8#�i�s{�c��PA9|������E��Ɍ��g"��}�67v���v��B��6^V�If��L}~hY{���X�=���W�������e[{�ֶ<(d�c�KT)��Cx>:������u�v7)s��v���������{���[���4�o���ݶ���^��jkO_��g/���+��E���-�j�d�,�@4�CT�ݭֶ7��{��a�w���1F��E�w�W�k���������t��a%�ź+Y
gPG:y2L���8K�-;d�U��ΐ�vQjm+�X*�ƙ#�z8s�����@/s:��2��}�}��0��¨9I�r���t�zt�vw|��V�)/e:{YL�쑕�<�<"�"�	��F�q��:i�����}�ұ������U�u8:P�u�2�l�x�*����+[0�p���^�{����i8��5�f���6�g�^iL �x��
�@����s��5tF_�����*���aY��V村t�[C��/G(�T�j��n��К'^�ώf5t���5��˾ջ����Y2�3�E>"}��QM ����w�a�} �Wv �S���9H�;�ЪN���|�d�䚘����v<��B���!1����Rq%�mZi��#5�A�~u��1��Y�rw\�,ic݇��5����Ah�|캠M�j�a��R�,�_)_�og�+�;��~9J�z�)C�����,��`�+̻�P�t�G2ku����J�x���-�P�$9�[�����r}O�mH�ی�����׮+YҊ�edsc������h�$�22ʕ2Y#��(Y�c\1z#�8�g)���H*�Ut��W&�*���A�ǖ��"zp�Y�ZuO'�n@R>?�i,��f�-X�g�D�(
CUR�J��'���Ze-�+�i���t���yj�8�޺�
����F��6<�b�N�Ӓ�x�OK�aP`�hp�@ �Sih�~ޅƅ�Id�T[Y�ɶ ���d��Vn���"ϩ�6{Y��%����s�GX R�Ϝn��{�ζ:��}��e�)�|�������`�zb����#᪝�B���0[	c0�?sX�ҭ�"���9�������S������ҧʧ��� yɓ�����i�Ħ����$q`�3,s���AL`�dK<Y9�{���}M��n�rwZeyέfN�N���*���c>�/@D�ˋ�(��\H�W_.V}�K?���Pqf�#�5�P��A�@(�NZI3h���N3a��n��~u%����X�W���e���m���9���o��Qf�>����22�-Hd�{�yy_R���73�l��{}�^��4Ex��+zna~��i[[{�R��*��&��XW&bџL똜#�7����F��E.����/&��H��(+P��&F�Y�+��n� Yy\hs��`=<u��/�j���o���O�]�����uD�1���|����h�,e�+OK乘�:��v�خ8�������,z�۝[,n��@&���{,�!ii�p*��	œ4��2��Ho���2�C�TWɥu�yp�3p��?�F^����A�^��c;8� =�o�iyt��&Qg�Wp�ǝt�tAe�8���Ol��ob,�8|�u�����&�lи��m��/h�5t�?q䪤������6Q@�M��ǳ��enml�������^a���I[���{�m#�C9|��������/0��=�O<�]˾���nj{��.����N��:�|��z���%�_j�����{\��{�������?�-���	��������٣�����M��~PF��:�,lG�^俍1�	^kk����|�����N��5�j��A�%cۓ~>��3����o1����Ȫw��<��фVK2�KfW��Ӫ���{mә��PR�@��՜@��jZ
��9������n�m~�����w�f �▟}Qonv!��G=�B������`l���*F*Wv|� =qE�­ Qx��O��O4ߟ�����>m���SvN1��Au(��pOzy@�5`T��/�_���t	m��S���$\^�4q0�E����BE�f�c`Չ�t�"1�0���À�ۺ~��t���Z��Vݪ�z#����:��ⱕ�R���T��P3f�,��cx9��%�Lh$2�Bϯ��M0��E�i�ch�:�i��������W�I��sw�R���e����Bz�(O+p�ɳ*v���{�e`r��+i	�nbF%����p%O��WT�z�ؾy����Uqx&OY��W�*��(R�\�%�<+"��ty�Jv�.�j�������o��敤�ͽ׹L=�ן_��Q�v�jdi`��9��Q����� ^�(Әr+�ߡqk����}�E��U$�=�,g[�e=��n帖�;�x�����=C�o2���N�:ҔaUFV��������Gլj�[�����y1&��^���A�ֽ�,��E����d�+Seh�glhk�J��>�K���~P��<q�����΢(磪�>�{�^N��ȗ��t"G#�m|�R�طb4 ҿ��"�+�鯜�0��RΣ�i`5d�S�NeZ������S6�'�T�s".V���l�u�o����Y����p���l�,�o�yz��Ύ���γ�@y�0wܦ��Pb�a`ah�n*�c��n��]jR�;J�<�wYf�Ϩ���ety�Pm���Uo��B���M� �)��:9�)�4�c��]��P&߯����/�Lĕ�p�AB�ۆŧC[Qvq�V�*w��8�����y��<�Qh�=]03�U`���n$�В�T�K�O2X������I �|�G�C��H�Ь���-K������v�s�iP���g�k������aE��i�o��usU���Ac���@���?��={�"�V�o'7 ��9�{^� WWV��͗�=N>�Y%�5W�^%mߢ����l):HC�sϗ/���bdih;f���'��wJ�Q�t;����@���a�jJ#�sx�ʬF�iL��Zp��<���v��[G�.�V@���駟�_��7��%~�O�H�b��ܚ�G���[�[~0�M�f��Ը�LF��|�{}b���_������}�Iy�(G����:��e��W�@9ЏvS/1�ں�=o_?~Ҿ����6x(gkk�<<���1z�q��"�B^�����n�"�#���P&�Tڃ�;(���X޷0\�ڀ>��1��R�v��7186bhh\��W�K3���Pu��C/0l��ϟ�G_��F��]��C�����}J���	��Bɧ���)4�<]���OF����3�ri�h={������Gy����_��_}վ����g�����'O�`�l�=������_a������/
�&w���6\��8X�F�|��r���g�G��5#㬿�8���|����5yyXF� ��wy܃B��3�)��N��Ǘ�!8>�_;����0��)c0>�I��Y�+8�$���7��?�����E�������<���B=s���h�A�Rx.��,�;u� �{����8u�C��n�ziE�alѹ�s�(����N"_2��w?j��?j����2�� 9�ar��������_}�:'z�x�*?�h���o~�v�{�����;��} �͒&��t �+�� ��_��'ړg���'��d��긽ܤc���Ϝ�(k7/����]��-mx��s�F���T�$���N�=Q���?��D�_��;�U�J���Wp~>^�,�e����*��%����w��ʩ|�N���B`������&ϒ+����.�}��3=3��Z�!��HFpI�}]�B�(�r�K�bf Ƶ7��i}>�soU� ��PP!�V�ﺼ�'O�vbr�]�q��\�����Je�|6I��uJ���g�d�?�u����t�@���#Wi0���&w��=hW�f)�{jA�
D�*SB������S�.r�gZ䈧���YYK<�*�j���Ɇ�|�<��O>}@�8|�q�
�%D��Q�1=
�2�����|��v�M�d�F��r���k"I�i]��<$�T$�S�+e����X���JY�A�ɭ��"8�5���u�==�ɵ����}Zg0�sⱻ�"���������v��q��g��$�U*��G�w"'ƶ-���:��b��$������	�c8G��([�s����|%�Z��nm����P��������>������{���mrv:�F����W�o����o8o)�����b
�-[�-�c1�xR<"�T����aq*�́�����Ct���=�rFO���Q�uN���Q���9���)�'����H�6�����)�'���\4�3��ϖL�P�5ͻ��4>T�� -��c�� �l�-�'�����r��N���p8�4�`�E�Qirh����By�}z:6�S�r���cp~���\�^���e����j !��e�`끳�D(3ĵ��ı�b���Y�p{�lLc'q=��1>2�V�wz�V�qE� ���փգ�u��^�T�V�N�#u�\Q7Rv��ڱ�	��f]����@�i#iB[���6H؋�\�n�Aqﻓ+��,u(rg&���H9����Ę���o����`�_�� o��	;0��ג���?I���C����7�K�Q�fu�b�S�Z`���b�8���h������|���?n?��p}	C��m������������h������:#��q�0qm#�@[X�i���i�s�����/�
M\G�~������,��>V!� o�*��wm����14����W_�&f�I����a�:A�-��[�;�78�_�$`�۰<08ڦg���������V�h�㸁���l�[��8��h�!?')���lz��qB��o1��W���o�6K�;����8�;Ҷ����8F�^�WƤ���;s�ͥ ��]��������6��P���A����?|D�|�>��0�v�i핫&���19�J��c��ݣ�2�!�G��W��^� ��mzf�ݹu�ݻ};iC''�g�4���o.��3��こ����lo���r��[h.8a����������mf�r�b�\p��,�0==�F��&OGA�`�6���9��4�+��@r���ה������Pw���oϩ��F��h#��,-��nv.� :@��]wy�g���_|Sn���s�t�-��ӧ�{�݉.>r�1Ґ���S�p	��9��w����{f��ĮS^���A�7W����l8��޵�"'�ui��~M�<\aX�ߞډI����z�[\Pr�l��q��vl���Mb�V����;�2p�1G=E�b:\�u%�ݽޮ�LC/'�6��c_��¹����_�'�:Y8A'#�K"p%�L��d�*��5He��lg�R��C
{�;YЮ�b��8X�Ͷ���ښf�����;?Ӿ�ѣ�G��O>(��!"U��2��Y�S}�Vϑ:�9�r%̾rm����<����W�M��<����s�*�{����8Y�8Y{틯_��gN�t�\�H�Sq!� @�B0L�ܨ�#���3~=b�`�u�Y8r�#�,��3��ݝ����#���:F`c�4<�S��c-��ށ�	�����3�<#��;5����\Gee2�8������ڍ0޵,!;55'��ƙ���F�n ��,*$[�u���odd�tG`<��b�}m=�����W���0��Q�qa�:Ub��r�� �-����#�W����3'K�P��<��sUF�?c���<�(2�yG�Ǡ��9N�O'kp��#�����,�Eɧ�8[��9�<�[/�C�l�%'K�q#-���|�Y�@Y���}�)�����d�-�NV�{���֕q�!�K������߇yv���o�i�qM��ut�H3\�rs�����=h���uȹ}�������[�N�@�?'b�Jl����cmo����mm����!���$]'��e�jy���A{�����{��Lۛ�q���O����?G٢��w���k4��Ttq�'F�J�guX�1��[�Q>FIt��ޞs�(����^Cl����'&|�þQ�!��b�dP�M/Tp����0����x���8<�c>qH�����i�FeG��2�����{p #X�'�@2�͏vpcqG殮eOш�O``ML8C������pSF�i  M���9x����
���{����5ؠ���]�4 0@Ͽ� ��ת`�]�~.O1�ң��@�����.�|{�ytt�u�uTx���C�R���A�3Rg9��إ�÷~�p���h��E��J��W��(fda�	W�`�h���E|B�:�ټ�{����Y� 'O�{�Q����?ӋQE8Bv��Y�Y#Y��Q�k�DZ�qJ��ot�\@�y{Rt�18�/�GF�b�=��ꘙOR啶���^0�dsh`�J#�q�Ґ�����r����d��vmq����V����q��o<��f�&"�_<������������V��|��ظ� �[��ݡ��w�,�޻��Y�0+{����������O���8.n9��&�Y�Af������m{��k��𜲌*��[��ҧ�1|��w�^�@=���z���
:oj�s������q�B瞒��"w�ݸy��'?���j��2�1�M��o�n�ӿi?������]r����>\�#E=@:���j���M�)�1�w�ٛ���u|������(���`��э�������}��G�����/�ۯ�����'\��>�S��[�� 7����V��✼M��<:3��q�][Zj�q��o<�B�]�����������.%�k�h���PV�������D>n{�����-�._q18���^wO�}�Xϐ<7$��3/]WC��f��|�d�ԫ�ˏq���	W�8W.CF�yV����޿�>��i:3�����4#?t��󟷿�[7��<N���\,��I������K�/��Eg/�:M^�PN�waV��	>B���͢ރYL<\�Eo�?(k`h����\C��um���"N�8s/XuU�z6��P�6�0e�b0�ۭ���~���vB{6���a�O.?�\�\e�=��m���a{���67M���Q��m'���}����w�v�`n�KJ��Q��dM�ɞ9Yٌ�<���-?�X� H8:�^�BQ|*K������?��&v~�~��?������M�]i0�-�
0��s��n<����{=�h��2��Wbv�� �*Xӓ�8�p�����q��;P=Y/�ڗq�^��d�S9(�#e6p(<t �xF�&�}	o~�0d�,��d�3?������t���EN�ȕ��B�&�4��A:�¡�����W���=q���0A,�iA�2 L-����� p:��c�m��r�N�u����G��8m�E������HG'k|
�P���ٯNo�^m�o��9v#ص��-���
��R N�i�U���)|�o�ĳ-s��C<��|��J�Ж�Q��B@P�@�p_���Rm|���i��g���Q��a[8��B��(e
ᜒ��3+��dIU��pVu���H>�tG^���wY͓��7�%J��(���tu�M���&w�+��>�\F�q� �˅Oœ�<̰�z_1������t��\G��|�*x�����⽫�UoF?�
�����:Fж�<���~�=����8Z�he�b��+�j�[f��� �Qr^��w��<j��A�q�&2f4C����p��&N���Ri+ƚ(�� �K���S��?ꑐ%���xѰ8�8����3�֖��c��ڊR�t7�\��g��"n-�3�q�����T*b�����3��Tr��:������G��3�N��{p����(~h�ol@��������V�P8���XMN���)��Jb1�����5�+[�k�ۋ��0{�&���	��S]AMCB}�#'��,5����&��C��b���������p8wr4���2��Ic&oU���8<
����=���{��1��"ZV>��I>:���.��4�*N��NV&�G��0�(���#9� .iV�SQXn��E?Wީ�KF�ݲg���ʽOM�Z;��q����dx$�#�P���CʐS�%����������虗�$M	#e�D|�|Vo��(]8�Jua����*-W��'���������h���az�>���v��|B��춯�~�����?�������/��)V�H�c�ZZ�d٨0ɳ���G��7nf��7���>���?���#3��i�)e6���7_�^<��9/�aX�SY�<�; \%�ذ`W|�j�=��z�֞x�75�@|���3'kkk?���ҵv���v����dde@�c̹Z�Y��D;���g���E��W��z[�^�.�SmB��r�JȐJ�y���E���Ξ,�DC���yl�v������滷�ڿ�矶��~��p�MNPV����F��?�U�������~�� �=��n��%�l���}�R{j��8���t��P�"�(;��}7��M�u$4�	�l�~�@W������*6�x�a�yqS��H:�_��Ŕ&'&#w�}�~:���.~q�W��\���iE�eO���f�pnё�;�c{
uP��t�n޸�c���'���8�Kmj�����`w/=u?���i?���h?�Yv���"�o���jcaec57E�Z.�|Ak�q�a�<�0F���py���N֦Q@��3�<ӝ~C��]���!6��B5��������ɆC�q�6�N���d:�pv��+��Uy�\�F[�EY��Q�,��r�ƅ?x�~������]_�v _����?�?��Z7'�������5'K(aJa�O��B)՘F	ϖ��9~�����t>PV�:v�
��(�.�N���+�!�[=0]	^B�-��3�6?��	��)���"���[�.i�'�/�5:��7�<���"<L��.BǱ�'�&|N�<�Ċ�G��S��%�~�z�1S<�_$ ��)�Ř��}�S��V�^Ǳ���:>�]=o��mp��?�h
�`��E�Q%
^e����,�@q������}�d,B�W�=H<���q���{�;C=)(F���$�$tq6� �e/�ll�Pa6�J�Q�� �~ΰX�*c�F�+*�R�u6nzay�i{ NW_�b<1�ޖ\��~�庫����˓��$_����'N�<�^zVT�"���܁X3��?�U�ϟg���A�_+�����ﻣˣs���J��(��y�Z�����������r�z��
�*��}[�<+Tm�͞:	�� �����Q������/{�lI^XZlˋi9Ԩ^}�=��qƀ�~�*=�\�!֤9�/
���6�|(��˵��˙�r��S�B��"W���t�<�ե�7?L�K<�K�U���Dy�AFQ��إQE�}V����$R���IY\���g�fØ=�e`#��et�s��ɝh+�����B��2��L��+3(��vmi�-�9�92�R�Isx:�`'��}�����;��cmgs�e�h�3Y�xv��Ϲ7�"z�z�u�v���}��v�����oc�j׮�i赶�`#�"2o�MO�e|�	t1��e�������U�:F��X�\�n�TcWy's��0��G�1���	e�s�������J�����qPuDH����;�i���~rx�,���ב��:�:��h�k$0���1���K;�6��m;����|G��?��E�h'��xeE9���t��������=Y?�b�Ƈ@h^���t��\��]D�,Q�B��_^�\�j�h�.��d��{������N>_eH��?��s���2<����:�����
�!M�@���΃����*o�C�����
��h"piNU8����U����k������^�i�+�bئ`�F����:o�7�~��mx����q>�7�u�wW�s��ܜ�b�b#`lj`��p5&����q&\��sg0�&K���6$���k���*W��zL���:1�8������0_"����{8K�N�=:�j}��uO��j�������۾y���v�M��od>՛�7���=�<|ߵ]������gCg��C�^���7o7�Χ=��w���"6����m�f���]��/�5�m�g����^�����8L�V��4������Z���L�dٹZ|������
�{�s���k`� }{�Ź��v���A�Yl<Z\Z�i��f����Ed��O�r�ɗϟ�'�|�^<Ҷ�7�t�U'~ow�l����Q; $�&|� �3��Q"�W�٠��͹����QD���.�N��|M�Q����A'�.��m�J~��a#,!���mW=4_�����߽0�cG;Z��w�qK�r��ؠnt$�#��'�>�eo���R���rh&��y���������x���됄C��=��{����:���~`:Yah�w���_�E�ô5���d!K%�A�d7�_C�,�� �h��u\��2j�~'"��Z��J"Ɍ���OG���F	� nVoA��4�U_lo�`m�d9	� �ٻw'׃�Q(C� ��#��*ϓ�?������ۊ�Pyy��g\��ɟ���"O|����S6�G#��{�(l��}���bo���&EvA�!8�!���@��Y*5c�1��PJ�Ơ��uZ�/�Ղzٯ�����@Vp�%ak���a'xdd,-���H�-B��qH7��&s��8[�TL)�h��21��Q���g�{�r�s�LLq�J�Vl'�,��ƴ�I;x��*�5J`n?�+�)Cン¿�S�q4F�z:�vn���@�t.��������O^^ֻ����S�..��U��l8+÷�:���7�>���� �y\L���{��C������=��Ѝ,�:M\h��}�G��sV#EN�*hu����_��Kep_�ޮ߼�V�]K�-{�;��ɴ���-�'��K�Ka<$?�GbP���Fe���$%V�y�8��}[��U��P+�V�6J�&���~wM�>�wi�z;8Yi54�3���dKrB9Zg����*��y/�H���+K\,��.�����!�i��r/"�C,�{���]������v{y�-�M�鉫m���O�Ƚ�=�8{*�6�!���C����S{;�'m��lc�lm���m๊��Ӷr�ݿ��=|�^{��G�N��Ç8Ww��;����mi�z[\�ޖ8Z++7r����#~�y,s�nT2�z��404$�á���zD�%u8� 4�E�P�����`�H�]Fl�ɾs,\�@�Օq�\��!��tZ��kX�=�����e�h����=V{'ߨ3e��6H��d����+:��I\��w8U����J���\�չ	!��&��4)�h�'����t/�˻1�H/4&?o�h���i������>߄�5��y��v:P[B'�t��S4�v%�y��꽻nںB��Ȯ��p�/������_�M�����Xg::X�|`�����ެ9��,��jn�oC�<��a�6`j��lݯ��7�4�_b�on���=W��Z��tƽ���Pp����k8
�;�g#v��Rx[�w��\��Kt�\hn~�McL�k"=���h��S�c�k8��'r��C౾��e�C�L'��pjo���66�/r�:��G0s��wdO��27Vڇ���8��6nX�=l�W��ص���'ϲ��p�Se����^��u�����X����T�q͑���,�A���mWG�'SG?� ���	B�x6_{��?��q�[���G�R��}��w�����5����lϷ=�5�&24���ƹŠ�LN��_��V�������N��~cw���OC{v��\}�]m�������G�ț�8�Q/�.qޫ���S���xг�6��m5���5R�R>����<O>����P�Wڲ~�q�T�t ًe�-i��@�#0��ё���x8ψ���P��v:8tsd�.]�����n(4�۹���[�ndsf��r{U:'k�=�ɲ7˞�C�}�+'��+�hq�(D�;�����D���`�0�j�TP�2Q�� �~#�x7Es��e���L�Ҍ 2��m�#-$=r���qb�hA�yC�5��y����'
b}�~uA�����*'kG'�͉�G��E�T����ͅGwM�T��e��/A������sQÎ��`�<+�����wz�t�\�"=X�4��b�''���:�t���(�H\!R*Ϝ:�`2.�����4��R�����XN8�����:Cx��B�*\e��ѱ8��5�����^�/�YX����1^��)�%��ɬ�TB/F4���9����cXI,&����r�U94>�@V��:zM>�T2�J)�JB]]t0HSүx�U#y�БXrKK3\R$f��{�ٲ�g�?��^,�	��E��}���g�_� �֥W��k/�t~�x}�Y5g��=ēG��Y��!B���Ht^b�P��4xXO��H�a-"x�/f��˶b�S�(��P�^kP9,�a<�n9��fz���˗/��o�nO?�p��Q����k���=�!�����>���4�J�T,��A�Jwεf�1�}�ݟ�Y<&��!�4�#����K��Js?��s|Ky2|��������A�X�(��z"�Im�3!�y����'�k���|��G��D\m�c������{w�G�n���^k�V����X�vIu�=o6,��Tm���նM�ùrY~[OmhC֨,���v[d]�D�NLN wn��}��Lݽw?�,.�����6=��F'����D������Dg�(�e��qRGR��Ju�M�ε�)[�1�4:��5���ب��0+(Z�'oK���3���1<��+�<9�q�&G��Y�Ź�47���Н�ae����.�x�@&O���i�'�M"��+�9�(o�S�(�#�Yp8�6�\����O%��M�҄v�!�Y��$��/ݐ���y:#��a��˵�+=��ޔ�9�3��4��"�Lױ�a���cהּ`>.x�w���6��ݟp;[�rc�充v�6r#j'7=�Ώ��j�������ز0Mt�zM>�0�0�w����4�B8Y��A.��_X̰A��ɧu�3r�`ғ��=�d��bO֎C�o�_�	�2���z����&�.\��m����c�|%=3��� _.��X�b9T��E�kǟi�����zY�$�:��h٫����"R����Վ̜`�����Α��F3<zpuc�ٵ �o�p͛7�ڏ>��}�ɇ�.���|*�@�K��<����ڋ����؎:&Ҧp[?��"W.�e�ݻ�~	Ms�n�����L/��y�)5�NX$��ï3�2dA�S�"+;�K��!A:)�@Ɠ��l��q���.�SKG�z	�����Ao;U!���8I�Ȗ'l�F�r+���:�nݼ��g���|��b*O��/�y��?kO�ykk�q�|��Ae�|�5v������wy��Ym-�˱�ftA�8T�����u�q+;\D���3�ʓj|��
&��!��L��i��HF~vt\�%�"��2TçrE�+*�#/�G*Bꁐ�R<��ccmaхa����<N�C��#�����h��mS���j�	s"O�)$�ǩ������I\Q�J�T�
�{��G|�O&s_�tT�qU'�9�p!��"Ac]"�	L�5��V].�e�q|�2���l9�����kA��$*,���l�P0N�Ȗ=Y�G��p���wK�*G��b��-�g��J�氼�.'�z����K���g��`m�����{E��]N+��|ch�{��*��u�|~z�p�n��Ǣ�.����!�rH�^��C.�:��m9�w������ü�ji � ��$U7�S�f�	��2D�(�t�m�v���{[ܼ�Ԗ�lͫ�
l��C&��K�X6���3�'��S@��}�c�� #"�c�j�ы��CA��0��WpO��gzI(s�
�R���ą�9U�u�;n��#� �[����㵾U�T�������ۡ`�^�8�%4\we�I�{^�����������U���8�^�Xz+�I8��RW]}Ep*�l�R!;�UC�Q>8<,� �ҀC������[*s�	޾u;��W������LNPw������oå_#�#��U�yX�}�@z �4H]��@�2&�o2OPc�2dO�ʻ�
�>��;���:q�&����*}����1L���I�O뷊)�`�B�!a�P�>����̧"�U����+:;�v�F������� N^�w�ߩv��\�w{�}��N֭v��B��B���e�A��P�l�űZk���o�d��C �|\X$<|Jn���x��:��y�ޣ����>��G��?hר��%�K�a��5��ln��R�qN�΄��(�{�fgk�����8[��1J9�qoG�'�����u�|�R�Y�(�;��5{�t�\�W'kzl�-�L���6�|D�`C��T�U�r�C���w������Lt���?S:RQ���2C	6�b��ꤜ�!��ٚ���\�ȯ���~�K�Z�$��	�G�$PV�>qt�-��ҟ���)������F��-���r�	li_��Up�0��^��5���q���[�H:1B#���-��,.�035�n �-/d�~���t�mo�/�x�!��o7c�
��:.~��z���O�3��37S=YYY�L�wj�~>�_��r��ǯ�q1��M{���(�j<]�SG��O�g�r(�K�;���N��� ���Dh�9C�=r�p"��ǡ���ٌZ�^3�z�6�w�YG̡��P�e�[k���E^l��p~���(��g���o���t4^{{N����Փ<3=��?���޿��l̉:'m��ry�g�^6�ط��ޢ���^��{;��UW��{�ĝ4���>p�%���\eoF�؈�A�����'��8�6T��C�q2�:O/e�y���9[�} �Y'Ȗqd��!�jG�ԩ8$��,?��x'�\��F�?�+�~������zv<mei�ݿ{3K�� �V�p�~��/�g��Y��~���8C�0ih��D%=e,�}l6�_�m���$�~��\}���E։�.|[Κ��������~�_w������x���,s��du�q�&�4��J36��Z7��֔����LVj\Y�o���Ԁs��W�ŷVn������b<����=�.��9�Ȍ�Fq����3�/��b��\V���:4B�����/����������������_k����c��1�	ypwk��WF��+pzm�[����n�;wG������q�E�d]��ٹ֜�g(�"Ub,:����~�`�2���<����©�=��X�M��k4u��N��M��ۏ��1��+W"h8��Y�	d&H�J�N�S�u�"xG��|�^�t�us�ݺ5��5���_j<��>��N{���v㺛 ������Ժ���.FR1r�7ݰ�浆���BP�* �k�%亞Wʭ�Q�a6����q��9�J�,xv���`e_e\���I����2���/��3?y��b¢_���i��	yޅG���烜����G,��9��_�u�^���a菳|��'�/��S�s��I�\
R#�F �iP���w<�*=���d��<㊙�ܬ߻*�K᪔�3%���J��a0� }�|3�8�� ��G������/l�H��T���OZ�Ut�w5T[��<]�)Wʚ��4?��>D�;���
-���!Z��A�А�j
����	��y�'��\%�ߥ�x��t�$�ڥ�-x��-���wf�'�l������O�j=���^h�0����pbW���_�h�8V�[�	{�n)�_¯�n�K�S�vx����v�.�jw���L�u�^{����O1�~��v���m�ڭ6�գ��Tc�T��4D�9�y��r}t	����� ]D8D�h�r>vq��g�3m`|��L�����{m��n�_�զ����<��x���ӉӠ�aS��Ni�J��z \ ����!��(���aG��S�S8�s��E��
��M�E����27�v�M�Y�Q�~.�쁷�s���w����B��pΊ��.���C�:[���p*yCE���K�y��{��cp��2�N�L����a���=�����ư�Qq��<!�J��ҶF�N�˔�]�Ј�`o���o��E8}�/P��p6h�V�Od
�	��憱n�����t�x˻�E=B3�Cna=h�u�:�*�脘n�@�/�+~6�#A܈��n �3��^xX^�O이�:=�Jy����\j�䈰��9:)���q�~_���	 �8َ xw����Fv��2mD�D���`!����@�ƿ�S�.����IZס;Д<���8&��q�������7����`{�z���h�tl�uێu��=W�ù����3�h�R!3�c�u_.m�Ap��v�eh�������]ay�e��>!L�F��xgfp��A��
��Ӯ|���Ny�1�r����i���QH�Y�A|� �#ec 6�{����	�9�`���q_w�?b=h�Q��@W置L���T�Q����ӧ���?o���/��8Z�A�0y7�u踎�� �#���,8F�ؘ�Y���yV�X��	��ɒ8S	�ql����7��4�9PI[}k�4�(M^�m�TDZ�m����?�<��o��%�o�F�f�1{;�����/+Ǌn�����_���ye��}�	G]C+\�=�?�ߎ5�1^����:�O8.�s�vV�xWw�����f �1�hW��ﹾ���e���k���?��������~򓟴���n��^�|�K<5�o)����j=�:��F�x��/AY���r�=�x��w�.ƻ��µ���P9t�P=
�~�C��+C"�,�d5&e���CB'�a蒧�׷ziHI2�!��QQ)�4�l�C�v��
�ڽf��`�c���շJ�k˔{m�!��#mv�ea�������e�5�����8ݖ�p������h�heȢ¯Zi�^.�_�L�7
�<��N8�&|�3��N�u�w���d.��^L8X���װ�����1*�R_�\��ϩ�~�������>vl������
y�?�T���^�'��z������Ͼ�δ�p��O����7�o��S�z�鲗?��Z�I��������ǜ������_�.�!W��$>�^v�#���o��W"|�둖d�٢�+�TW�QNF�;����1��m��W�G�k�0^Z_;T���/��L��ҟ�w�޺��}X2�<Ja�'¹�(�bf�Ζq�H�a}Y�:�Ş�Cx�a��9$p��,��w���n�~r���{wۣ�7��[�my|���f�^{�V��^>�M{�����+�Mx�S�>�����%F c�y ������T���^�������`�{���p�Z� ,${�lt�|�#q��ĵ����N|��ᘸ�Д�
����ӫ���\�Yi3�7����@�[��fV�g��Թ�v;�b���t�V�h�l�`��'�{]�������#W� ��aP��t���m���񦐕�Sc��<N���	��8=��u<_��:mW1qz\'��+�?|7齊é��Js�8[q��&d(Ut�	�+u���C8ݧ��C��;�'N�p��a��θ�H!q�E=���i�}���le���|���Vz,>֊��5"����~%Ct!C�x�c�'�F#�FCyS��0R뀇�ӽ=1ܷ���Ͷ�~�]Ҹ?"�}��ԩ��r@��urD����<�{���~u�4����SAy'[�P��G���O���\�NY�&otVS�����&�اib3�"��MaPFT�:��m/�1��`mC{n�*<6P�0:,�o�E�b#��d�ud���d�"���Fdt�<m)�*8�[P��b�)+6��O���I��o�Z�u{M]������Ջ�m��z;98��5��G����A��82���/��O'/U������h`����@�`��P�c׌����v��J�|���Y�𽇷۽;72�t	g����a9�=��8Y8��Qn1t��_��ҿ�8���W|�?��}}J�.04
�ad�8W���u$��ˎ���rA�o���u��/~�>��g��~�޼|��n�:�h N�+��:u}��A��*��`���8Th����;Ñ��C<��*�����^�E㹟�S���3�� �AF���0� �c{�w�; ?�f��A\��Yއ�-�zS'Q�v��}�fH�r�N6���b��r��Z�C�A�᧰,��D�n����]<3�B����>�ޘN�w�R����ef�����onl�a�K��u�ٵ����N��@ n��pA�F|�5�n����
.��	s`��+�y.x�g�eltϿ{P�z���d]���{���:��G��_�P)se3�J�����(X��(��
:�Koq�$��8O<���Q1�@E��p�_�����~��J���"���zg�b�+�ҥl�^�H�(5�c�������/.��lͷ�7܋Ca4��5���ϮW�gs)�ѮW+�Ӟ����W(�B�"φ8P�j8
5��ǳl
_Yn���U�z��n8����ǸԈ��e$$L�|%��F/�����q��]<�J��.�.!�\ϻ{�OZ�^8]ȟ玟��kB�����}F�y�\��?�����\W�>J�h�T�>�L��W�E`��_[UU�:@�Wc���Tg��y@:d.��~\nĩA��b���әܤr��~�=�V_�O}Q+/�e��a�w�����|������R��\������	|���k���'�;(Wnr�r�g+�Z�i�Ø�UϞ..�8��e�����ɡvmy����F����k?��C��{܍c���2=��5��>�m{[o���m��7m�Փ���%��z;�w��Bp�Q�0H���NQ)G� #��s<;?�n�Ñ������{�k3��o�H�(������p�!��3��ժn@���n���︡�4�����6�C5����Wn��k����;mq�f��m�p���P�f�x�s��g�}��\��o�b(�#/g�e�G�c�`p�@_�Xq�����05�n.͵;�2���R- 2�p䰫`^uT ��=�4�3�,g�z8ԩ���N�O#doGc�:p1�}@v������d�f(�,s��˟�i�.A~� /H��ق���:j8\��q�}�"h0�%��S<sDC|{V0V�0N�P���jq���Ս�����_}��������g?�U��/ݾ��I[_ߊ������C � ���L�zs��z��}�v����/N��#�:��׹t��:[G��*���q��.��I^�m1����@�6���yK4q�]����u�dRn����M��w���D���o̞�Џ��q'&���Ts�{�Ж΁���$��w�Q�$C��o�jV"Hk6�f�ׯ��Ʋ��C�o���s4Nm�B>��	FT�/u�C�m�v��+}.�S���ġ��>��>N������?��'�_��?n���ÿh�ۿ�������O~�~����������xDf�1H��S��ɼ�7�;�Ydj
�2���7%�9�򧒌�\ N�/yH:�}�U��'�㶽��^<{޾�������������g?�|��ϟ�m_D��������.�G��=^{�]���*��d��zt��2dYe�,�E�̗{�ѹ�3���{֤�؟���8Z��r>�!i����f7�ׇ|sH<������JY�w�R��|�J�6`����8��F��aM��FĎ�{�����?w.�K]>quA��@��	�X�R�4H�ʗ�!z[�v�r&����J�z`m���M���F0R&�g"i߮�57]��ti��1`F���o�_���_~�^�������=�n�-�+ח۝{wڽ���4F�-]�� �\ڧv��N��rŃ���Kmc�n���mc��HZ�=��+C(<��Av�V�VX=dfҞM?wF�kٴ���9�u8��k���C�\�"�/k� ��-	�T��R��T�[f�]:�!���˚^����@�1�g'�]��`"g�_i�P�j����8��Xc#��!�>=1�������)� ���-v�CX�
,2�"� ���-�&��c�k��mjjŀq=����N`��=�	c_�GM�t���m����/	T�5� j˯-d�|���6[qm=(��(9L��4cd�4^C ���ܓ@
��7�!0�`�k>T�����m~\�Y���)h��\�`'�F�-M�#<)ۜ��?�r�=p����@Y����;S9
��=	��>|�^ةSpח�wT�3�2~]�a9}0K_�|�0����;L�o���ַ��`�%��i�$���V8��3ot�M���,��p�t���]	Oa��X���.k;�}_�c:���n����M%m˞U�.�X����w�C��p[�y�`�>N[��z�H�|!���_�p�ϱ�D�`>0��3� N��
��u��������Ud�Y���<
ZMu�ex	�}��`��2<�3�>?�X�;�8�
��O|�q۠|k���F��dȯs/��������ۣ�����x���m�jo_=nۯ~�6_}�6�|Ӷ�>���v���?��#��	n#��mX��2���U�7<wby�9�݃d�v�anf�=|�}��?h����j�ݣ��1�������$�8���'�O�ԯ�䝘��'�|��ɋ���6h��X�>�uex��C�na|�r��ƛv��3WJ��Q�8����Rp��pe%<�!���e�T����D$F����la���St�%p8D�c����@�q͌��QTe����8D�Y�~�����3~��ʐj��C]˄�^:Aߧ�� N����*�i��b�<�!F�4(��O��[��EW�O���v!�g�2�4j���r��aO��_j�gu7�Kп��:�n�O	����\�A�@Hy�k#w}'ok� #�q�ca�D�_�����h��<�ۍ������Ͽh?��g���|�V߮Ʃ��Ё\���.sԅ��I�c�Ч۝�������sLnI31�3�[�X�,/�	�t:���u)�u[xx�s�Umt����	��<<p�<W�;l�������|�>ש�S��qN�N�$�CW6�f���0N��!h�$�!���=�3��mzn�:�����/�o���ac��]�m��po7�r����,���hGhkK��;��ҁ��3d)�f���w���ڄ��C����n�%���VۗO��ǯ^�5�����lQ���ҁ�m�O#FF0��(��g�!$)��> 7��48xp�>�{�>v�kK8\��_~�������p����޿��޹ٖ�\Ƕ}�r�mn촫ɸ4M���-s�oh�*ϑ룃��72� }F�eCa�=��h�Xڤ< g�S^�Gg:�Y�w.!S.#+��\9�BC��������W����}������*�[:)�H�qִm8gG��u>�������{���0X��I#�-A笝���<�gJ�����l�x�w檱��6���<��ô�U���D"�lB�'Q���'�m�G�kfXΠ�B��G�m|���,����R���@������ß�m�d��.xD��d�`�2x�I$�p9tʉ��C���FDU+�� !�������a�繶l�1�."ɖ%+n{{�=y����ן���_�t�-�s��q�+���-̷��=h���G(һmM+� 2�^"����3��? f���mmk��O�Vt�v�L�9���ā�VJwT����=.��:ξ�Gb��
�����5�#��UdJ��k�"x�U�!$�<��hlJhԖ�/��=�Y��y�sI��A�
j���K�ڪ��X�*��:F<�d����p��c(ں�`��/ce!X[�4hN�uú���Ult�q�_(��
�9F�d�_������õ�N��T8�ZfU���OL=�H���#F�o��G�4 �����}/@���M1�l�!�h_^���W�0]��H"��#!N�q�Ϫ������ག�;�����8I��8�}�Ξ{���"�q}�������x^���k#��ż�2KȽɝ��Fҩ_&J�q�<:b�C��uZ��9O��[8� ఑ݝm�p9#�hH=�
ij���O*
A���9Y�#1�FfI۶r��� @��Z*7gtH����t��b�:5�� ��l�c�?[�t�z'*��NR��V�T�i�g(��Ƿ������ ��Vy���Y����mq����[�1]y��"1D�K�G��E7t�s�V�	�8/�d�}�f']%p�}��^���w��A��������1���A����,�7�x����`���GǴ��`v<�g+�~; "�f����[w�}����fA
<��}ėqC9+�_���������#v��?�y�!ŇF�J;)�~��zA:�`;��)D����z �y�β���ƃ^)��G�Q/�˱��-��Щ�5o� ]d�M�/ƒ�׵�'؋�q\�'�e���P�'e&��S^�����3Ϥk�[��}���r\�,�'�*�O��JW�����l�"��l&1x��s �#xء~#͹mZ�Mr��]�B��s[�"���(��3-^��ao��B��X�a��\��
	E���ng�t�N��ql�׮6��N&Ω3��k�!Cځš^�7�ڠ9�S�g�zuj8�r��Aʎ,�ŷ�Y'�N��@N�6���@�m!�leW�W���6�omi?)q&��[۵W���&��1�S�8{�����%��� z��Ü"8l\��ͶG�V�PWq���S�/۳/ó��^��llp/)�Cg7�Pv���FV��ƪQ���-xf�����XC��k���r�um�M�K�`d�����I[]�jO�k��|���n���mg���:���pb��X��b�i�B:�ewgx/��ىؚ?���S�v޻Ӗq��y�0�n޼�n\_i��Smzf"�%�`=51�;�R��L�M���^��vx[> H��ӎy���!P��Td	���3�u��V@�Ï�SLW���+��9F��Ӯesz������)4���}���`[B��V���$�%�����in��{�'6"����N��盺���r���8��ɻbՑw�Q�UT��.e�0�<�G�O:.�پ�r��Iʁ�%�g�iOփc��67���m~ngB?^p��7#>Dp���Qh�܄AAak��֡%�
�v��:Q�Z dI u\�-TV�ޤ^(�{��)�C ƈ��i{����o�o���=}�mmnS�&ˤ5gjf�ݽ�}��G�����QE���C�H�>Ғ�X�n$'�'� �v�(�ݙ������N\<�{�1�s����|��AB�Ȫ8~������Q�vM�fȚ��`�*�^:[M��QZn�:
��9W^�祁l*_T�pl�à\QP'+X�/�,1��֕s$d�t	��(x�ɪnS��1�{ibbl"N�c��m��hڥ��٫Ɏn
缳L���2dR�w��d�@��o�5�j����]ŇI���2��x�$�O\q�m&���,5�/<R�O�-t��8k[�9?r���\���ԙ�#���B�1�
�\u���ĵýL��\�?�y���9"L����Ͽ�#e�����o����i<��I���#�,�[�Y����j�J�R��#R�7iL�A��c	��[{k�G�a���fm�ʂ\��B>��@'Ǘ�=m;�g�P6�|�6�ꡱ����-�QX���;i52��Ѐ�ՙ�EP������d�e�W�U���,�q�A\a��4��S��e�_娆��{��g�+�֋���P𲱮�'��+>+�K���
���675��\_j�cx|�ރv����47�Ɔ0~�6�ƛm�����B?�hQ�٪ZN��h'�s��\["��2��Q��PPg��y�Ɠ���L�̶k�o��w�;���eP�A�}a�e�E;�<9s�ȏ$p�γx7��đRNk�/B���ĥH�	% ��Τ��C���:W;���;�w
�9�hvH��B��U��ּ�G��Й�_��c�%F����2�op��!Q��p�+{O��9l4����n1=e�嗾�t"�ĝ|T�(�$�i#��N�Ys���F�O��u-�H����hlg¼xla�����q����5I���m��n�ob�y��I��|�=���g����|��?��e�	 ��6\���*r`-rA��HÔl��Q~�����=�D��$��/���lS��Y��at�wa�
�x�Z�W��@9'�׻��P,���̜,�C����6N�2�!}򖋰��6��jo�.�U�.�(��e�c��1Q.���v7���iV|��i{��	�r��(;���r8��L��e��j/�tu"�'s٨Ӧ#;@ҹ=N6�N���-��ח�H�بii��,a�mn�da�>}�ެn���ضҢN�����_��Y�f����,@O�m������?����~�>��Q[���o�S8U��9�.��xPN�Ώ�>���Ȭ�;�@ڡ���MG��e��޴�3����R%�E��g���x��_3y�U�t���W�#O(�E���-x��kk�s_�����������4K\eqx@:���м3TO{&oM�4N���߻�Է��u���)�+��Y�^���I�;��79*N}w1�dɏD�`
X��+�1W��?_��N�N�X/y nt��j��kg��x�\Y^���ٻ� �����:YT�i	:Q��Cf�pF8)�]࠘TemeS�P'�/DLp7x��W0��c#mY9�'�k�hm���W�Z��y{��e[_�cIt��GMʹ;�G~�����l���G��c�Ax��S�����ow����w	!q�OV9Y�d�ӓ����|UO�G���:K}�{�X�9r�j$+T�1�&}`HW&�!���x<�\;�C����9Y2K�R��/~e�)��R�N����|'ю�߾ե�/G�[�\9Y�:�R&8Rw�o�j}����[珡������h9s's���ug���8�k/4���P�w�eW�; �����OV-�  _1(b��c+�e҈�0$`l���NA6	X���g�J��T�P5�c2���[��dI�(	�v"��Yգ%����)��;y��o����?
�ЇpI�yv��C�]"��}"u�]�n��J����:u�]���G���@;��w����q�Ԡ���W���J�[�՛�w�+�� v�p��j 2�B���Ri8/І �� �<ʭq��W�Ώ�rMDW�L��
�����������8Y�"X�l��1J�,k�����Z�ԡ��[�#�D���Y�M��$J��z&/�Z�9y�N�s��7SO>�ly�ҖW��D�^5(��U
�w���w*h���!{�&�1tf���+�;7�=7�\�o3cC�2J|o�m[{����~�v7V����rB=�.yg(cǓ)�q��(�֕#����,���:._��nܺ����[���$eq���q�a�r��C�\��y�B���g���[d^�X�s���ީ��3	Ĳn�ho��s������u����~�^�GZ.�Y�JC8�8����q�����\��w�RWD~��s���8�ܺ��;�Jǵ�'$ǻ�	�%�"I݈�'�I\YW�0�R,�20_����\�c|�̣j�ɒ7�/�I��W-���OU�	�P��o�&�S�r�0ab�L-�T=�~_�4�-K���K�KcA�pE6��e��j�:�N�{f�����(�1(=;=Y����qكj�����W�g�^*�ʽ�4{��_kb��-?8�g,�<���\�@k��}�2��v`���ޅ\�ݡs��J.N���3'k(��J:y[�M�)�8��>z��"6�]2]������
�P*@��ց�կ��H���ǖ`U���!�9Ls�S�1T�������٫���������S��S{�z��Y�!���2e�	|��3������Ǐڧ8Y|�~[�>�0I�A�	��!xV�N[iO�G�>�̀�8H��g{g�z$G����(�\�륓���?|��
"�]�;�]� �9��:�[�m��'����F2������6��F}y��ᮃ��� ��xm��L{���)���KG�H�)�E���`�J�����o��)G���+D�R�J��R��7
�����c��@�aC���8L����1����l�0ӆ����3\�9Y����SsV���
~�<(:���;u��������`=C4v7kԋu�]ضX8�YS���wp��Cql!�UC����ٹv�:J�ރ��'��=lKK��"ӂ�1�2�0	
�V\�qD2��Y�'K'kO'k紽�8J���6e��B
��UA�DLX)����GOTƖ�e��\Y���̘��}�Ye�3����dG��q6]R<+�y�����Ӑ�.�F���54Ľ��`�9@��z���)qχ)���L6��Fp)����:�?`�Z�P�T-f	�q�#�N#(��~��"�Q'�7!����*	ǋ�xIZ�\�a������jG���4���(O[ �!5�3� ūM6mvH��a��*�ac+�b�Q���	��+�ِzQ�.U6
����N@�������N��K��/G�U�mz�=E��wם�����F��w���w����y�%٥i��z8�gH���壳��G`�Ρ0����q�|�+a9;��U�~.��)_ۓn^i��l� ��
��ނ���Xv��ɿ����� |�+i7N�=�8X���k���z�͛��s��m�Ei��{���
�55�x!����}x�k��2I���z.n����)y�+�
}l��FY�6���P|L�*��B�d<���W40:�\�R�!�O������߿�>~x�ݿ���'Gp0
���������'mc�y;��n�����`�v_'�MK/�'#��l�"�(f�C��Z�NL���%����v��{m���6;�Ԇ&�S��)��%� �x���C�絵H�.�O]u�Px�d�g�+�k���WŃ��Ş�7�U��X׹�r̼����G޹G�c����.�H&z��U������<g*CgdeH�F��,:�<Cϕ���[����p^����(5�\T�.�4�X6�	�UK/y��<�7p����!��C�<����?����R{�|�9���	��� k�1X�ieS�dU�/:���tH'��	��z�����Q�p�:���J)�
��Ti	+��
-�;� �@~J�߫��(e�.�zN:��;�Y8��Q"3Eƙ�!g�j~n>��9T0��u�a�P�u��'(�=W�λ�G�p�d۱5�HY3�̡z�mr�İ�h׾�v��.��� �AtN�+���i�����lcc]O����q�[�mݽ����kcS�k;=(�M�Ʌ^�g�z�t��7��!�%�t��&�6��T�ϼ(=�-9Z�]��G�YW"v���q�\�+؏G���W�����-蓺��bEn���*h%����^�
K��˹K�3��ѣ��?��}���ڃ���������XM!
=Xo�?|;��� -^uf�G�"#�;=Z���)�I�C�CT)u`C��w�E��Xz����[I|�>�8��q �v�����������Q>��S6�#c˱Τɭ�l��lXz��9q�-�=��E��ӊc=v<nZ�P#7J����/�<r�g���3�X	�1%�[w\%���z�+y׳|a}����>���H�����S=�%O+�e�DN���/L��M�'k:��f�?�����NV� �_�4�$#��ӈ�'K��ɒ�ҊdT判�*q5_9I�d��̭�%A['��	O����j�:����V��A߭[����ڝ*�Yx k���n�ի!cW�8/�P+�� ��mk먽�<���]�d�p�3'+�&aS颢#�����NVUv_���X�mE
�%��xY
�՜�^�6�d��û�s̬�9��r7=p����)�A
�"�0��؈���[��(����\M����,@"��� j���0��㪆��G��o�V��-�^}��br��Fa�u-*1ru�0��p�����QǺom������a��8�5d��+	�!/Y��b)��U1J���\�a>��u���V�r�Қ)J����֯� �(x��{$�<!N=ٓ 3�+X=�����B ��B9���&��g��� l��]P`�S�(4gZEk9L�2ɑ�ʄ$�|��T/���Uz=|��?�a���<�|s~�n>�e�S�	�]C�\�L'JA,�����zd� ��{{ke��1�*=�
;ɵ�nu!hY�d����YMDw��gU�C�_�y����8Y�x������N����{��PM9-��J�U��������
��U�w�W�8���Yy1c�)��>��~�=$����2�8S.rqc{ c���mj|�-ͺ��|{x�Z��{�ۣ��۵��6B�w��������%�7m~nG{�u�M��Q�KLK���*X6V�KqalJ���SR��J��`���V�ٹtÝv��Gmn�F�$�Ɣ-Ãq���~���U����OVA���]�������՜���qT�ЩN�s�t�����#�{��*7� ���j�+�Ў���)Ԕ<��L�z�Z�Ѱ~)տ�'�L�I(�&M ���Ll����\��#6H++�އ�6Re}^�2�lyE��6�q�Ͽ ²gg6�H)N������S����̵�3�(|A�/���yX���B���І4_A��G��(/O�'4���I��m�<2mΑA6�w>L�4k|h8��
�m \��
_]n.�]s�]Uo,s?���1�V���Ó�����Fo�.�-��K�߾�b�@-m�X���2ҍ�Z���(�[8$n˹�;{;��wʡ��\�����_�El\tъ�Q�*��]h״<;"%�z�1�E�290�G<�@���>��GvQO����JZ�_p*�hwZ:�<�)p��ep073Җ�����R��=Y/ۓg�귛�
����mb]�>q�	򝶕{]nׯ/������|��u�-,��Gk;��m��M7����ն�����������۶�f��l;�C�����l���rH䈛�S����p@�ۧ3�,E��(d����U�q�T�i����#�=i��u"�p�eW����#'�-!�����r����؇��8r����_]���#
n~ʱ��%NJ��#��ta�{Tٽ7��Cx=wq%����,a�G��O���Cz���������T%����F�#��u-�ц������RwB�ߚ���M{��a<:Y
++8����P���2	�#�Q�� �1#a,|�4(y�X����#Tb�q���isssmfv'k�-,�g����T�{�L���
F�B���� �y��D��sxx�����8�av`���r^V�dY����������a�.��/��0�v�����)���c{��������N�WS-�^���r �Y!� �{���8��G'Ke���j�3�%]Yh7o��'r���x�d�W�a	
Q�^��I�YV'��q�,KZ��Q�\GY4� �;�_�p��q��lmo���:aA�6���6ζ�:��#�Tۚ]KO�|!|-S�N�[�A*���[�y	X��B)-��U�q*d��ʯ�?���I�2�?�^�(�j��y�WZ)�̑��:�"g��"�@��ҽ2�$����\>+�ѿϧI[�+^�����?��*#������;�m��e�r�*�G�B^���[�������Z�ԩ�B�C���QF
�Α&��l����S�Dr�M�WJ�o��y	��B:p?8')۳���9d������<N֛�y�.���s�m5/�OC�;뫧�a�蹖򺣅�O!�]����xX�幯�z��J�*iCZU��J�Q�*09���*C�8YWp�ZV7݇s�צǆ���L{p��ս�!Fǭ���t���6מ��5�M~������0^��Q�x4��!.�ŗ1�,��'��o�;Q��=�)��`���i+�7p�����t�J�F�/3*�����?�@�pޏ(0��-��������a?7������e�E�,J�'kGtow����F���z���2�Sշɀs����C�?s�/�6Fϒ?�
�.2_���Je��q�	#�Pf��	L�G��Gz<3����!u������<g�O�1��\�����Sag�E��AK�1$)���[�"�)g��3�z6��ॢ�N�9+��|γd�<s-l�%|��o���٘G9qE�F>�i�.�!�A�n�����)7��Yh7n�h�+Kmz�Ց!!�l�."uqͻ0��y�:#~���v{�4�E��_ߋ�з�����,hΡ�q�H�!f:X�3�4.=���oѡ�:��;�I��(�y
��Gգ2|�mh����L������p+� �VDᔲ[nғz������{a�^�hWȻ�4Ӯ_�Ŏ���v-�����ܵެQf�?�Z�%z�zT�kew�0�C��������v���69Y���e�/_��O�e���y�NX'�ݶ���ސ��'/�+�wΟ6XqI��
�q����D��nmne���o��֠N�t�E�|��-mWo�4CY��8g��4"����~t.���a��t�r����ԑx�:Y"�7�zȺ�z�	�0z����{�&�ôr]q��J�Ay.%��}��0�X]~���u�p^+w
�gǅ�|Օ�ţ.h��Pl�N^$+��ޕG���K\{����.�-/eN����r���� ��,	�9YU}�;�:�C'˞�=YY��L���!ˇ<�bTv�"�HЮ8�ޘ�9AaN��ζ�k������Ν;����a���m�"�س"_[haQ��F���jp+��՗�a��ɩ���c��Q[뜬�P���c�]���B�L�sw���R9�N���(�b-��0�X���Į��NA�١6v_��	�X⍃e 1˧c�3���LbT�����ztą;�O!�������:�
\㉻c���{���$��\�u��d^K)x�Ñ�Q���j�,,�Lk(l�r��c�w��;6�Ǝ���ĉט
��܉8�u� ��R
_aRuܯ�gK�m�}S�hW{�K�۴�H�:����6?������nϝ�8o*F�8���
uoѡ�~�}�ܣ�#뱞z�B�_�{�}��Y�i`6���8<����Ҩ��Jz}��!L���g�����Σ��8���r��U�*�t�_���3f��jA�-�ٺ���6�w�bq�<*���h7��j���krr*�;�̕��6�a$�;����٫o5s�Tj�K��p�PyR#����q���� u%L5t��]�F�KC���o��(^�,2*���]�%i�+�J�toT�'/�p�*��:pX��#e�.�=ʤ�ٙ�v�Ƶ��������������ᶻ�6޾H��^�s8�l�(��r*`J��[Ɠ���:ᷔ��!�|����}�l�E��Q���J�u�~�y�N����&��,�!5JJ:[҅���W-����5��wਣ�1?9w�;th���K?M�>��@��{���2�y���l��lOO-�`̒�^� ����)ԓ^�no������<�K�-��%O��^���4�l��=i N�WΗ���x��%w5&L�Q�H�1x���#b,�P��r{]4��9v3W���r�2ײ���<�B,�=z�����񧾗�!��������U��,��/y�!�u�k)Q�U�	C�42���r���/K��+��J޲�R�}j����۵��v�j�p��
��T,�LS�y�wǬ�$οrć�nh�[n����+���B.��{�\��F
��"m2�lϊK�O�;j�вϑH霬���ˏ��W+L�G��w��F�>W�e�[qD%�0��xn}�	��:%w�Aҭ�5��e�ی?�pk�m|d��\Yh�ݿ�n��n�H����w޵׫k��Ы׫mk�&l\���/���^kYpIU��;??��.>�����C�LO����>{��}������~�>���\�̽y��^�X}���������g���B2�L�%�遏����PLm�͍���v-���4� ��8*{RY  ���.��Ζ�$M�th)v�r�84��Y���d9-�߾�t��AS�)Ik�3��K�LG�v*�G���m��(�5��w�So���z�wҜ��}C�z�2RV����|,��
����uo歟=�x6~]go��O�4t�k��̕8�Ʀ���$e.�$NMM��E����4P�e������7q��ɺ��%�+]�C㵜,��ʳ�Ri�Z]4uVaR�T�b���w�V��mEs1[��F��{r��J��|�������ￇ�u;s�l�qe�����x�z���"��M8���P�rX��/��}���[��Փ�;���ɲbS������=�Y�*�{��/=��-�y�F��"��[�Z�ߎqDt����"�r�������:˽�W�\"�Q�W�d9FFp
�%uuF{�n�Z���o�Ӷ�4Q����q7b�,&A�*S��Ki���7�C�F.ZB�Tv�P�&-�T\1'sPF{�(��	�\5t�-����M�x���g�#�0�qpB��އ$���Z%m��+����"|M�\c�QaC餂�0��3d0f
0R�a�`H}���C@����֑���]�7i�g�%0{AR��7
�|h�y�����в�P�_�p��d���{��'�Q�Nw���]Ѫ��}����pcN�Q�yt�OP:Q:�*deS	i�,��[�/�z�T-ڜQǝ"O~Č�E�������ܮ]��t-=Yʌ���8W:Y�.�V�p�r$�sFb�R�4>���2��9��a�c��RI�tʀ�Sq,�4��>��/��ߩz,�����`}#=]���v	�^�X���|��~��X^�iw�\o���A����v��R�nG������u��q�Ͻ�%Li%'�6_6�侜+a����rO'��I���ׄ7uI\W�u��k�n�۷`��l��yWH+y��a�����܋�2�.�����x�M>�����|hy�w�_W
UK$�:�J���y.l�����z��ˏkЋ7�)xS���'�,b���>�;�-)s�6^��W�����m�PG�hUs����~6�F���t?��z�L���*���da�ka0F��3 ��@��]���<���|���(ꎺ������	^��]JY٠>r��/b����>Cf5�5�I���t�|�*1x->�y@
��OҪΕ{f���Vf�3�3"���q�t��9���H�e��/�M���ޝ����m�kG�u���*mY��i�6�j^�s��k=�K�KGZ��%	#��1��܊��*���l���	��<�8�~nv{����l��\�9���F'kd� �q8�˷g� 8����0�qd�84_(*�g�Vo�2
�R�6ʸ�f�(�F���|K�q��|�ûw�������G�mwn/Q�Ql>y�E�޵շ�?k���aV/��`i1C�a�/�����N۵8X.vq��u��j�Z.���׿��oۯ�E���q��ֶ�+{���nO�hϞ�h����u��������s��g��!޽ko�����<saI0�����q& ����kB�(:��8�o���m�n�7�'��8X*��֬.u"����Gw��v;v����g���x+�BxWSv�p����������{���఻>8�o,!+\��/�LG��^��xѕE�AM�Ƭ�G�
�t�;dj9���`"7M7��"i�Y�t�����_SS�`��K�5�D|���t��o����㟯m���'ˍ���txR��*�r\�4qj�|���dQ�)|K)J{���8Y|�0���Y����{Ri��֭���?|�>��8X�o���|������S麘A�0
a�KGE'�q��5�+W�DRz�`,';��8s�6_|k��uQ

	Ɋ)����H]<4��<�W���+�}p��t���<������@���!�R�QN���"0�KN.5#.s��Ͱ�}�5����[�Gp��������҂31^��Wi��ތ�e}�9�eS�^e��̥�þ�r��Qf�P�p��?�`9��0��)���eƓ��w>C-�f}����PT*b���%tq"1���k�U?���: V��O��g�Ԩ�U���<*i[\z'��3�9��:���M��SWݵ��>��uPS��>!�6�`Y=G8����GZ��Σ��D��^�6��������Q�ї໹�q��y�Ο^L!y{�k��k����MZ�{u����^p��1X��K�2*�){P�{�Ϝ�B%��qX�4����;�歛��r8��nm�U�^�_���F[5{�GmZj�;q�G�C�P�D�i��⺌���� s2�
z���V��(��zP�����"�A��@��	�8�:����8w~�<=��07�޿�>��a���G�6�Cɶ7Wۓ�?oϟ}�6�_��mү���!����9�$Ō,5��O8Q��YI��\��y�jT�'������]s�������ͻmhv�! �{坎�r�Ƣ�>��%��Sݳ�W��idC�g]�G�2�N�}d���w�5�g�E�q�:���#=�"77�Ӄ��eA��9I*�>�Kq�y��������Q���m�NO|�=�,~��2��pF�۰ku9|���j�l�K��|.~u^t�Mҳ�.�vA	<�ʅ�\����{�x�#Q0��u���,��x���-����b�Y�R�' ��<�bwu?��7o���J�+��X�ZuȄ���������^!�6`��}���	z�����h� NM������`=�w�ݺy=Ñ�|X~ձrΧC�v�-.�F)�8�G��^N����@��n�\���^.��Y#W'K�*āCL����+��+������<M�zw�TדU_��\�����h���ɄC��<S��^9˼��#��q�8��J��ߓ=)��HSiVN�.��`{����G?�~��ѝ�^,G m휴7o�ۋW�	o���΃<��$���9����z�`�6�s��߻�>���������݄]�W����q���~�>���W8X�_��lɵ�����6��]��X�Fg�=�t\�#ĥzK{�e����ً��8���8WS��W��Ûvv9`6�"[�N�8�'�<��}���V}�V/6�=��nP/��v}Y�߅�5���gfQ�Us��$=�Q��M�ݎ@��F��z�����ݮ@�˕*�nʍ����u�{N՞q8�Ќ��RiDH�m��q"�$?�G�$�������^�+�����\x���tI9�^'k�MR��ԍ��,:YK��r��o�������N�������j{������C�
�HT)k�8�E�.Sd3E�*H��
$���Χ ��5���dO;���|�>����o�Źئ&��
Yt��	ht�`� Ą�q��0�N�����@~��8�c��!�`����y
��=����ȫ?7�si[ӑp�0�S�!�W���=��j̟Jݡf `��%N��v�\&��]�����+�ѡ���d���S[�e�#� ��� ��Ȑ �`�S.+P���D�f�i�#��%E\'�:6|nv�-/L�����ʂ+�4j#`� �sZ2Gjߍ�w)�L�7{����c���a�n꧟��~|��7@:R�p!�+��Y�ԣ�ﻙ[�4��iQ�R��g���l�(�U�7�%a@P��z����!ޓ�-�A1�+=H/�FQ:�����Xķۼ_L��/춘��(o����u2�%F �*��sA�@ �H��g	۸�����ѥ�OH�e�eUyK�
]Yn��)��4�&F�߼;��e����֦�ֳа[5H�|#FM��]��
<s�Kñ���?ҷt�'�[�JS0��z���>��!�}�{���,r�-���������@A�'G;(BWd�S��,�L��z:r��<� p���s	�("�R�rp���r�Z�v�z�{'����rh"09�kc�m[}���
�x#2P|Z�����']�@��]�;�9���/⤹[��-v֡)@1\��3�O�+����ԣ�L6j�`r�!����<ql�C$U�6<��eㄼ��C��k��A�>�k�����mj�J���|�~�����r�y���_�W/�h/��v�ހ��ل���C�.�˧���U�c�&Z�8y��,�T���hx���GENyE���6�t�-^��fo�+�8X�����&�.jMMX��B^����;���}ܳ?�(��,T2�s�2�2POq*S.y�t������i(?�+[���ڛ���5�|�|��CJ<��~��R�=G6����ꪄ���Z�O燺T���ϓ2���=�����b��ha�wI��Kȑ��T��%�խ���!+m�;T_����D����[�Bc���%
-���++�|��#oFVBG.�}�������:��5��m:���+K���һ2[�~��uJ�p@�ܓDc���.G��|Q6���%�;�q{�߹iهcJ#١�n'��ܦm�Eo�O'�h��\]A��id�2����70"g��4F%J6�S�ݝ-�񚋣�������ai#��Vlw��Oe]Ki�q~jQ�
�-u�\�G�O�A��	�R;�9Y6��&�rx�+=�`��1��"��������HV����t$Я��"h��%%yJz�P_���$�l�s|����_ŧ�h��A6)�q;O^���1�����o��O���9�x��/;ck��j�}��I�����󗯰at(+<��{�A����	}��nAW1�gڍk�miq���+C�:I����ן�����k_}�U�o�А�.�_Y.n2��:�	�a�ù���q=EG����yt���i�ܲ1���O����E{��Y����Y�H��X�VؠDg/�w���.GO[��TF�Q���
5�]Ɔ \��^�ؔ�
�=ϕ	֓��|Ĩi@[�R{��/�q�6)����0U{�t�fgfq���`�RީI�q�I�)�'�i��^�U6����B[Xp���8�9O�*࠿k$��Ex)���>p#	��~K�G���P8Ծ���9�.v�6��U�#}'=�ث����6
�Y�݆�q�uaq�-��R�ԙvK���s<�H�Bb����i�ɳ�Ew��7��@�I�����d1{�ڵ̿�}�V[���Dx�5�it��޿K+�Q �b@ky�*D�aK6�\��\5�dh	���P����A�ٌ�,��a��F�Z���g�9_䩷����I�����D"J�Bڐ�`����<����X<�F\X�"��3�l�x��r��u`׬+�)�&�΋�j|{�4XA�}=���%hT���+�S���R�[�� Ͻ,\��lA��jG�&�~A�ZK�1���w�f�N�o���0L;<F �ah`hd%�3�RM��k�4�Ʌ�ըD	����0�������L&߸q�ݼqa�0�������$�T��B����:p1[�%мP<O��V�cH�T���QO���M��J����ӫ�J��xT~�T�(�J}wF�u�9�(����I:��C:��EY�Yס��������O�_�;H��G�T��gw�ٲrT�H��)Ћ'
��B/���UWʁ::xs٧	F���O��௎QK  ��IDATq�������9�!=)о�6Px����'/�sA=�'\*W*AQ��0�#���K�o�J�+���_�_�N�u������ѹ�$	{���gpNf/Pkk�4�o\_n?��G�������>�8\����o^�Ǐ�lϞ}�^�z�ܼ�Eq�/�{����F�Ȳr�Ļ�MCI'�sHǑ�.�i�ȋ�j���U����
���g=��ѡ�p����A�O<z���u�N�t��Nŋ�p�B�Uݞi�9�3`��K�+^��J[�&�x���s(��<�V0�ҁ֑gt�<fKq𭑏㤣�#��!v����b��L�`D�a�G4�m��'�=�� ��GS�ˆ{J�w{��S��l-w���~D�)K~HK��V)Oz����ܓ/(�F����8K�g��g��k���ғ�G2d24�&��zIk������= Ҥ "@ݿ��G��s�c�	{�@�.�)�r�\����R#?�0���v�`gSa���
���l�]�`!��5��mnm��I�l�{�W7���@��^�v����ZYY�^gӞB饓�!9�ݹ��y�
�H�q��FGkc�;L���:_�K���f�{�|�=g%�.}�um�;T6#Η�ޫ����\��c�л�q�z��=�y����b���ɋ�S�K�!����}�ױg�V(�ڐe�8I�6W(��{/�3��>�9�1}�v���/�W_|�~��_��_}�޼|�a�o߬��_?i���/�8X���͡���<�o�Cߛ#L�C�u�\�g�O%��cgOF�z=?̽����a�>�M�:�i�{�,��������k~��v��݄{�������������Ç���k�=j|�a�>�3��O��˞Y�FޒW��ءx����\kd@J��`|����Gw��:{������D� �r�q�#���}G�yB)<C�ﯻ�2�w�O���A9�D,�{��.� ��� N�@�0ƻ�*~��F������z��~�[�]gE=�!��S24�zNH	�ჯ��%pbLq.��=#�W�_]x~��{����F��Z%U<]�줗]��C%d+cة?*=8	��ĳ�gT���|8�a)���+��r����5�ff��s��e}��ιr	�,^��ϙ�ٕt�)��u���.��c�mɩ���P`�5r�����5>�B��T�k�Γ�qȂp���Fo�څ�(��Ͱ��)�/�_����5lzj"�7����7u��q}�-..�U���v���Ί]��t�ۊ�9��u&AU�����'���w!Zν��M��>E'���E��G�q��^'8�dn!Fk`x���h��O��i�[��Sldqx!t嬣������q�:��}�}2�縘RN�,�'��r�\��[|��S/�z�v��{��o���š�]9V�V�Wŵ`,�Rm~��w����a��4n��@~���P��T�9L�t*�����׽��ɕ��}Ց2�{��r�6B�ۋ�l���ÚN0N���P�ym���{��I���ғmw�={�M{��q{��yV8s2:�u��0u@�!��Y�p5b�)6��W�FN9�ԝ��BpXߦ���Ajc�Ζ���l�B�xK�U��������'�Ԏٳ2Vƃ�0C��WO�U߅[��*c|i����!n~���^q���:�]y���R�)ߜ����ur�Õ�p�O��ĕ6?;ܖ�sF����$w��K;m��u}�^ҫ���a`��:��N�y����s"<��Jv����x�oF��ݢ�G}g�=,:���r�Ꝇ}�xw<�ϙ�F���q8���#��i�*�����ޥ�+�N�b<e��>u��k�:.�a^�п�ח�w>��"L��g���>a'?1�pQ狺���ˋ�p�zI��=:`摡\8\��^qb�b>4�,)�i���D���9`�-/���3�mn���>�FOCӼ��g<���W΃_��L0	�se�{y��:4��R�l���钏
b@y���u{��y{������r&#f��딅�32�P4.��e�|B�D��|0��2�.�@�f�f��{H>�ۛmok-[W����AF&�|�5���o���g�|Ӟ?yڞp��_}���'�~���o/��	����G�>���j�>��S?%��u���5���W�wP� J.�Iq��?NZ�Ƿ�	P	6jHS�S�ɚ�^\Z������k�K�������|�`���8d7��[�۝�w8�"�u�ԅ؂�f�*���ὡ�w=΋s�,$������;����{�p𤻪ԍc�������z�~��;`����K�ڣc<oJ���┡��RƵ�`r
~�%���9@Gmw��lM��D�8��U�*�����"��`(h�C�Q�;�@�J��Q~ϑ�F�@�i����}������O��ud=<>�[	9
��\�0��0C�K��++��W��1�=+b�wΖ��B=�#��4����<O�k�s:8-���G�dY_{����1q3�ԡ�qf QWq��/��k�x��Pt������ᄇG:\Ё��0:q�}8F�c�j�w�t��ҭl�;��"'�-��k�
M0 �����U)�PX
{{*������`yi�]��Ԯ����ׯ,g� ���V�@q^��&h�H�UO���t������On�V��w�zZu�h]��@֦��g��E�eZ���`�� �� �pq��Sh$��fSL��P�^��z]W�T���V9{(��8����ws�+~���4~�A�<{n�����4N:'˂p�q��>~S
F��ܣ+�?���ʕ��߬G�q{#"t�@}��p��7��qE���eJ,�/��M�G*�+��sz␼���{B�MՕC-mX�¡���\����� q1����63>���Xj?����'�{����m�����o?�e{��EsOB�29���iނN|Rx������+�˞��Û��ݛ��ˡ����Иc�2������>3� �<����G��s��9�`��;��v9gì�-�ĸO}[���PC*y&�ro�bV�!n9Z�)��~흭�QW_���+��?�mV s���췑�c�� ��H��,��Ļ6>�߆�l�hm�G��'����0���ڑ� `��ܐ�a�P������V�-��1���������.�$���O�W���rړ>����s�흢��� �'�^|}^'����[匽������9D�к��+q��b\iܴ��8�䥬�!�]d
y�E�8����z{��M�����A����ٳ��9�=�ܫ4=z�-,�ht*"O�+t@]�ц4fɂ����{�І$�)C�=��f�p���Z��Y�e� �T9PU@y�OL+�T�~.��
��_��7�pj;��l��������}�Ǘ~C}�H,r��AD�i;�Ό�_��]�Uv&�v���Oo�\k�<��}��G�����+�<���K.���?�gz��d:�E�\��k��7���~�>����/��ӿ����_��z����t�n����.�<Fd����;�O���a5F����o�^+D�s|+���z{���W���	�F���e�S��@��s�i9w�*2�iZ�yա��{�lyy%Ι{�:�K^�.���3]B�)B_�oݟ?���<�gޝ]wR�*��}���D�Tc�6DQ��9�0g pCw�<������@��,�)�M��  +���MѼ<�w�c�l��c�y�Se͛U��|�.p���o
��r�7�obl���IPEd$Ev%	,<�����*Y]!�����#�@�����yũO��a�}	iI�*B�D�Ԫ�!o����0z>��R�A'�W�+?�[r�#a ��--ε��Y��eD�o�u����ب=_86�j'?^T��w8M5+�r��B��N��U�r��h���=-N ���r�^*�5��q��r���q��ګ3fD9YYT���vL�@zv����^`�1�C�ܝ��Ѵ�/���l���ZY^û�͙�G:�r1��R�g�WD��Q���{ƭ��PyE�r��H�g�^'D�`�\jD��( O�Ϡ
��Ī!���+φ��{��Y	Ǽ��X���밸:5����C��[G=������۳x�:{���LЉ�3䝟�'pa]��4�xf�m�բ'㓏<F��/3���4ĵ��������p�J�@y�E���М��[y�t�7]=��yU�c��'{ڪo�t�<�
~Vg�+>JK:V=�:�UGܐ�	�j���z�oې�����βK��6=v�ݻ��~�������v��
�~{�����i/�~ն7ޒ�XBc�W-˫Ѥ1�A��, ��SҊ��3_��@R�0ro�5��	�rB�8iı��{rl��0���_�ly�<�b.<�O~��j�+���Fb|�О~���k�*۸OUN�t�����3��Z"�ԥ%"���c� t���!�tHÿ��Q
�S�>��Řj��6��ۆ���� 2t�][i+�m~�y.ȡ����ެ#�y�G띛VP�#���z6_g����B,���|�3{�Q^c�ϲE�AO�)r�2hL��׹��}_��JkҤ�Q8���^��|..Iב�GZ�����U�ڋ�"m2���1꡼��Աꇋ�ӄ5��0��;�E��ip�|K�n'�ffo�:����C�Mҏ��`mmm�����}�ʶ��J+eg��3��}�����.��1n)���!NB?��|�cJ�� �K��sq'��7�X2�4����+�?L�g��b����e�����#�8I66&RlSe6�[SZ���q?" i�bw��mn�dናC��F́6;1�޻{���?����W���o��i��Oq��;7��g���T[�ž�!�fo���Y��q�^={���o����/���o��Op�>kO?n�8`�a*���8ʌ�3eP_�w�H�wqz:NiR^�oz=�ԃ��/��r.8s�I�v�|w�'�I�]gx�FpԢ"��p(�C	�z2>�*���a�5��8luzF�L�nq��¢�2gK�LG˵z�B]Z�'�Ͳ[�<���g}	z����u��>���(�y�?z�Hz�=�y_�H|h�$�?r�D�~��vHN-p��*x1K �y�s����R���z�!�d}FW�|����ŋ���_�/���}��Y�km�홠[B�1��Q�rD�L�aշ�b�� ��a�
��<}0��B]_����w}�쨸|CeD��g��s�ҋeK�p���W�Y�u�
VhZS�y�ޏn������Q��Ί�S����s�Ĺ�-^�w�k�,,���t�pXA�F�C��QYxC%��Z�%H��Bޡ����;����J�[�s�����B{���&�cEPqV����� ����`šw�U�,m�:��!'�祌���g�'a�0�=h:r1n"�J�i0�Z�B�]G��L����l���;t ���=qI�:�g�Pk ���,��x�2F����y�cp!��v�`OF�mnG�˵�rt�H'�V�M6�L�MmX��<OPQ��B������u|�U]��//�	GpByK��CW�#k�{ST	kxh@����C�w�-}�x{L4*��K��)5��V��9:��1NW��j���O�:����(�#FO��x��Ψ�1���֐gߺ�_KD��-f�u�B8W�8"W]���e��h� �?���Zj���}���v��|��!��ɗ���~�^>���WK�0�@�cF:M�k�`��K%��T9S�4�^a5�|v�SM��-q5�jX��W;�?x���>$�!eE�B�Z%�:��O|�E,u�з�z��㪬�+�JZ��F����Y���Y�|␆���?rdx4�}�Iܵ�`��8d��u��!߇�r�:��C'Λfz�c��>u�<���#.���~�׆����@[�k7�'ۍ��8}�M�n/���#�q���G�h(�	p��-?� �hJ�X��r�8xn�A��u�8���X9��8�UWד�vV@��.T�F���w���T�2�?w��(�"�����4����)Ⱦ,=��ųj���@pVʫh	Gpo���
��l^���Qx��d�mi�$p���}B��!� Y_�4�0=�R���'�VtEE8��LU�׎x �UU�i����IO�J���!��Źn�/���wR�Ѳu�Ǫ|D����_�����:q�lr�z�H!72�	�F����K���AK�!}��o�����/��#�|��K�w�Se�N�i��q���꛵���F�ElA���cK�3��of����������������O����>m�'?j�����G�k�~�}��G��=j�?�ۖq�\�����~�����i{��)up�E;K]f�H��dѡ�[���l�N�t20��B}��g���r�q=���<�_p"��+a#�}��Q�t������O���D�"]���[�6�CrO0]�%�5~��e�@	׷`��ɸ{��u8�v�s�Y�V�ӽ㿇�[�.:_I?y�i�#nF�����UF/�F&~!�[�|�,�F�Jd����$.
i��M�SX{Wm��}�����8.K
�l�L
>[]C�Ϟ�h_|�e�����o�s�d���PW�qxL�� �;qc1�v�t�僃Kmg봭�ﷷ�G�}���{��zZ�֏{=.8"�w��!�}�>ɕr����!+ZUV�*XQŏi�C��}w�v��վl�V�/��Ͻ y�[-_�.O웟q�V~S�U�ۃ5;�P��v���5Wtq�x>WԏHӐ��s}���r�Α�cڕ��y>��]F�G��A��j(1pZnߞg�:M�snL�W `�����-*�K������S�>:Qm˧�X�.ء�S�j!��3<�?�&C�:\���q��L]}H��Ri������/��,��	��{�[Z��H�<�I��&�B��@�r�i��	�.��^�<��-��X��C?��%�Ic��.MV�H:q���L��+�NM��sh�? .����/��h~�)��{q�S��k�Y���a���*����
��K�vNwG�������,َ���BYP�bS2�<t�/�a0�r�/��a&���!���&�n^����Vp�V\��@hB)J���"��[�/��;���G�ٯ�f*�x_�m�Oz&S���8R:oY���Ҹ���8��^^=m�s��n>��ngq���`g�=�
W_gn�eh�ޯ8��G�t4x��>�#��Q� _���`�KE?�z(�}��z��\Q'�\#�Wfs��<osKmnq�ML�a���> ���Ի��3��_��]�#G>�'}D�_uPG�c=� ��`y)��t ����[W�|�����0YW6F���#
�!U� A�ø��儕f�҇�c�:��l�t�HXR1�	h���@*�9�B�L�>��G��hR���Q��u����l"gz��N��[�qP6i^��؅x�**��{�{y�V�T�����&q��>���m��T��i�}�����@!�����/��$�-g"��v�:�����C%~kq���q�Qh�፵|���l�����|?:t������$:h�*L�q��i?r�a�
.n�C�t	��%R����_�[:h���.�e��C�w�&��.������Q�F�=�S����4�s2>��e�yǩ�IvaС��ş���`�� �r��<S沭J�	������܌��se]�(��Qp']�g�az�f-��l���������������8�M݌�9��͡���76�g�.�C�^r�iז��nj�d��AJ8En%1��S�v����g�����dA�͛7��"S�N�y�c�z��\hZ�+�{%�:?\�J/x&�sz�v|����x���6���<���րϺ�/d�|�p�����t�?�#��!Sڕ'�Q����hk:�CȜ<h?���-][��k h�9�Ÿڂ:��DH�Om�M��Z{c��j��N�����#a.�L���r���|^W�:;��a������Ш�V�[]�}�0�ځ7,�U�ːǹ�Y�:�^�A'�}�@��lF�% :XCh[��pV8�p��lD���Q
YN��$	f�C&3�q]K,k�l���m����A�֞�x�s�U����7{�S�D�}�,��M�iK���\�R�Q2�S��يR�G��7*�J;h�ӶIw��v�d�"���*-��+x�l�D3�R�8�X�/Cȇ2K|�����:u�Y�,`��HDc17f�v�'��FG�g�z�`�;�!|f�ʲC��̌-�|)�%� �1���P��q����ش�����;�@p(�l�R����D.SGؠ>a������3߅:,��4��L�xJ�g+l��7�Y#[e_\�M�->�ǚ��4�%v���cݜ@�����l�X:@K�c�i��»���u�]���@1U-٣�c�oM+�u�|�g��RB��*ϝ�>d�'��S���{BuDs��.v@ȾdI��6}�K�F��g��(�#jrٗ���|{vܟ��礛�|U��J�UYŇ4,>��ʃ��9 �X#�lB�⯧W�w&�8*����
�c���*?�C����`�q��0]�o�8�A���Cn<b�!�
q�T)�ƪ½Jy�OB=n�n�\Y���#��zh���0U	��Ea��w��\!��ϥ��#C����X�s{�=��ݿ���w�mo�m/�~�^�`9K:t�n��1�O�yE����,g�3�sF���xH%�ux����뱮b�'��#�L8ϼs�R�b��/��9���6BL�ӳ����ٵ���?rt���>�y�Q���� ����}���޼ho^>��z�:���)-_j�(��s�෣�'��E�ޙbe/f9�i>��P�O�f�����</��{�%YZ����4\!W]r?��Iz��R�k�(Q �l�,�@��Y6�%3����q���{�����MW�p%۬f�ux�/���+4�B Oˣs�P�4��O�i�}�t�u/K�D_����*��8Qf�`���Y#Pg���δ���������s����E��760�gj���v�_���n��������Y�Ǩ�j^rL�k��Bw�r� i�lao�Q��6���ԐDt-�t���B]jåN�8��dp`Z�!�1})}K�հ��a��GElp�
�ں
ޕ�r��$}���y�:� ���lD�nC��l=??;�f	�J�Z�$pK�ص�ߴ7o��_���"�ɸ v�B�أuL9�[{T�0��1�o߸֦'Ɛ����-x�e���y�j�]���nݺVj�rǛY����tx'�'Y%�y��ViQ�L?<������(H2���5��,{��)��x'NV��Z}_�6��ԛ����l�O���Jg���#�w�8�А�q�86�P��{�J{љ���{���i��:�2�QWKc;Ю������KAK�_ �Ggvww.\ǶJ�D��U�����O��o��7���S���p.-��u��߼N��=����t	����w�Z�(�j��;�cH�����V��D���og����߷����_���h�W�~��_��p��?�r�����~��������O�>��g���gq�LW��aS(��2�Qy/�N'�+g���+�z�M���G��g��o����
4ԣ��Y�����p��%���$z"-�WH���B�A0�c+CMp�c��a[L���<����,a�zn��gy'[8T�2�-J5g�6�W%��J�Q�{��08�X���n��ؘ-|m�q�{q�"*%��bk�8v��mq����&�Cᄛ`�qc��l��|��r=���5����cp�9Sn�aB���5õ�L�5�������� �{��Io��5!�C�?�(�"S�::��:O�ѡ��mx�E
����e%pm�3ޝ�Ȼbػw��P�y#��r��=Á�hP|J���r�g�\�>{�;�4���ك�u�����9G�SH��=WʚzK�t�iXU+j����}6�����Y_�8.�1k�Ű�	Ұ��`�0N��������0p6$�x9��,ʚ��Ї�0t1��yN��}�I#W~m�H>�r�gu��j�B�^����v��J��f[^��������œ����mk����(��'��#�{[=;z��,�/>4�b�1ҀE�؈�CV���:����򳸡2'�:2�1�#���4�4��y�3�� ���a��*XLXV˅�*Á2Y>B�	�Ӡ������ޗ��Ƌ&퉈|<{_4o�gA���+u�t�\SN_��t,�K���ԓ��.���n�N�-��.W}�:"�	t���Q��1�I�=z�B���x�ۇ܎�b���}�2/g�oT��6���D��Q�X��x�w�_�+�J{儊oeD䃩�7�P��7<�Po��]��]�{_�<��u����O�������49��U���t��m�����0����^��v��}?�toϞ��4���pC�V����Q�;���~��?�U��n
�JI@:��k�ɧ~��]��L�j#$��'�7�W�Cy�h���������D�
�6�U�_j�[��ŋ�훯�`��>�]�aY�:��hp���m :�i˔���p����K�A%�q|�/GR�]�N������'�M���ա�6==ږWfڭ�������r�ug	gk�ݹ{�=��������/�տh��_���G?�4+�@X����:�Y܁�_iH#�sr�g�������Tw��>�/�����τ�4����+]��J�\'�P���S�<�AEO#!��"4�P�_��4[�b�SO�~�+�ځ<��j=���y�-��U������+��(��L5\�:3�#@Aa|h;�S���G=�8�:��[��J� 9{�kE(������wB��t�:O�<i?����Op�~�ӿ�\,W]Q����N�W_}پ��ӧO"�$|��������n�&^@�Y\�?AL�_��x�?���?R�� �۳G�Q8���aB�J�^J%!�LH|�q��
2��U9T5T�k��D`Kl�3ӵ*)�Ҫ�2H�΀.�'/��,�3�^�%-��n���d~��'tε�Q9Zn>�ӕ�)�Bd�+��
p\�!��ؽ�Ʋ���Ɏ�hA:�2�-_*%����KY�'��z��1a }�w�X��ťᑆ�.J+='sh��)�\���2��n�q�JQ�4�Cj��3��2�+����y��$x���Q��sH3u�NU�����hg�,W���_�:8W���*���-?�(U�a;�!��.w����:ZM�ђ�o@'y	GWS� �\���?����3o��;�vߜ�w�*�k�dG�V��ay�dN��-�Ơ�UFU	FC����C'1�1bl)��֡9Ҍ�.�d8��yo�i��徇'�s׽�V���~0v��"~gw��~ήy�4�g�yD _	���
RM/�-j����n�911��nn�XnK����/���8WY�g�Mݝ������m}m��{5�
�1V�Ȗq��'��8��L=���l]�]�oz��-Gp�s�Hk�uC]X�>d�±Û���?p�&�J��?~�S�]<��n�ҊSxW��xsNH� �'=ÿ08q��\���"#8g1R�vN�>��v��S�6D�@��h���x��q�+�:�:_�2��x*�GHW��lVŕ��y��NG����cm��1B��0do�=��^�,tQZ�q�<2?��O�ٖ��s�v�g�� ���hO�M|�7�З84�Wt^<�<�	$�
^W����o*Q���z���K�u"��&'�S��#eo���8Aoq��oެ�i�oW�_���{���3e]���2����M�=�E;�w�N����ϒ�����ܛ7�q��#i�7N�Y#x�ui�W2G�O�N��%.��(��{gͣo6bh��)N�+W�4��VE�%<,������;��l�w=��obc�dy���1�wΕ� {���rE���Oфܛ�/�G��gO_�����h�"�
�5_�{M���ȩ�Xx��3��̌�����?p.׿��������6x���mV�s�A�J����h�	�{{�����u���;��C���9�}]�~)��G��c�#��~���`��n�yN�wI�<f�.���(�M���-���>iro>U����~��K<�Ì���L�<W�zt�(�����j���"�Eɑ�o�;�W�����d���oڳ�x��(Q���S�ӟ/����0�]�� ���F��X� �T(�L�;�TeQ�*dg&'��k���۷ۭ7�˹��:�g��P�����!��v��F�9,le��ԯ����s�r��;�#d��q��S���V�+m��r��=ikۻ���y9\||���� ��h&ҳ�՚��<�q�H��ڸ�����Ec�V�Be��^�V:k�����^	������
��dB���r�%�V���H"Tq���Jf�VG��C����̕693�&'Q�CmE8b}�.�<�^����_�o7W�/���f�x/�>L�Cm �j��\�}dĽ�t���U�hZ� Y�=/2���w��e9dg;�l�?�\
ŉ���[�l��'{������%m0������̼�h</:=v�BU�+8fەg~��>"/���c`'�ԫ�):!�&� �:
c�������s�B8u�AC/^k5�4�)}��E����X٥�>5�D�N�b��;Zk�����:��?�B�j'o����v���yh�I�mAR��_±2=w}��Ѧ�*8��S{s4��������{�%�d�0I_�	�|ؕ#e�\\*�d�|*����*��8s�W7t�c���z����nR)�T�5y7�=��e�k|�5N5�<q�%�Tr�w�،B���w�������-r�� �g-��=�i�'Y�i5��8�p��	 .q�aX����o���#)I#3�l����LZՁ�q�q�5ih؆��_a�K�^9iC��C0�c5���K{���v��T�{s�-͍�A⮿~՞~�Y{��Y;���D��@�}���P��vLY6Ťe���C�"ژc�[��u��(�����U��������Z��|��Ρ2���m�tq����6;���smy�Pe�6����A���r|w���?z.�Cǵ��מ<2��9������ �O��12������o0�_��v���d���F0ab(jp�H�3�<Dj���Ro�i@��M�8�<��T��hU>)�a��NG��� N�����B��f��ts�?��|/�V} �s�n���G��T�(K�(9Y��x�^]J�c��$8đ���3��'�S��+ī8,;%�!���֗4#��|h���w��ɀ�U7DJ<9�Ά����֑!��!K�3c/-����
����;l"�y���n���S����z����"�۫�/��'�5�G�i{��9��K�l0�HmmnfZ���z�u�vq�Ї������54�I�G���~���V_��/]��Y{��e�X续����S��\ViHǪUw�����Zbޑ�0s��N���!���vZ��8ʝL�'��:%���z�N���=��՝�(�)o��W�)��cGA�NGG���ۣ��o]kS���@칧/_�g/^�յ��k!2�W;��y��}7H�RאS�G�d�@��SZ����>cT��.��ݣ]�2�͛b���XM��1O��gml�kj���ܾ��l��ml��P7�G8M�EJj�W��Ѻ���mbx�{�q?7Z�d�`Y���Q��=K��#�S�j���Cĉ��z�a�3Rv>&�`)_���%v�������U���"Q�Rپ������G���Өm]��T���K.�Ws�6��re�K�cǂ�ֈ5p �s�p��W&�l��^[a���㛄�z�,*=����z����#=��`+�R�rV�Ѿw����㟿�ў>A:'�G ��\Ԙe,@H<N�tIoU�L��ڈ�#�7�Cq��h� +L��J6����������G��[7�go�7�g�I�g=Y��%"����>���ܾٖ0�u��L�R��p��Q|{��o#Z�F��o�̹�ka��'cY��B���R�ܓ4?g]��&S쪎
�k����Uq �<��͛q�}�q9wF� ���>%���$B{�4$i����=SxS⮡B�� q�Ǔ�������0��΍�)��e޵���
h����n�wa�珂F�At�ԹJ�K�OP�8����$hX�ٵ���ر�c�C�kIe�BT�ll���EA)�MT�J%fZ5|��+��&[�;�H�_�UG!	
/[����=o��L�����������#�U���e!S���)��cG���E�Q*����>�ƭ?��z�AU��ސ!�&�Dt�x�NT,YNYZqq*{��kՇ�]`���H_Nh����<-���DM�'�֜�	�x`��2�K�s$J~�fŶ������ן��ԛw��^�(�g�+B���Ojl�ϬCWc�A�޾���pP���|a��}OV��N*�I�4z	�??7߮_w��kY:V'K���g[7ΣT>�C���'"�F�p$���3�R�ֹ������!	YC��T=�[Ґ�X�3H'�.�ʙ�S�A�X�z席,ϴ��W���4
�][[}Ӿ�����Q����9T�H�}ﴫ{j���K�`���0aޫ�䇌$ �2��m�#iE��M�X��T�w��B�_
��)���c�o�힝]h��Kmjv���\|l'�V�˫>�譢t1�������������̷��o6������}�#������M�щ�~���L��Q�д֒���;i�0|����~�(i$X%։?�a]��|[�11�I/���E���a�S�l�P5��1�4�b�P&���=�"��7B���f�ҹ���^(`���H��@,S�}A<�8��f��4M�_|�����N���A�3�~��tȇ�c�S4"�]�/�֙�u	������is��i왾�dO���;��m{�߾��/��gO��gϟ�:�~��,{�:�S�&�ʝ�>Go�
*�W͗�L�Ԫ�S8]�]�Y��^�g���Y�;�F��g���j �a��j�(�T�i�;'��)�w;��P_7%�&��S�� 	�ԙ�?�A��8k��w�he�zUzⅵ���	͗n�vJ�ڛ~|���p�][�m=��>��.��r�	2�������r��W�}����i����6�La �2�vY�����<�p�c,t�����t�Ƿ�8�n�<�ݠ|Mq(N�%�X����[�= J�<8q�$n����g"���L<g�l:�6J�Hi�3r�Ls�|�x�@|T|�}��m/(g�aV	%ZO�JF���H	<�i�jă�Ҹ8��U?����Ȩ���,��|f�]d_���C�lxY�t�|�͵�ohQ�i?UJ��2Wў�Mi��d�װ�4�^Ҷ��.��9Է<M�	L���>�w��q+����5?���H�<���n�����ʼKic������7k[����;YY]��N��S=YT��!��dQQټ/�sntD�y��H��*�U�0ʯ�������8X�[�������`9Ѧ���$�]��<%�Z��Ν��G�ڇ��n߼��g�c��$�֎�Et��t BY�w�p �T�mm�b���������J���J�����L���7`v�ߺ�9�&c��p:s���r�WM����/�%��O�R�ZO<e�\�~$��iAq%�A7~�=	F�p�|6��5�9#�2�iSR�J��^��v�=	K��6�/N������4��t��T`�G0��\07���K�a�,�q	�����/!�[��@��t�lճ����T�w�o���<B��4�u��)q�s�;���+��Q��Z0�#�}7�,=lm!\q���ev(@�i�#�d��"\���՛e��'+5_�iX��b�P���g�Y���W֖A�@Ed˱
]G��ltaE��J��k[K��R:��0�O���tr&�rB���W��p��i�#��fU�<��d��ٳ���қ�G�&��Е�sNfsᬠ�*l�d�d��0e7u?���LR8J���ܡr����Z�R7�R\�pUං�?ǝ[���;w2�cy$CS��鐞�Bb-F��E�EJ۝M�/��j�-U�1Ɣ��!
^�eW��s�/�ʱ*��������<WA^�����Ơ��*�k��ɉ�8Y�Sc�=n;[m��6F��Yn�=�s����������2Na~q�M�/���9��4��B5N6wX�(���S�B���LE�_	N�Ys��
��
�@���Y�@AY� )����� z@'krj��Y@��"�u�}�s_AJ,��'������H-����츐������C~�5?����z���ϑqo����u�q..�=Gfh�iDԆ�Ǒ�B���|5+�e��BE#�� @�e�����C��:��5�����Y�״��)V'�
�z��@@�����u[|�W�^?K�7����o� ���\�jxur����'z��.=�@KT���~�Z�x�x��<v�r_�������<���3����1��M�]�"_��^y�|*G����x�ƍ��������w����r>��V�r�-��#�����Zk�]�j��G��:��^L�p����yL���*y9$�-qw¯�s�d�u+�dQ"�%�+o��칑��1��{��8O,�s�C�Jz�٥-Nu�\N]޷f3�)��ـlϜ${�$�8�Z�O�P�mH����qfz����v��������z������W��g�ګ�o�Q�`�����Wf��p�:�6Rh׺���qv����:�:�=+P��{�m��^�Qz��յM��^F���) �"��S�����c��g�T��D9(?�'AK�e�չ ?%��.��P����=X�0��euA��W|'?nKG����<�C���f��BVe�m�nn�g��k>ˠ��G}����,�Z}P��z�H�|gg7��ʂG9׆%�Cp�/�X��]��������B�?Q������;��X)r�.tV��9V�ٓ�6	q�p�P��1�o��E'k���У��:Y�"nA� ���ꂇ�d)x�0�@e<5�#>�Hл�nA�T��+�\����o�wC@�Ric�mn~�- �K�*�-����K���������}���{x��&1ګU�Jtll$v��C$�����.N�=Y��a���B���Z��]DS�l,6��T8���w�,�r�.]�=N�ۮ�3'F �E'+�"Ε���z�����`	#8Scc�Q��ؓ5���898Y�n�;=���YqX�*n�wը|��uZ�҂�bIK�1��9X:I.y��35צ&p� @�z��KY�ۡ����C��dYo҂t!��2�p�Ә]}�&��a�
]�MM』���(0�"�\�q P�S���bb���5�$�J_�J��Mw���� }ˣ�5yCz0e���`eu�8Z�d�p���杳�����N �o����
��U<]h��t�'���v|���Zg��h���l���A�g@i�\U�Y�ђgm	��H?�Ȋ5T�UD�Y�ɓ.T�rE��S�\l�%���M�g?��x�/��|,����(��+�t��ϴ�0n�5���Ke`�<Wӥ�Y�r.��]��<y�r�--/Ei�H��%j��|���_-�@ha�^"�a&[ 3N5F
iȌ�K�8G��ϪB`��蠇�sɎG|�LqA�A�!���YW��1x}vf,�4LO���Q��vE�m��K��d�v�f�y�n�{�A�o���nsm�u�A�~�n[�q�-�\�67���5�&qp&&�������vw	{�	pOil�ИU�:��!G:YN�W	��T�5&r,�.�ļ���P�5�I���'�!��z��|���o�ߪ�8���󛳫��9���?��z�;RW�u(�.6߶�/��?��%�d�_�S�l�	�kk�6 �^�B����ˁJ������8�m� � �	#�E]ڠP�|��Qd�������� ����F��h�G���r�Fy[J�%����~�m�|�\�����B�4V2�����_�AH}��7�����G(�w�Jc0�t�����9S���a��S9N��d�Cu���2D������-�%|8����ֶq��R�*W��
,��!WԨ��ʅxv��A�"��l/��s�WCU�Q�g�C	��7T=;�/���q�8Y�͉� ��Րf<iў,j���fA��ɲ.JT��<��vUBxT޷�ӻ%��K��M�b�!��a�9�Cp����Gmiq�}��G�~�Q�}s	��洺)N�;8n/_��g�qdq,�w>k���QO;4�a��{�v�sj/�۞��{G�)�Mc�I��e�ņX��\� ���F{��e{�-��|�y�'O]�Ì�%�9,������!�O�������pĩ�=��A�D�¢u����|��t�z^�͵���x�ҡ�9���T+� #w_�����nm��>�w�ߜN>g�� H�\\�$K����m�Z��N`��o�;������������@���ٽ�ԡ�����cx����J��*�����5�3ДUW.QwW�[6��M���/�Ѭ�]�F>��5�m{kFSY����8��{e�p�Îxq�,-J��^���˨ ����ПK��y�|�ƠG�s^#~q�W����"�U��>��]#��H�k����U ?����8�)�%H�1�BE)(A��N�����H�c���;������έ�1ӽ{�H���	��\[_l�o��PQW��:���?h�~�i�����'h����䴡�Qʀ���0M��+H��t��Z�,��͌d�n#���R\Jg&��g��To�;�]5��i�GB�`����R!��R�.����|*�ll�S�=e�A�H���\���d��@w��x��9�л��8�V��,ᱤ�TI�o޽m/_9��
mF�g��J���1k��r[Y^C�C��^��i�\��
�4IKm~vK���� \∕�=w5!	c�+���k���f��jG.GK����alhQ��8��ǐw��Y`�GBe�3�<ذ��[�:G�N�q�7��_�� ɹS(#S[�XS[/��s�L�(��PA��m�W�/�D(F���B{�nb`��
#��3����C�@��������ýsΥkhL� #E1NK�*�Й���.-G=�<�������k/u���v�S���?n�[f\.*)�>K�NQ����Pk��u�2%=e~$\d�
���ǔͫ�FY�C���+'��l{��a����gT]���i_z|���h���5���.�^c`��#��K������">�(3�Iん~m�b`��
�x�@��h���)��5����rj���əv��
F����S:��g�}���矷O��i�䳟``}�>��3.d����ƽ�Ɲm�ֽ�~�N[_��V�60����Z^]k��kT�\/�*܎�����C}r-U�[����^,4HP9T�oi0}�W����~�ԛN7�Y��\*%��U��G�W�#��=��4_ߋVu��>���� ^J�	t�3*p[oQʞ|۞?}�vw6c�L�RhL��MG�UHT(�A��s���m{�(�N���Yf��E��(�$
"�2���^y�x��_��� _��v�p�t]f�	Ƌsd�#Xе��9�F,�+y�4��2��U�#A'�y���oLK#�O3�)V����mr�N*^d���T�2���Ɔ�k-��
p T�[\t��r�0�(WF]���|S"�qQ��ɬ�Rz#�:�]���7��n��P�R�َ�ؙ ���'nL�l�ڬB>^R񦂽����*G��@�R
>�Klܽ��M����J�n݊�+�%��8]��*�F�S=��t>#�4�!O���2�*�]������\NCe�	F��c�Jy�'����F�t`���֙r>�7�9��rmn�Ѣ��Eq��u39y���]o��?���������nz\ݎ���N{����/��4b͓r c2�A,�&yZw�4�`P]PO�6X8��r���Mu{g��e�V�Wov���_�o�}��y���'�믿k�~�=j��wt�#k��\�����早�Et������ft�l���|R�?��<S��������u G������7��z��;���aœ�	��l�OzJg�7ye���������@�H^�NJyQ��F����L���4�����L��5�܅S]�,Gd��|F�4��A8/�65���>I���.C�j��g�P����.��2G�4�=~�Y/��?�l@Ddo�يKO@������p8]��q~�;S��T��y�gy#
�{n�k�MUf/L�p8t��#H>{5nݺپ����'��O�O~������;w�D��7iR/zpD>*$4d Mal�+������9	Y�x�Ĺ�y���A��cB�i�(sW��Qѳ��Nط�@�@��9ժ����
A�Zoa�h�l����n �b�:_�ic^�2ho�D�����£��!�P5�&h�9�l�s3��Q9t�������"^�>��C�[w tv�`��>3%Ĳ��Jg��;]z"�5O��6�����D�Lb�Ȅ=õ�" ��w��z;.FwC]�}�������Ԛ�ݥ����P+���N_�����:?�gx�/0�.�w��������>��4��+�#�s�Q��lx�F��{?����o���;�َh��r�B�tV>GM�\Ew����Y`@$H�!���U��vx��W�8��^7��K�ǽ��Ӱ�� {�UlH$aL+B_�z�� ��(�N3��������g���/\�{�@Wː'e1�`�4�6��D�i��U��R�)�.���F��p���Ԟe����ٶ�*o#e�r�g���/�Y����_��O�Y����	F��{>i�����J�6�H�9OD����R�]��:��Ɩ�
���'?k_�������?k�g��}��?�P���ݸۦ�Q�����y�W�+C�A7�p����/�xy$�jMƔ����!2=�{��c��u�}�K7J3�R��5��4�k�������zB�cܕ$�s�g	�8�{uP��nTaϬ#�pF���!���Z�fo����E���$���<5]�yV�����K��[�F�J����A�D�nzF�
�

�	ak�F�h����U_�H�����1K�<�8Sb��[��ѯN��ڂ�������Jd�i���F��@�W@�2�O;�=>�SD,a�H_ʲ�|cG
�D�K�/Υ��s��HF�z}��S0>��pj�A�y�_�x��R�NR�s�y�����Q�s�J7�ШR	�L'���z�w��ͽ��*���:8OG��>��ݽs���E�2�EN�����g�}�<x�ҷ�r�"�j���[X"i$���Mޑ7�w�/������������5��hم� ��ĳ26�?��p��b����q�����M�n2�L�~C�N=���kcS�Ғ�����C��.^U���t>�|R��1�w�r��+-e����b����L��}�}������������_�����������������_��_������?�M�������w���_�_����髬��S���#�|��]Tc:H�aי:bh�t8��f��b�l�L���3�:�^����s$�s}�����~�8��s?z~x��;x�t���� G`�����q{:8?_�W	�����+aH���t�D���\��~���|�k~��|�8���7�߁*����C�jI֤���@��Nz�xE�w魂pPn�םW��)�Z��;���@�|�*SZ0�>����1�����݀���#S/(fPvG7\�T}����B\�a@��!~���w�";����L��q�n��W9U�ʸr�F)+�Ù�)ϵ�Q��&7���6����Fw{������A�;�L�Rxv�ِ����Fష=�=_UR<��N� �d=���\[vD�85	L���C����Îf9�"�I�y� �h�S���Rݖ_�����A�G�o��އ���i}6��fkd�����e,|�륷�EZ�Qn�����ي�|�#>_���}�ni	IWC��x{�T��%�(�F�`hq�8��;���x׀:�fNU���'�Q��u:^�Ff�~r�iIN=Ҁ=�p�k'VG�\(�x�wch��6�L��)
x��H��.$�k�y��}g G��}��%�C'�E��u	�>u����(�weX�0Z�G�q�����J��O�g9����;�>���pFِ��k��$����5i>�=x�aJ����5�Π�M�P�i1�Z�3����M���m}�5�B>��ݽ����'�����>���v��Cd魶���r�!5�Qum�ܦ����\�8��R���umj�ML/�ə�6��֖�n��?h|����������������'?i�o?hs+�9�r���鄮��ѷ��M�k��
���k�u嗎�1�P�O���)r6r"F�8���2V��l*D�/�z���3ސld��Dж�ȑG�ww�2�(�=����rƆkآtJ#�T��I��\7��l&ah]ww33J/6�����:�҆�S���9��)K��=��}���x'��!��Ea��a�5-�R���#�5��M8ʥ�g�a�ᨘ�+4/��L�R3���5�~R���]Z����/���wNx�(B~!�ܬ��+�B��FEޔ�5��ąy^�T��w��A�]p�_��d�Q��eӶJ�y��w�y������+��{yV�����}
��&Q����df9J�{�WWW1��/>�I��O�����,>]&q���~�����O���O�?F�Z"��ONR6ׄ|��G�#�$G��t@8
�r�i���Swi'�!�Ұ|�O���}�[Е�v��ɰ�A�k,����Z˄���P��A���t4.��^퀂��{G4��t,/�	�W��_�L4�[_D%}�څS=���.R������sR.iE�_�8�0�Q�9��r�b���?�����;�2��΅�=o�}��}����7��7�=o��l/��n�^�m/���־��1��ܭ>j*i�n����m��H��{�CAj{R�4z�5%��uM=���#���������C}ׇ�8���f�f*���u�X����mW���G��y���n`����0�ʋ2�z\���K�n~����gh�|)�%���_��_E�3դ�ϥSׇ*��J'�vڎ�ݰ`Q�$�����6w�~�K�C���E�E��H���I�a ƞ	{�*�\(0 ��ap	K�vbvv�-,��<7(=5Ǔ�G#�F��^X/K5���8{�_���&�J��_���p�UWW��F��K��p/QX����+�W�g�"[ڋA���h�,woqq�S_�̎7���T �;�R����L_e �
�`�F���"���.duFnvv"S�W���r[s+yw9��UN`>�+{j���y��u�X����P�E��Оl¥�R�%l W�BYa {��V�}�;x������R�y�N��A;�C�2�Y:�6��»\�฽���}��:�f]e�F-4.-xp����F��jJ��a�k�z�ϩҡ��k���+0�;X{�o<{*���D8�G��I��X{���1��r������s����%���=�uZ��W���fo}
�Sp�]�y/N�έ�X!N�vM���r�$t�L�]�H �U�G�M�iTy	��n� �f�8&��9��|Y�[\�?\U�35v�d�P�'��S�o����T�a٩�����ܾ�������?i�Sg|�n޺�Luڏ�̐�9 l1��]s;t�������N�h5c3��1�ÏMεY�[^��|�Y�􋟵O?�Y��ӟ���>l�+��t�=�0�:"cy(m�E�(j�ſk���үýB_�u��5�k�4�����H�Z�^C�ý���{��Yu:��7�W��y�����v��溚ׯ^�W/����M�9��q��"��rP�;-�M<P��*���i�hl�r�b��s�3���k�P��Ew��{䛻���-RwKmzn�#z��I����J�dMZ�AhY莏eh��.n��B��������u�2���?o�ZK�mue��)���HY�,�#vӐ��,���R��B��<#VC�x��C��;8qdZ���FW�J>�2�+~$%�,�yM}�4^�ȏ��xc��Y�|7m�f�7ST[-�w��i��ʹ���v������7n�V�e:��S���ǟa���}��O��o�}���:;�S���-��Y�t���:a)�*Á��U�k�����c��bi瑣r�1��"7ĩ�\��F��x:���艄1�餳NE�0���Mg��||d����tf�NC�s䶠u������N�T$��*ߑ(J$�u��0�Qg�ܹ}����������l���ߵ���/�_���]�7n\�n�̗�������}����)��.�x������^���6eK�k�^�p
zm,�	����M�&��;�6�}��?�~�I�����wVԏ��u��{�t"^�G�]���(���΢���i��.5P>�]�h�;Ȼ��v
U{DU�GeQ����@:�0	V�F�(��-=������=цt*v���(�%2�d^�^�"A��q���?�~" ��^ɸz�� �x� �޼��K �Te� 8:�'��ˋh�9d[ʵ�m5@�0!2A2T�4T���l���_gZF�I��O��\�:1дU
��Te@���nc[#/�a��Z��J�-�\k$������/_�gn���Q,�lyM[� �|��H�M�ku�V1u��s�`*��"97;E��D�����]�]g@%kLi���t�߆̺S(J*���{�	��qT���IObK��U�67�p���zvQsZ�iF���U�����a/�
&R1&|MjFqU� |]֩�|�������Rw>Wr�K�+:M���;P���P6�W6�pO�cu����9xַvMY�@�ҘB0�x<��3�v�B4�e������p���=N|�Ph7ց�V�m)�8�i�
� ~v��u��PB��=�|����� �U(;%k3�ŷi�Sʥʭd�J�^:
|�J:�|�0I��N#W��7i:��뛤s�z�m�"|���tF4�'�AGA��_n����.��k���(e���>��ݻw?����ih8�1B�;�i{ns�2=C�����fX)������)�O����9�P�WV���w��~�>����ǟb��E�Z�I��)�("���R���8����h�F����vS��ͷ٩McK%"!�ͫ|8<�}�g9+�z~������|�@^q���P=��흽�*�/^��ܳ�����՛��>bj|ˀ�'�خf���v�-^D-#��+�^�(�!����!�\#�����x�ݺ{?����{H�=h7���v[Z��Z���5UaVq^F�_��(ԞKxf��U�,���[v��	tz���Z�_����!�Xrf�<A<׈h��^�:�Z×���T|�����=�ն>���&,��u���@=D~E�SDܪ�پU�tg�q����J�U���m�Q|� �A��	O�uC����l��&Z*��4�i�-�Nml\o��=h~�郷o�&���
F�<��3|v�n����w�d
�mG6@���
�%��}h���)��e�F��2�6�2��w�,S��yxq��R���z�#TƩ6�v� ���U6ڹ`[��/�ɝ*���;�n�Q������[ګ�?���(�	M.�_���9!���8ӼR����,;nΠ;r<
�f���������������m�����������?i�}�i[[_K�dǬ#�v\8j�R
0������*hW��Q���6��m����k�k�_�E����0��C]�R\������G~^G��v�!.�������xޙ�pJ;�.��W��kD�f6]��U�M���s�r_��:��OG���R���_k�K<_�0��QG��O��*x/H\� ]z-We�i���m�A��2jNÎ�O�����˷���p�}KLj�FO��a��k��1,M��C�A�*�I����L%�1��"�*�;L�s:�J�1\�PU��BI
Xw�����!�����E;T���ʤys��%��|���a�WzC T�������nӝ�.���y���18����?e��P2ˎ�^�^��m=��*?��ZeTyBl���x��l�nO�sc�'=�ƍ��R8�Saq�G?�ɝjt6�3nz�q�����یv?N�(	���]�<�Э]evO�wW��
�
�JP |E���<����}�+Fpj
!��H}��I���薎�^�A�.��2k5��@ nIS��l�dgA$��"m<6�1uk�ḻ����	��V.Χz#���Ã�]0{p� ?t�$�r�f�z�J�u�y�|�<�YYS�t8�1V_؋�ҙM3BG�-���(�2r��z-�pd�6�8m�p�XgІ�qr�:�ܞݭ����-�UbP��_)��=xi�� >��8�`�5v!O���*Z��Z�h#8�r�+1ˆxeT���t������(�8�-�O��,ÖQR���0�P��_�h������%��l�mxwΎ��;[`��!�bS#B*�ES����.x���,-�7S�-;"^�p�à���ʵ�#k]*l5������Ӕ1��~���U!M��>�|Es��;�׸r�����YþjK�Smcu�ݾ�����޽�>x�}���о�D8��AD���'���lT�Z	^kk�9^�r�Qg�0i t,}���+�W�r
�8�Ok�k�;~���Gx�������F8�1*~"���˅Үi��s�3�:�� �g�����v�\���T�|�_s�z3��.����i,~���$o�<o�|�����w� ��Z�Y���)��@e�IG�����8�[7��=8h�F�	��p�B�tj�#��(�+�nJ���{��a��Ï�}�>��c��P��a`y.ܭ���&F�+k��.̟Gn�{F�J�� sF!�{qn�g)/�6��l���/*!�ą4O�Π%E�)���.�Wҥ���+u��A*���V��O������R��Wq�>�/Ʃ��UnR���J�r]� ��c}�w�Nt
_$͢e;�\C\��|�CT�8 ^Z��.�wJ��2B����k��.�Xow��-�r0Z����^�*�Ϊ"j;q�֭v��ڷ�Le{��I����,~Rf�c��]Y��C�p��$���Y��g��M=�a���j6#s&�p�dwC`9>�Q�,�l��4]�B��3��t<�,�E�e�q(L�q���+7�� �c�NFhzv�ݼ������:qũt����~_~�-������N���&���q�Ip��S����wo�?��/ڟ��/���g���e��O��s��[��wb�Ϛ�t�Y["жk�M܈{���v���v떣�����9�������O��W�Ho�&��؋h�_���W�+�	����Z>����Fǈ~A*�d�.�U�����*�@��I/�9�û2��)���������o��su�����4< Ĥa�E�\Ӥ�p4gY9���g� �Q���t���0x��vd00&������F��}BQ��zLG�g痲	���������Z�2ݼ��ܙ�����o�����O_���uuwA��H�*����Z{�]/�H��� Na��W�ͧU	Ѹ!{rrv�Q
γu������;�P�����d���Ϟ���/�cm�c�!=*䄵��!ޙ�b^��C�� �4%�������wA_����{���)e?��s��W�%���{�ih5�g��Ή@U�Y*D��/klz$��a�P�8:J����_x��9�Ps�% ��s�U?Xxq�S�{�����������=`"w0�@A��xO{�4����߶�ͭv��׎$N��:�Q�r�����@ڛ����y��H��2сkx<�rP��_n%����8sچx�$�9?'��==!�创�7�đ-�E7��/?Հ�	{U|��L�O�����mc�F�ԙ�_?��W��Px ��b��[�
ʑ'߃�C�3X%�άA ���W-P�:�( 4�<w?n�*��6�?�l��w�1��O��=�4D�T�jJ 4��]�۷���P�Qd�*H<�kg�;���z��H�`�&0�]( A��[���Ma�?��X��¾znP����6��S��H��^��kI������(V�P�ĉ"^їQor�&
�i� d(dS�i\��"_��,�񑸃&+��h���M �86,�� wj���ZP���P�yH�ӧOi�7w�rڟ�/ʲy�/*���r�jRTed5&��g�7�y�d]K	Lb)x�Pv�t�x�AI[��D~��4ʹ�N���D���L]�o7�r���{�����w�h��ǵ;򵽸�ȏx�l9ǟQg��iwgĄܕy�NՕW�d��(¤��E`�ȅ�a��<���i��:Q1���d�2�?��m߇RB3~�(�\�&���2��_��0\Y	<�f9\��nȴ@��X�C�.}ӼC��8����f������W8�Sh�hE�:"w�y�����������m�yA�Ӷ03M�5M} �
e줬��ȁ.m�_Ǯ��#
��xQ����}�i��Oʹ��������}�>���Ï������v��g�~���m��C�Hϩ���u�m�x�6n>hk���;mn�F�^XkS�m
�b��F�j�f�A�P�t"�N�;{�\�9��K^r�Ƒu(�ܼe�����cTÀ��9B�q�k�׮���o��;�0c�;�DeD�Yw5��(_.��q;ͤ#y32��JN���/��m��R݈)eT1��-YRt�IK�'�+�,�p�Ff����lp�#;G5d��;s�����nz�Y�O�?mO�=Aw�F��mk��m���������˙Z֊��N�2?�/;g�M-�Զw�.'k<0ލR�|�s͝xݘ����]��.{�e���Z�{� �%y&�(ԡh9�|ls�kм�U68�o���:e����R`3���e5^�y}�-"�a[�t���������U{�������P#m�"�vN#?N��X��=��i���Y?��c���>ո�^�+P�m��3�0h�շ�t����S�p���<?I��|/�{�o�4�V��2����v:��v�ڣo���~�е����"G0�C����b����}�y �$+�S���(-�WhU�
�52�C���$��w����-�<��Y4�_�8I�u��+���N�qD޵�R^=���|iǲkċg�+w��v.�Q5��(WFG�D�F�tL>�n҉�����^'
��� y���I��C�����fjD��v,�k޸~�ݽ��u�zpiێ��o0�v��dadm�g�F�J�#��Is7:{M��]3� :� ��/4��U�t2������'o����̑��l��_��헿�u�կݾ��ۜTn/򡇻��+
D�`���LNT�;(I-V�4�<<p��ɺh��'�'5���e�OP�-�l% q�ʺ,��JN�&�k*Vda�w�}� r���-N�2bэ�R8J���1-�|�����,{�����*��۫�*Ij��(~��OF�h$�d��(q�m�a�^�j�l0�|k���0f��|/f��6��N\M#q���~���2.Eo�9SB�Sfu���aPѯ��d�K1�������Xk�o�o�5��U�%����r���#X��BY��� ĩ6҉�`C>��� p�w��Y�b���H<�A��{FF	�/���n]*D3���|M�[�1�
ש#�k��q�>b���f9�B	-�*h��rW^���V��3�s�凂K��7�uM�k@q��(�P���Р�^f�s�.���\�����w�*[���}⋋b��$(Q�?q�C�H^��<��g��Z�\U?�㡛��#%�o�CY
8�Z�`5mP4���	Nw����O�5�ã�=�^�|�v��2,�����ڔ�S�Qa�YJ�b\���"�Y����i0Z^�
eGm9W�"�m���;�-�7�<�X_m�n;bq/���L5�G������P�)Õk�����Жu�}��K��o��	��R����?��`���1^���7g^�q7<�`48��j�0��]9�� 6���qJ�#I�Q�6]�#[��ɀs����/�"��~(w��>;��n�(p�ql�Z���l�۾��79���]��!��a�j��4��,x�ze�y\��j��RR�G�Hʘ.PO`;��7n���?h�~���hw�}��w/�9��PЗQ0��餱d{"�{f�#)Ό���g��f$k�-,-fV��Q.g1��Pu)o�yW�;�/��S��S���}�΁=#�����S��$U�R�>	N�5�	)��T�taV�/����c\x���F�� �3-�{�3;��ݐ���=�a[#]�b��x�8��(i�J�S�τ�Y� �?�v�'�7�Ӂ�״-Է�O��y0�v�R�r��u��ӧ5B�L/��(�ԛ�����G����gV�ӵ�W\(^u����-;������{G�m,��TiWǘ�\��cN�âq�dR�G�d�i���C�f��ԩ�άO�!��'k;�U�����aЍ��3�9����z�]�'��>�ݳW/�k_��ލ՜�r��$L��YE8)�wtңen^_k���n>����Ci&����j�����7�Y^^h˫�muh;n\���C��2nݺ÷uxf^���w�!�����0����z)����4�`�\vWo�n�<W8�Ӄ7�	7�Hg��r���K�E˕�����^�6l��fgJ�Th4��S
����u�8-PCI#JC�{g,e4U�t0���AN�tZa��9���C�֨X���X�pI*�˯�7��aNz�
6ë^�{������)��B;�cY��t����:W;�b��H֏YVm@"+�������\��\��xcA�+�ʕE+�qqwA�=��s��L��=z�}�O�7��~���-V_�����wvbيt����YϾ���4'"(Z����4����kmw��t<Y.Σ�����Vo�
��-¹�,Sz0��G(��5�?	����:z_Dn"*��QQGF�FΥ�ui�TZV�J��B5�Z(��P��ux,��L�Q&��=�XEӑ��RJ3-��X�p�}�9�aC� U�:�#���J��G�4�k������hd�7e<Ӕh�-8	�X)�L���Y�`��Xך3
^d,�C�ȩKKKp��s�W�j`9Cx��='2�F��=s�-8�%�R��b8 GAd�7-��	��k4BTPl�4p��x�s��|֣�!���(�Y�K_�ѹ믎ݦ�:��r�j���sG�jK:I��I�6?a���� �+!�˼�Koe����S�qJ��h�cF/'5��1�,G�Gx♆�U%��W�YZO��w!�=_����;ӤR0ң�ҭ�/&3Y������N�>UP��2��Y�v-\�pw�LϜQh��A�2={�=����W��@�T*�H�Dʛ�t/N��r\���w��P~�g�U�UI������ ��g���Dfz��\�B1�sc�ݻs;�	ܻx��4��6B�A�gd	��yF\6�_��S��:���\�RJ�AU��l=Y71�)z{yI�Y֙k���Jp3Ы_pߒhn�w��lCjǆ
+��l���H^�"��I6�+�j���j�G���P���5���J�N#s$,�-n�Rxz��^<{Ծ��W(�_����6�r����p� *5ă�Q�J�*�z�,iԩ�Q$�'m,�9r��s�N{�>����O��}��O1��$�f[\Z'OG�<�{��딉��5x�X�2�g|:���Vc�^\w�\A֮��y�N�!,V�`�ò1�����tӌS�f�z���<&b�;��w���W� �(�"�R!��=�+�*>Fo��s�����v��Gŷtf&���N��:�B�߆ހ��,:2��5CY5�XGm��i�4@�ӈ�'�Ƨ��)󶥅#��J8�D�S�ˑw�;�w݊rj���� �#���&��~9��iy�U�	�X����B�5H����m����,���j:��|�OED:��6��!�+���L�f݂���It�b�^��,���U�,��HG��wӔ;�0hn�A�l�Q�|gG����	F��o��� ��ԷxO~��t�)gye;�R��0��7V��;7۝��(/� MFG�@�yH��3s�����r�u�F�{�V:�����k|�0�����u�	����;a��I�  @߿6��7ߴG�����]��?��+��4ܝ�v�<Y��I���^�jd�OC�B� '��ԓUFB�]��0�C�z�K{��N��.� ��\j0��� �q��׬ݲ��3k�	�8оr1k��T��k�`ɋ���-zx��=���r�e��\ԫ��Fɍ���׍,ٖ������5���ک)m�v�v#�LH@@�"#Y(�Gܖ�E��!"�LF�j|.�����)9*k��s�����I�Z���oޤ��7_~�<���}a�<�����]���	��+�K�X�)
*���<�

@��GG��=C`�F�.�,��G�*�
��U1dH��5.|JE�~��*)�$<I���w<JcM���7ed�h؊�Z�'�%�6�`Z@��Rf*Fd��4�*��"N1�vMF�<N���O�N�SC��J��[ O8e��4�j�E\�۞�/��B���J!��ң�B��ŉ�q�v��FV\`�Bd�N2"���C���8�bd�~	#��0�>T�э��:d�γg�8��V�4{��\{s��ow�u0�pv�S]�����%P:�Ttl�T�9=�1��.�!��%uuI:L��y(�P��)�|��ЏPY�d�t#k0���R����΂�.�Lߴ5�����@��3h�����}�xW��'��s>�H#�z����c��|1.��
pJ�]jOyZ����+��+_/F�5�# �:~@>�N�(��/�0��m͢� k��a��I��⿔��Z6�4@fM�6���k�\q���pV�@*��7o^��8
����,Wdf	u)�_��\B���]�IT�N��x�t*���v�6e�!ʅӭ5V����H�;7��}��h�?|�}������пk�Dn��&�:b�h��*�*��*�ht�^S%�7d��y߁��U��)����Ha�C��,l����Q5l�t�:6C�a�Tʷ
�����u��x#���!���xa"��]Z�a��3?�K^��*������需J2;���K�������j/�߾�����_�7��g�2
� نEiǻ}�)I��S��F���!�Giy�X��>�6P
?l�����>��L�[\\oS�K� q�J%���Gd�������IT^y���v�9`��ʢk�4�f\l��)��RA�#�B9it�8rڛV�lO��Ҙq}�U���]�2k���(��kT��_n)��h�H��d��]�Π#{�� ��{�2��\Wb�`uW��cTYt��I(�1�/q��~"L�1�!�"��.�x��|]�e���Dv.,�S>��A;�m���6�4ܽO���ݻ��.ϳ	o'_����7�����Wt*Of�	G����
})��v�`2�9]FF�����`t1׿jdY*���*�s�d�W�?g� *@(��ˑ�� p��������ݩo�)��@��������Oᙩ"�Q��m�U>k��>k/_���U���G҇��$=Y�6�F`ҫ�8sc��ٸ�,tX�G�l������v��u�����;�2v��-����>�G}��q�Ȏ�t��Ϟ��~�~�믁�u��C��қ#dVZ�$`.���.]�m��y�)����*	�;Kb9�Ȫ���*a%c>��s*�XF�������u6d��	��&5�9TDQ^����JcK],�hk� sÌ��L{C9/=�Y��Q�_���6!�U�^SR��o�_:���'�9�d/�'D~:G�]��Ŝg/�ٱ������
>��?hd]n|�Q\��,���
�>��O1�UxU���U��oń2�1By*Sqn��h�-c �08�e/�g4�Ý�W"3�L*㺦K�teO���R�7�pj��5
�h���{y���ȝ�|��jdQ��l�,��*F��}��B�ϗ�]��W"�/�E�^&dY�4�Xeh�t�-�,�)x�/f�8>S�P�5���AA"��kd��۫ú��k;bXٻ�i��3]5b�4yH�̜DD��BW;����<���FE#���v�҄� 3f����קME�V�����CF��P��o�U�D���&`�n�j�z�����Jz�j�jk��(/N߳!Q�Qq��Gq���������4��*��s�S�����a�e3���3�58/�,|�Ry>ɯ+�$ië?��.���h���:����邎f��)�-��$e�AU�-W����	�<�X�fY4�2��-� �S>w[ps��8mЩf~K�(�9�&}{��{����l�+��T�(���Z>�F��Y镁e�5����B[��x6�*u�Ϊ�{���b�_��^�����P�̒@��(�X�u��q��"4�]0}�N��Y�޾�\r:Kd��"�T=uA���g�7�a�.��p�T�\P���}(*���9�\o93y#�h��m}e!�'>h�|�Q���ڽ{3� Yȿ�H;j��:�4'!G2F�g��F|��2N��t�wF�U��$<�p�J��@�gG��j`UҮ6��N��A���չ�\�p�$�eT��I�K�!��[H�D�L{�PR��;!ͻ+e�X�V�{�x��>u'�6��i9����ڄ�9�gϾk����l_��o��Oÿ�(��� 1��/�g�rA��L[�q3��/����j���������ڧ���}���{�?n��7��y�`P��'��}.��4@�kd����?yO>��L�ƕ����lOm8䜝Q�1���5�ȑ���Ȓ�e��T�+��O��@6��u*�`y�q)����K���:j⽵d�ا+��T�]���F콯x
��b�Z�}gۣ�ԍ,]:����5�I���eu#F'�� (�z琰�s������
핇��'?�9Y�anx��L�6gh�ʬ�����d��ƍ�m�]sIC%ϳ���c��;���Ehd.儔(�d�k4[�^ݍ,��f �#]�d�&k^�0,�SM[���x�c�+K�Ȫ2�S� 	������Qߑ.jz��]y�w�C^$J��J2���7�>��~���=ʿ�p��1�^�'.1y�<���{��>���j����^!lN�U_�^Ż��Ƌ��`~}��ٸ�27��[km�k}}�{)�,.ډ���q7�Nc�=s���'�������o����˯�G�3�rO�,q�o��ů��;��JVyӟ���B��]�X1N3��2����!�1+˒�|���<23_I+�:l��-��;�F~���8��H����N֍�2�j���z��W֡�C]���:z�kȍFH��8���!��Yߝ�]Nx�|���C�W8qi�}t���R�$p͢:��"��`d9�%])I~�,OO�J�_<V#KZ�Y�#����"Z�ӣ4_"��s���6�0}[����!{8e@	����շ�V(.�޽��:�u�`I�A�4
b�]�M�*F�v��C��h*V#�����GV��&�唏�hsdS���e.�3�<�3r5��AP�)��Ѭ���'��MyU�bl�Z���1���Y���S�OPf�L����E�{����c��9e�:�3G}���u#-�Xa�R�G���!����������:?ZC��@(�����^N*�^�}���&�&���œ
٩,/�/�_
]RL�	 ؐi��(ݿ{/���Kˉ�bl��Hj�Z��Ű����"��!�4�ҋ���m����Iø#Q=C$ҵx�w�󆦦�&�6	�J��[�:�A��6�As�W�,�u��ed�b��s��2��;�uMZ�"�G�?4��)L}YwQ\�q�F�7�6�d�0hkb��^�q�z�'쉛�%�N�3��J�Z��l��H�,��׸���
[�\�X<{�<��ሎ�@�mc��J
��*҄��O���76Lҝ4Hiм�%�ɺQir�)�ko�w1��f4�5~�e�
wt4k�|���M.t)��}�\��k�Z�g�C��^��kF��x�[k��͚��W�f���B{pO#��.k��)�9�U~#5U1vTB��;�% �OY�=���zC�]��	�䞲SO��2��8t�Q�wG�4�4��U�4�FS�8�!�F�I[���B[�)2�E�{�ʥ����on�eY�+W	]��Ӷ^�qQ��r�H�so��%߳���UvK6ȴ�������o0�����}{���=d��#��SG_��A�+}zUVɧҏʝ孩\�$��
[In �L�_Z����}�����e�^��^.��4@���fٕ��M�"���M�o��w�^�_<_(#�z���,�����h$��-�k̬G���zv�8�J_{+$���:�'hj�歬�N0��J�~
�N�����?�x��
�����!��xϡ�!�C���2�#�ʣAz!���ed������M��4g�[7��Oѫ#}�q����r>��g�۳�χeﲉ�W{�U:�{�]^��՛(�n�TgG�<��9�=}�|-sꕲX�1�g�m�t����R����z�ʺ<�y�,����I]�62
�r���ӎk�b$v���N�C\u�c7�J];������X�*T�3�$�i�榑y���{na�B٪���)n��������8�;bd�G��������N�l4��ϑ-�bJ���!���E��ܼm���8e�X�L��f�"ry~����e�4۲n�����o1���o~�~��7��k�F��y�]���TtE�U>�w�}����ҖĐ�W>�3��\�!�//N�s0��+%EAϏ����a���'��1����R�c�ռ�(G�I�5�U>S��p��U�^k��k��j�)X�����q�M~0�ղ�,[�������fΑ��2��7��p�=t}u���8��-F�L3�����N�.h�}��%�ӫ�����o�#~
�K��;��U�)~�L~��Ͷ�`�bJ���@�"�Q�@E޵fo�<D�Bm�ܿG:7�"F�ʓ�)	Vnz�
eqc��wt�`_���u����3�
u�U�����tk��o��K�y�'_�,`�C�ۍ,����B�ˆ�j� ������(�1^ciciaq.~n�w��)�:�^���w��b�8�3�P��q4G��r���Ҙ��zU�n���ᥑ���� r����I�*�
Sa��ф��:�0��V(������>�B�Y�4����zM;�q#��F��TfQW�r��naXmmncTc`�:�W�I�r+aϒ)c�^W��o������c8lm�Y�F�4FV�s�qz�#=*0T_5���:q�A�z����#+S� �#���}��D�5�􃐄ХG�
a�k���M"4rU���*�$��^����"�E�)���cHf�I� J��#~���ܲ�v�2\2��8�<:(I���c�����KZ�&�k�����Le-��{�~��q#�0(�̳
i���i��� ����Ls"�s��xǩ�ـ�X�R��j�(�	�x #i?��/W�
S����<oI�.`Ca̡*so�g�����X[�1w����!JƇ�;w�l��&�(6-�k�3:���N��;�z��ý�s��OW]��~1H|�a�{�)/7ո�� v^�wV,���Ec�9 +�ƈ��p�̽� 䵝%4�A�>;�o�q¤���y7�_IS�&��%�ܡM}x������8�D�	��k�_>i������o��=�e;�ۤn0��͞m�V��(WN�b����-5-L*��m�Q<��O%����_Z��)�~��v��'me���@0G�)
3D����V�|)��!3�'��������pM<=��s>��h)�
��xN�>�<IX��ѯI\%FGl�˗U��7uvL�idY�c�:�qh�Ѹ�"�:�Y^G%xG�U{\��>��-iR���ZF�;f�fc(�Y���^�SR��ik�?�N7�.�>#5��ـG���mB�H^ֻ�s&�#���ſz������]��˯����W/��W��&���em��lg��W_}��.����G��'��~��Ǐ'a�N,���ʡS ��U��F�A>X�v�i�;+CC��,��iP���1�c�E�w�.�d+��8�<�ŵ�4b��9�_5���9S��n�4?��w'��8}6�&HǵS���@�a��	��pz���n{������FF�m�pR*�.p��#Ó��K�mn%�{�v@:Ϟ�l�޼A�?N;�:W���v2�:e�g��#�O�%�:��3����2�n���W��oem����z�܌b��΂���^���*��kj;:�2�t;��(�y����7#�	�ːX�K{���D�ߥ/y�d�~yqS���p:<	#~F�팉�.��UU��YFV难�Z.;� �.�|Z�f9���ma���|W|�������e' g-�e��t�h�{�ux؁�T���]��=g����i�&��$P�0�:N�UhX*�2��)ZA�;t���o��˽���A{K;���̯�V �(��- B?���*�(X�z3r���
��֋˫���~�ߓ�p-�ɷ�]z9�7V� �CR�<\z%�K��Ҧ�r�qvn:F���B��n��633�jnf&�=���
Okw4�-{�4�l0hh �Z�UʱxMϱ�_Z4�To{#\�������3\0��.�u#���6��Թ��v������6�
ͬ��@��^�Y�%����J[[Yͨ��O���6�.�vʽ�ݶ3,��Y�W˭�5�l@z9CWօ��a�C5��BRWոW#[
\�a�Y�H�˿\�j���^��#�P�PA�货��G��2�����.�� L1t.��@)��W�p�U�Cj�!J����Ǝp�o�u����\�JW7*��%��//qD3}����Xc[��H"GJ�6��Q��������g<�(>�װ�K�kk����F�QvGx�{��u!�4-��EuM��l�8�T�����+��6��l��-�"�ݕ�b7���s��ٶ����\_˦��~�Vyh��1է�ѯ�U�e��ҡr����4?����*7z��(P��}0��Ebzy���V��1�i�V�;��~V:q����
�=�����u���N�&J
��~;��j[o^�����������;����v�:�ה���
��g�CZ/o�EG b�O@�N��zWe���������ۯ��o�l��=j;�Mg�2zR|��c�m�6��ۑ����I�(t�S�\��,�յ��޽������Qvt�Mբ0#�-�)I{|Q6��>2��t��\b�c����
�G9RyH�A���ЛHr�c��-�g�����M`۸�ͮn��j(�c(�*�1p�W�IR�$���65~��!�g������N;�}�i���>%�4,^� ;R�[f���k� ?N��2&�f���>G#�F^\�-�htt?�xe�48r^W�-iXZw�'t,2��z ���Qu�7�rX��\NW}g]|��I��(�{X�f�h���eeTE�	�w�뼨|Z��qqh�ҷ�$���[��ʄ�J���G����r+>��22#����9�s�%��:���\9�C��MC?���Q�FR�u�]�O5QƵ�u�hG�����mz�H�o����G�@��u��aϳ�(g�m� �:��3�¬o����q��7��_����_��/�_���׿zҞ>9h�^���Ϗۓ'����^�o�y�=F�[gȨaX����4��y�=z��}��wY����b��̱�͑ϖQ�\>&���q܋�~�^�W�iQG�.��6��C/�u��}�}=�9�+��0vr��Vv�׺w��a����hUu\�S����8��ώG���Z�1��,�������2�
��|�r�������Z��&|?��R�]D|�:n�;�dix�.�b2eZ,�l|�9U�d���P�0��D�A�Q�W���EM<O�v�A������ �0��C(��!A��]"�k9}����dg�̻w���P�1����'M{�E��s�����9�H��=�H���X;��͞B���h1!����1�sp|
��/�Jb���#Y����AF�h��
�=:u�г@�~�J�$M
Y�� ���<J��%�~zuu�--�0�9�����p7OۯQ/-�ŊPU5��wZ)Z�Wϡ�7�����u\��q�$6(a(����|���cq�?��;.p�{�IC·��(�=N��:;5��+7�����%LE��JO��Qۇ~T���j����l���iD��z,7�@��2}�"Ho�=�c�3{T4ŋ��2���X}$�t����j��{3ZQ�)���wx��Q5	��e'A�_�ȕ#YNt�K�v	�<�s��+WƅW^�.ʑ	4�1���'�0�<8�̩e��������ɚ��njG��.h|�c�,S�yz��g���j�L��'�P�C�i��+�a�r��#Y����20溭��x�Y�,{��+�˂a��K��4T5�JG:���)�������G~�nު�%\����.;��9Y�"��\P΅�HH�J�ʧ��O���c+�E����W�(�����y29� *,�mq~�s.�?��=@~���=�2֡�\�4�B�y�4́:�ZO�\�������E9_����Vu`���|����n���#7�Ⱥ�Cٶg���ꈗ��Hx�ڨʠ��v{�$��3ʉܰ����rʺ>��b�%�)[R�A���Ϻ�4�'�t�R&�aX�;=�����I�ۓGߴ���b��b���MO�!g�Ń�N��T:�E�r�o:
Tr���c�K."��ե�����W�{>��ɷ9��vQ"�3�X�few<�i�T��\�����������vԈ8����X�X;�줲�f�!��v��<��-S��tʸu`��	�F��c�P���|a���-W7�H���,H2�`R ����,䅆�W��P�%"�-��&��9��bZ�Ok��[����[d/e�CD��N�JW�oh����<�1)� a{h�s��9�c3�[�B%7�X\r�7��F��}�V֌.-�dѻw��7s$�ŋ���o���7�;qa�i �Kބt4��u8ݞ�C�b��n��K:��/�r{�v�х��t%�b�BRo.9p�k��$@���D�`�����v&YOv �L�)�L,�Ӵk�WF@RQ� ��&�o�h}�9�7ӡ�쨹(
8�wO0�޵��`��p��a?����N(����yq�M�[nk������[[�{����C��i�^�k�_�n��>�.���m��`=�p��0�����G/ڷ_?n���ߴ����=���r4���E��@�y�[�����f�������pQҧݔf�#yF{#�ţo�����˶K��� ��N�O��T���t�}�Q��"�ֻ/���n��P��'�E��w��A�,�L�(yx�e+�^e)�ay�!��>uaxcV_<�s�W���"���3��Q�-e7k��6��#������7� e3 �2� �l]O��$�� F(�1T7����k�a��h� ��Ynwy�˰�P�}� 2%r�&g��V�;�����)=�袱�R���'�.&=�)!��ǝ.�-�1��^1���BC+��X,������o�^�Tj}�BوU(��Նo
�X�Xx�,ù�e9H"V/���p����i��Dd#+�y�)U4���q�A���L�t�
a�UX*� q��@����1�kd��y�E'�<
k2�ArEq����{�O�z��;�8�uA3�>p�ؒ{�\���>&��Y,!�Z�b�e}e�U�jgw7ƺ��;<��`�
�s�=�%F��*{���r[^�vz�����A\����r� 
�Ą����S�7�x�U
bD�0�z�_*W�&���`�us��W��+\h��Ҹ#R�|����4��J��+@Da�4h#j�J璚�n�ۛhgF<6>KC܍,{�'f�a4���+�NѤ`�����]�a���K�n�:�=#Nʜ�ߞf�$;N�?�o��h�����遇�Q��_��%H�45������ۃ�[���۷(�Y�qpʎ�TV"T.Ç�����w0*^�w)z ]�2|�ڼx�C]���Cc�Ml�v���%���L�}s�}�ˬ���ǳD����T�)	�T�/�}'|���Z%��I��{���zT]��K�S���(U�ͷT-r�u�h�#o���N9y_���Ϩx��;y���>�G��X�1;N4H��YȀJ�YS���E i面R>SO�9�W�����}G��lٷ7�7_�l;�޴ͷ�۳�(t���'O�A�z�B�a��+dZ��=-E1��y!�]0��ԗ2�O?��3A<���݇����-������yHK�cy���[�!��{�KwE��><Գ�����w�_��{↧��c�eBN��}x�Mi��#	?�'��@��m{���Q�*1�:�r}��	���)~s&L�keWW�C���xx��U�l��Cr_��������Gf�̸�8Fҏ�H|�]�z�x�D��'L�{�S�(/��C�*�Q����.�(�v0��k�4�ԑ��a��v�;��Q��R}-��+1fl�^�z�cp������.��D{��a�N������=mF����N�½�b��Q����t7d$N&�^�*O�VFi1\�#;��>
��[�|��)k^擯2�5j���A>���?�{�}��Ӥ�샶�83=��<hO�j_}�=�x^N����C-yu����������yf�g�^���Cd��1z���V{2l�����ͷ�g��g/��7n���޼ގq��ɫ��W������׏��ܿ@��٣ ;��̴=雼���F��r��m�>���{��ы��׊�'�p�I����?���4/�L�w=����e���P�M����#!We,�v�W�`d�ܧS+�����L�]���9����^������Ӂ���#4��4|�.�7�Y�	����l�����P��L�������_��i�����z��u#��%"Lcl圥��F x��'�ۣ��R��mأ/�,�T轹��"���IU�j��5�]��,wɚ�$=�DUO˸�(��9����W�͋W���ghn��b�ݾ}�t6P�]�f.�=4��V0+ x���0�<��:k[{�ed��yA��`�b�5f�?��y��=��)*�cZ�Ƶ:p����e��Hl�<£���ѣ�����db�*��g�R��.�dz��S�V��9���Xm�;�g��;�!��"q��Bם�S��i $T�Je�pxG�2J���8%�c��z�@c��w��
����Q{��wD>��w��s��p�F+Jjqd���@w�n��_���>:�J�;�8�����������LO�F܅�
t�؜Bۇ�}���uL#N��`��@#{� �q�2��O�ۈ�!,5��X �)5V5"�C��YxCD�!��8����7y��Y�T�A�w�cb�R��#���f\�0?��,h���u��5�"�dҞB�m�	[��n��;w��G)S<���ژ�?g���f�����O�jlyL y���`9�ۻ�z�mM#��`O�/�4��d6� '�Ĵ+�eɶ�(N��5{� >��;V9�?C��t���y3
U�(�!��Ƌ���ۃ�c�8�)�6

u���D�K#����Am��Gi��Aҕ����t�����3h:unX���U�x���S��q�<��gj�nt����<��u���o^�h_|�Yֵ..,�wZE�RC��q�F�g��9�)uF���W��\ ��N�ū<�{I8�{0�
$��+��ڮ����N$�6G})��N!q���f��ߎ2.{N`��G��␦����1Y ��<�Y�Ie%ӵ�5�G�����
f��#Q�%��7mw�u��ポv�tG;�� y���w����;����Ѵ��E�z����������٣/�c�����K�_��o� ���	�A)�^�\�@�譇�(ևp"���$H��X��Ǹ���[Z�����w�����p���U�QTp �C��uV1Bʇ�[�a^��:*
�c���(�>���<o�cG	QT���{肌l'J��Ó��
�r�ΰ��َ0Ng��k�{�/�BI7�n���q|]#�N�
&1$2�<�hn�� �X����Q��D`;^�
�n�A��p=�4���,���)��\ۭܰе��1�ԥ���l£��{���v��N��G�B������Nw�s��k�w1D���¹˝��e�(��9��J����{�Ƥ�n���7ߴ_����7_�޽y�1xď"ʽ-���C��ѳ�ЅrC±���\�k$��bR9���E�u��k�5�;;f\��Hо�f�T�gYS�-٥mz��'�m�R���٫!��g�!�k u%g�l����?��}�Ž���Ǥ��q:�4m��̻��o�i������ͩe�k�..��,�h��]n����W٩(~��<�E}X�Ʀ�w���n3#�O�>mO?mϟ=ko_9M�%�/�ӧ���� �_��7�7��㈌���n������1�7���k"}[��xoۖڒ��z>ZE�%u��NI��Z�"�|��uO�	�SКzf:�m+�?�|Ƃs�fuH���Ś�� ua�zW�������$WV���>��)��ѩzxγ�����U�W�5˸��b���{C��T�����U�p���D(<	�ptXt)7�5{��*��s��αi"^X�֠i��<��
=jh���D��
+i�JEr	+'��ʳq�7\�\�h��K7��K!�z��t8�x"���T�<w�vk+��ֶ#*#����

�U���wﴏ>��}��G�M�]�T6N5?�{a��5��RF|u�).|�,Q	"��}��k�*�u{�ep���C����j�`�S�U���x�6�'��4�#p s�=m���Ƭ+t�X�-R9ѫ��b�_�lY+��a䆇�+�Iy%�(�0lz�^�a����8쩴!�fC�qw}�p��������48��~`]L��c��Y�0�@���{�
�=���DGto�v0�в��`@ (�?�*��K��Ͽ�u�Qg`l'Nz�-�z�p��8����8� �q�zx ƍ�1gJ"~#�i��9=���(��h!�.Aky4B�C~��G�T)W���.\���S��uxiF��+�V�//mJ����͗k���|[�?�Fyi�ttI�s�j����p�_�i(�iٽ*�����Jp{�b�C�9�c�o��ap��T@7H1���E�R�F8�T%�����2J>s���x��}�*�JG*��(0>?�l{�� ����˳ma޵����@�F��\�./Ei6��d�3�3?������~�3L��C�rN�ŏ^���CX��O�o�w��?�Q	z��a5�1���p����iED�:%	�:Q�8>t}�����c��oړG_��O���Q{��Q{���O�iO}�}����W۾��_����?������ڋg�b|?jo�<k�;oH{�6�8�_�Ǥ5d�J�5��k*��v�Meg����I�\�dQ��i��vR���U��v��=�]��67/o�Y I�zW�WY�>uU�ׇ����?�E���|5Z�������K�\�pY[݀��3ZS�P��j�0�;y֦j|���_@�mee��@���NלrD�?�k��A�gj)����<�#Cl��9r"� �I_\�S\;�lyY�4����m���E�����QJ�J���t��R^&?#�����z�������޶�̖8"���52��&\k�s�k�Yy�h��T܁�sE_�A�۷��SJ����P��o�'��Kx,w�WX���Q�^�F�7�x�^KIu�kɠ�Up��>����R�����æJ~���/UuX���|`<ۣ�,byyØ��6]z�������kx�9|�?����5۶���vJ;��ʣt8� !�����ZF;!��>exG�����{�}����������ū7�՛wVO����o���_���������_}۞<q;yw:ܣN4�-q,Q.��6y�� �4�"a��:��>t4��8*G(�%>����{.�~���O�!J�� �����{y�(X�T*���x�	��J��K����G����t��Uk�φw\��/z�zA�k���M���2�v�K�U�S:��
Y.��n
�p.[��LS/�g�kpV� �?�6b:!�)���G���2�JwG��u�}�FxI#���@|� �I�h���>�����_�Q��?�'��)��#a�^�-�a0��m��$�@=I�'A����U
SAn�*������y_��?��$Ja��f]A=W��7�w�o|�bF$��B!�]����z�e{�hdj:�
�A���?��x��ސސWa���'-_�?�V:iڸ�3R���%*���Hх�3�5늆խ�ݭ�Mj;>G����ö�#|s!��{���F�ì]��|BXw�2>^��.H4Z�;[m����)w�D9u4cCk�M ��~��
��h�F�Q���(�͉�T���k����t��|e��A���4>��E��^Ư�)���]ml�$&1���J�)�p��<�g. ߫���4wѴ�e�h�1�ܦ}z�C��Q�<�rCc�2�p�#n�%��|2�f(�]]��\����aF�����"V�Pi�] G�Z/�IY:�u厉��ޱ�[��=;)!�ӧ�]y%lN�y��M�Z7�������c��}d�%OiG^,�ғ7��RWUG^V%CE��d�+��k�K�xw�@1��b1ݖ<��^m;*2J����͖?�%��c]�����?��W��L7���u�/��2K�Uo�-;8��2	UE�s�X�Ƨi�3����A��C-稂NҺd�gM���Ѽ�)�;���ރ�Ͷ���l�A޼j�޼ho^=m�_=����Q{��;�������}�k�/y�}�z���w@����Ǌ�!�/�����eg~ 	G�F<hd�S�<yH��E�"���)`���uڼ[���;����meu��ώFxW��{&�+��r��z�����{�cXu?`?^�?�{�0�����m�m��8�X}m2Q�k��P��}>ǳ	Ɔ��nf�Z؇gO�~Y��3E����-y1j#@yT؈�*�؈�N^�'Uҝ��aä]�W�KeK�V�Vqmҫ>=�[z�q�w�P2�t�{�5�q5άs7�q��J���pY���zJ��I�bj�����4v��*��_��C�$�'���3\M]��C{c
�6��u�p�iA�v�S?g�2Ȏ���.�9i�Qf��!��N�IǶ1�h�l�TVkW9�,AN_;�.\W�:�����E���0M�5y����0��ڛ=�^����tpL�_vhd���t���/G%fj�2dw@�4�y���4��v
�C���!�r ����`��>���(>:D������Gg9�-Q�tqe�.����`Vy�Վr�D����84T�}���߬�T���9u<|��YѶ?�U���?iDMx֢�2�l�(ע��W��?��]�:�v_a�>{����iy4�Ee�xE~���Cc�y`Y,m�,���\ﺱ�cη�܍�j�Y=�@x�(���B`\�KRM������n�&ސN��Qx� a��R�+=#E"�j/0�܂���-�)$�A�(s�#����>����?���O��?k��?j�|�i�w�~�Ntg<�*�""�mh�%n��CA�Q��dd�_���wW�v�w�~��˄�J<U��
��r[�h�r�E\�h��J8�TC���&�J㉣<
[��&�0M�.�L��1��>?6���9ep{��WX����v<S1�Y���:(�|o20
��yj�=�h�#,�6�������+��ְ
�Ӷ�u�9՛Y[�v�����V���&�=�uBx\�Y�*鵌��@o������N�H� ��[�ڰ#-�L�� x�I�%~�IsҪ9�
J���(%0�SI����}�f�w��\��F+W<��������tL��#�'g�Q��0��O�n���U�-�CG�����<�%��'n�в�H�#_��f<��y_���]n3X��+Z�4`�(3K��iO������TD��� @�2�J�C�)����5��߇�A��`\�rY�(-_�_����]Y�k�xy�Ma���οj��\�VQ�$ňw��7o�F�H;�VT�Sv(�P�-�[>p�,�E:�8�0E6��a�W�)yP�0���鏮Es��Q,��l�N�#{��p�r1�u�v8MB��5��Q�R�*oR/o^� �P����w�����3z��Uc�C����J^���k5��Q�&@P�ENS?�ě w�������f%�2:�qtP��$*iϠ�ϸ�*H�����)�͗�57�ᘚ �s�]��-d�;����~���w(Mo���䐽�/�io�	��|������Y����Q����sn��4c�x�]��r�/C�zw$��-eKpG�0T�WVs����:�	ON(��\�%Gɂc.�+�����U��틮��N��rUy�,z��Q i�)�¼���r�R�[N���)�8��&���)�Dw����Y[@D��L��Sm}i�-�`|����+ϩwG���]�k�ҕ.#���i�y-��\ʣ�bmx1��5��B����]}��������)ys�}9x����y��E�O7�qꯛ9��X�L��޶[٤s�v�)2R�='�ֆ,�Y8
N⪔�7z��'L�I�?@
�xM[!���R�ۗjK�j����1H4Llw��N�s��08�hp�L��[άv��妝�rB�z��� �qۛvD��\`2KF\��&h�Ph>>D�o�Cl���J;[4��R��)�k��w�'�D�t*�z�m�<%.��F��L���O�,���E�N�^@�҆b$:�c
���,��@S���
�>F�#�Ǚ�vŃ����gۮ�U]y��N�y^�����Q��=\����Е���ǥ^|Ï�F�m$��R�u]����^��u��K>��Q���ϻ|�_\�R��e\%�ļl��bܙW��a.�
���y�ݑB����U���n��|��U�0]'Y03ʝ��}������n '*��5Z�WN�R x/@���y�}�ͷ���Wٝew�u1οD	"�,�;�Ǡ��/������'�~���?�Y{��(K���Z�l� �Q�3��
��x�w\�K�"檋�����e\���D�û�-^��G��ʛT~5�u���Ŀ�4ˠ*�jh��S�@���<��pOOa�|�]8�1K^��t(�0R9���T�F� C�S���W*/���"����Në�u$�s_��i��0�-��_����I��q�#�a `h����c���V�~}o7#c�P����պ����oo67�[���ݶ�V���;�o ���ux��'(U�CҴיpW,����Y�̔��i@,檱��	P>�$eW��Gb�`'���v�KӞ2�֦�60�n���j3�7�5�/a��e��m��r�w
D=�#V���z��h�K(rKW�Za�iX9z5�Q�y�OvL����v�m���;�4����/�|ax����W�%�� ~�,�qd$�!
�R¬`���|n���'>
��4�䳪[��`���F|m�A�(�vX���W5���<3]d�L�E��2p�l���<�@/�y�/ �ƫ:2�P=�n~v�-�a(L�ޅێ�cT��y�ω����M)?Ey�ptw���uU'=Fխe���*]�]e.� N(��8���MQ�3�8����Խk��G�g0b���ѐ�.�N=��
w s76�w����&�a�"??��I�F�(kk\c��Y:������h�4��}�C��vq��"�s`��p�I+�Q��Q��_8��5�-Q>���Dޝ�@��ɕ���֟�K��4ďu�᧮SҠV�Ӡ����R���\�wC���|�d�[]����:�����6�\r��%���ep����D6��rƢ�P,�-�g�����x�X�l7����"�ƶ�v�"���8m�[��:��tr���Q��͢/�� �.z�H���찛0�����t�ٖ��Zp�����{ۃ�����+�2��p�Pb.Ҩ;~��'���ڊ������L'�;��1T�euT�>"��[�2�c�
���q�FF�l[ԉl/�3�q��U� 
���{�ѷ�P�����A�Q��S~Qߡc�;�s�C�$p��\f
7F�x��p-;�j�*�.�\[��"��'F��5,�r�E�`�������P�mw�T���F�g�f����*ʏ]3f�����P��W���>x<$�cp��t���gl�����j9���%�.5N��-��ȱ6�K#JY�Ⳝ�V��� M����"|���b�C���~e����^ڭwE��NZ'��8*�v���Z�:iA�M���K��ۡ=�������!���\t毻Q��ȯJ��a�G����zƙ�D��7�88��w����C�o�6�]��G�����1I� &�
Xn�<|�����A?��@{5��+����j(���x�T�K؍�����r���_מ<y��]��A�逎T�����t[[�hwn{���������
�j�_B�.�יY\m�|�7�F�2au�yŏ���%%�G%h��陇�������P���F�������D�_=i
��٪���ّ-�MLGF���*�̮���X�u�	��ȩN�#�>[���]+ۗ�1�N1�NO���Y�p�g�����8��2���4��"M�ǰ�S�A�(t�P)>��m�������vH�n��5p�����5���n{'T7w�"^���Թ[;����"��}�ᾆ�:JN�7�>�yJ3*6�~)��MPCK��Vb(�*LM��'���6C�E�N#�M��h4<c(gQcSE�@m#K?3wc�F��Yo�S4���[ �y%��~X�o��	�<CZ����<~A�A�k��8>I�m6�x8�A��(,��2�֥Q�<�*�\˭83.����pE�8��y�qoPq�S�dZ�ѽ8�XO����Ty��oC^qM^+[ª�@kY<����d����tyX��v)^ą�ltR�|�2 �Sdq|��R�U��\'���ʄͷ�Q���e���)�M��D�`|��h�Pg(
�3iS#�\ULL�0w|.t������l�q9��2��������Fh�]�4�܉�\�LwU��oy�6��b�P�T�]ˣ�Ɇ��q����Ŷ��B۰�]`�b74���*e�p��T��e���1?�jD���s#��,���B��?oͦpQca9S���M^7�����Y�K5:��e���ز��� �ȲP���E������A��1���/�լ��ʈZ��a\��.RG�15��	wω7p&]�Â�h��;��,x\��j�+������� ���TM�3�1���J�|C8��,) memz�I_��[v(5o2O�L��ȶJY��"r-a��1l�@#��݃0HO{�~��β�J/��9��`�էb�9�/_�h/�?o/^��Z+�ގ:��Mx޽}��ʖ�M��
�#m�ʬ�=pi����w:/֡����W7c�
�ߓ�`�<e���:Ix�^� K1�r��x��c�O��0���h���`���o�q�#�)���ȏ#�5�]�r8]ؑ-�\��)�1t��)�{G�g�CK�s�<�+���E��GR�R��#2�:�?�)}�i�N��F0c��^����v�DN9Z��#�����F�G<�ѯ���ACK�s4�YJe��O��{X�e��Qf��h-C��2rŽ���m :�������n��kp^�����K(C`e_p�:��w^;n+m�E/���4C�q��t}q�^ٖߏ��9\��m�z��[����廻��n/�eY$���؇��dy�?Ҽ
@�,�$t�9zu="/Tz����-�!]�UE�4�]8 �̸k�_��j�����_���y�ER0�$�픅ӡ� �`<��i�hH�����92��I 5}��k���3$|Q�(��
�^ȯ�ǯ��z(7���A���t����6���W����6��|��T=��i�t*U���9���h8�H���ʢ
��m `t�x%�ț�uV�06v���v�|��|�v<]#'��wmwg�����u��}
���x��|��V�t�G��n��������g��v��v�w����wӛWʌ�Fp#�F��� s���;n�����Fik#����9'=�0���}���;��04�G�MX�����M~* �h=�cg�[�G�4B�h�Q)q����\=�\��f��~��P���uIc�LO�wW"����U����mv�F��g6hHn�����O��	l�g�a&��!e��uK�5<�s+|#�����޼��.�t�xi:����|��ǁ�G.����3�}�/����T;*��+?�k�]�zK+Lߗ�ք'2h��2�o��0��RQ0[a�>�@N}�V�FSX�i�� ��)/i��]��w��P)ܩй��;4�5�����y��,����mZ�?7]��9��T����M�*.�ĘY����ww)�F7��Y_u��y�T�xO�=d}UބG�F$)���L���
?��R'��O'�҄�g1��%CJ�aǓӎ�:�G?��h�蔈{{G�ͻ���՛������٫�����������f{�f���m���u}�ny��ce�A�}�i���o�v2��Nm��n�S��,ƒ;NcNP��U�P�Q��Y�
:���<�mn��y(���q�C��S���n��ҕt:jo~��˧��븘l����G��u��+�t� �knf��)�Y��c=���
����%����q�NQ�YG����
Fm>8u{|G��T��5Хmy_ݢ�s�t;lepϟ��#�v��h�aSL�
<N}8K��AI|�<%$�HG�)��<�	�Oĕ���mul�$�g`il)c4�]��ٳ�C���7����ޣ$^bd���܌�e�)W ��'2цKX7~�*�� �rN!���V�ӂ��K��(唩�r�z���_�[��3Yb�vy�.q�:�M�Ͻ��d�/#�¹����y��٢�:HY�j�L:o൩Ye�4~&rbfa�M�-f���L�9h���eMç�x6�B�h+�լ-q]���4��Ye��Q$��9FPFI�{Hy�b�aT�X�o��k���G�F�W�㈕y�o�.>uJ�¯�cA��}�)��R4��C�}��t�s��K�Zq#����ᥑ�/����KLo��jR�&���w��p?t����z7����\�*9h-媲��:ߧ#eR]����o�l�����r*��3��7z�wy}��𾬼��K��h�!�P������_���/�������=y�m���]�Q:E�d$��1�^�:!��H��w\��R�nx���A�h���8a��2+�z��b�����l�o�Ziy�ҟ�K��G�V�k�0��1x��Eé�嶻�g����F�g�P1MS��"��h�4@%rG��]Oض7�p�j���q���i�N$j�zv\��
�#am��׉#Y"{Xʘ��� tE�iOs�@
OmS��ɹ&m�#�:��w\��Ȕ�`�N� �w<�ct��˧��$�ْ�2��Q��=¨Ұ<�~�]��y������N���k��h���TA�ǘߋ��4V���r�Q�0�W=�*��K�D�wۺr��}�N{�EW�5�j.�|�?{�y� �lI�F����;�Z;����(��׵qwE�H�h����B�B���6���~�w���,`���o�)���^z�Y��y`\�i�(q�c�|�^)`������IGA
�Wxs�p�����\��Kw����(C�6��kh���E�ėܩ�Jl`����K����5 +|d��&�RE� u�eeWon	ͣF:�!��H;�2e��E���nW��D��m��N�_Cq��g1�ڒ[�#�f10�ә~���*��Occ�4j�VS�IW}����u=�%��`B1|��^*ߢ}饛���?���Q�u$K%��k)]�z��Oe�D�ӻ0B<@tn	�
��]1!`T�kٖک����Hו6yX�F�퍾66C⨑F���tZ��ጝ���������Sm�99�h����9@�"�4�4���N�V�*4�q|�������(�n�}��� ���v�EG��Iе�oz�{h�р�� ��C]���+��wy�[&�օ�λܿ�Y�!r��W^zt��/T<�U�Tm*cO������&g2��Y+++˙
�z;lX�E��`f�w4���M;�EU>$���Ox䈆��%��.z�;ro�#��8�.k�[KZ򥾕������6�*ePf���k�e�2�Q^�%]�V��6�'� ln6a��wn��'�Hl:5���Tp�O}H���N���Uة�x�c�)�,4k���
c�W��z�/F|�p!ۨ%��9|�1Ky\\��8�)|��M� �O���oh�i�ś�J�X#�Z��-@+�w�ĸ����4��#�̩��C���B�];z���"ӄ_`�4Op�b��i�dV�����:�A�8����u�1$n$x�-��+&�q�z�ތs�{��>�:p򮌭�n�etRc�khY�����2wإ���V���CK��F5L�WȚ����{���n�X�m�|��Y�uw��i�Fpy_/�?8a��g:��{?-����4�����7ߥ3���*�^��g8�c��o����������u񳗛��.)�!�+2�ev��iF'�@�3�O�YyG�ԛ��i�TŔb�y��������l��u4�Tһ���
�ǳ�V <P�<�qJ�/+bWМ:�I41��'C��ݽ���y��m��=y�Ee�v��D(��oj�Z�B�k	��w8	�����*B�)M����e�a^ޏ��� �K!+�S�L�P1���FAE0�hкum]�y.�0MӖ	�&�lP$:�$�ދ*G~��K�z�T��A �ô���q�b��VF�lP�9������9�:=e
q)H��F{�r����&#;�A��]8욚�o߶7o<�ͩ����ꚤӳq��8��u�6]���!�s�r��0��i,�#�;p�wr�$�B#��fSsО[�����t:��%���AɈ���
Wo���i���pp!�\
���撄4e�8DmO�S���0MҨL�Ш8���(NM/�!��h8¨�N޳N��]wO��s~zz��i�+I2e"\Ѻ�cᄫ����H�*H}����H}2���4��
/��bt�뮩��Ё^~+�����|{��Kի�Y*���&�#e���,��U��v��Ͷ��E�z0�["�fk��ݞY�7��>L�Bt�䁴�w��>ߧ|�+������M�,d��9�l9l���R������<$��
9fꚖ�嵶�q�-�nP��o��b���c��`ǿ��<�:�G/t���^X����~�c�5��<�>��<�{#�����������}󢹥�9
��0�2PN�R�1�y��J
�%���9���ѡY�_��|�g�yX���휈��Ȣ{;u��ն�>׮gk�U�_�@��su�� _[����n$���u�`84�Tp��8����L'�p��q'5�I�;eh�5%3�/h�3�����+��Ս.Tg�mV�~>|�4ո�v�:��a�̌qAR`z��VWt�}��|z�:L5�%҂>a��3��p��R���^���݌Fjt%=ӗw�L;��͝�������}��!���|e�K���w��4�i"~|"pl���z@�-1��� ہ��G��`0`�OY2%��M[i��&�T����!<m�G�C�keNr�ܰ�xa~Z����>Q:vʿ�}��b}m-��We�F���޹�n���͛9��%��n��3��[[�ѧ�[LJj��ݪ'E��۲���S���1�o�������Ae$Y�Y܈7u?;�(Kխ2���ND��Ȼl�E���T�$���	�R��F�XYZjwo]own���GH������כ���뭌2� ��̴��vD���4�Evh��7�/�U��*8�s߷V��Đ�V�p��R��|�E�N�7���D^�$yi��7}��۸z��U_�&���M��ni���u v�Sqm��)�����I��I�ڦ�j�4*��h�b*���`�:� �|��G��x�r��p#c��T�<_���p��k���/{���H y��^닗�Q���$��n٤?��]�J�sfޝ�]f1�6F�8}��F�y�F[_]��'iîYo������	����I�xR��t���~'Hb+l�,�d�!G�P�!�_ˌ*�2�ƚ���0��1������.��x��5�F��59e���>:��J�vd;�st�r���}���q�w�5;N5��
 ��TF�/ї75���Cȹ����I.ɏ�|K|��R��(�F/F�r\y9\�;�Hp]�&>�`H�?���(�S��38�<��U)������1�������k�@�����B?ӽڣ����;�3�XeQ�*%���Rw*�
N�/�1��P<�,� k�� �,��e�Ɓ��9J�.�w�G�6�����[�ҵƃ�?�a|���;adm��<c��Q1�����߇��|.G�N��%�d(�|�H��� ]���c_#P��ʱ?���q�L����K^F���|P��J���� ����S<Ә9]�s�<�#�Cb�i<yࣾz�5
Q4	�i�n�c��l�a'��y(D"8S��%E�x�"̡q�<�y;PB��"%b}�>�(shFz�>���z����;kRa�j�R�"�訦F�v#��L�w�-�^h2Z�̩xp﷌��`:k+�˛��p|uEa�~�"a\O���k��͌t� �N�	���'��?���E���Z��\<e�:��C��)�ܬJ�|����V���<���IEMY�ڂ�I�\'���U��G�D��K���P��%�ux���\ç8���>w)�4D^f�F�O�?:p�%F���m����a�n����� g��x�!X�����TQw��|z`���/����
8WNȳs�mqq-��~C���v�ƭv�
��{�֝{��������n�^�n�	�����]�8[XZ��ښ\E�]�((F��:0�U��Yy:�!5=k'�YG�S{�]_��-,��(�SQ�]E��4����V8�p-�puUq�|����&.��z�����)�
*�|x��w�Wm��s��>x�\�Ϣ�n��v�����p뙀}��QÃu咴_y�f?*���Ȟ���]{���v��H�sڭ��gv�#����pV�
ra�6?���E/��S:�0�Ż����8z�5Mȟ����,�^lSm���rg#g��l�P�Cy'�bt�Q�G}��޽߈���ҨҸz��Q����dT��'r*x�C��=>���A�f ]� Mݐ�HN�����2�T�����Ω\`vj�r�8v4U�hd�zٙ��Cئ����t4^N��2�5�s����v����.@Gҿ��%(����ͻt�-�;�R�R��)����!}���]�Lҵ���Wy'����p�Ǣ��O��봮���Y�Sv���r����IOY*=�ҐN�+�ZI>?��5P����V��{Gz!%>�n9�\�S��p�)�NA����M;�u�2�>�dn}߿~��:������0��3���-~��䫔/_*���;�7� ?�xN��G�Q�:<��,���xFy�f��ϣtfB?�ಥ�zS�a�?�YO_�m�_m�m���6(�*�"O`Ul=�$F��4����KEt�$L�e+aY����O�^�Q\Y�ј_���bYp��j>n��������������ѓ(�O��l/߼lG0�����;W]D_Ui��!�m�?�Ⱥ �����59;�(�ɒM%Ɂĭ��"ˀ��|xg��R#+��}5x��IJ����ʗ�Jr��{᝛����g�Js���FE���k��(꒷�I�
�-�:���Gp���i�a� ��,b�/-��L��������V�I��B_�і��ڲ'��	������gQxHG�P��:0Te��)��aίA��eFzrҊ�2_���C��zh�g�!m%�Q�e7܎]�3��x8&��ã��x�v+B� �����y��0OBc��)�p��5�0����?7����=h#�X6��4�jX"�g\�*;�(��=�'�Ӕ�!�b�4>�˚����FF{����?E� ���� Ҽv�(e��^k4����EH�Fs�P&�Z��i�i��Q�\����<~��àݞ�w:�B�/�ݐ���_�y��x�$�҃�p�i�k�O	.�z�~�HϠ��>r����6��*���,z�DຎO�<�>�Z��gz� ��P�TpI�N�;� i9��~��ܸ}�ݹ{E�F�%9�%���x�����՛�c��R�B%D:L����B�v�(y�R��n>-��������J�S�g�-S��ȴ;+�m�o�(i㮱�zp���ru���j�s�f���'Rɨjh����Rz-�"��\@\��U�l�� ��e�3��(�*��{)\,�#�B,��'�1�3���wo���g�|o�M��	��q��F?J,��?���U��Yo������qۂO�0�U�<�{�d�G#hC���v�at��öz�N[Z��Q�%��ŕ�6�l���i��9��Ц���mBܵ��)����6�r��w�|fM�����7ﶍ[��ƍ�my�f�u�N��8RF8�f��s6���).hG���8����7�O��q��z ����@:���J�9`�*{t򐼦B���J�o�?��G|o�.]���28�]୴C}��Ç{mk���s�����n��z��dl�5�5NƯ9�+)���H<CQ�v���)j㼟!.t&_��D�yB ܺ��Q�e��J[hK�T�rz�F��IuNp�o��5�2m�B���v�)�<(�����CǇ\��/��-�,i���6[3v��y�ċ���Ў�)�ې?}�4#So^�l�{d㒀m�{pzq���M{��e���/�W_������Y�j���YF�qQ�1�)�(^�i䒀�3E�����dV�u�*O��q�F�������ǥS��>�"�wV:�.�v�m�m�-����^;Ǐc�+���i�[��n>�������yC��z:�au�6�v�+d��W���|���o)�>1��=W��6T�m�-'�G�X���Ë��z0@XhH:J<��0�0;�
^���&5�ɁV"7��L��.���֥.��i/�9�ʽU�چ�_���|��N�jE�<�B�:0Ե����,����4�l��.Ǩ�1a:�)��u�AޫÕqm{D��,\ʚx!P_�~{�*��<�ʻ�',?�ő�w�s�w�xupB���W'��IE��N���t� \C�PF�+"Tq*�#7��|�9@1��������(�-�[�hK�q��������?�n�=y��={�.lND��ȲV�@(�9p��ʝ#Y6��dY9U�18��	� ���<B%���]g�r�qQ*4�Hd�*]��E�o߼i�6o߽JźɅ�~����[�^p�#4$�ps`Q��@�~� F�=j;�\�Q�����z�>���!�z�[�����o0I�eX����>�zmK�^*'�gF����;�"P-O�X\�\T����C*I!�����^w�r1��W	�����myy���jX-~����Z]mk(5�K�W���_0.������J��9�5��6�گm�;6�!�����SO�.2y�G8�%�32q\�)��b��Cx�#�F'c*��t�E�bd�}��C����mD�E,kHL�c��c�*�)|5�ݪ�.P�il�4��(��e���tZ�l���N�]%�fy0��)c<��H�I>|�l ����Jq�u�/��.�;%8Bx�(�*�y'.b�&^5�YS_�ȼTRw���U�+'\.V_e���
��PaH�J��J/
�t �2��f��W����mw峷У2u8�w�a��9"�$[��x���v��W� �$\�?��������.���Hw�t����/jG�w�2ꙩ5X�4�TI�x�FQe^���[f�����9�l�99�i<������t[Aip!��rI7�٧�'�?����FD�7k&X2_���葯�8ɥ^�N8��������-y�Ԍq�_I�4�g��Q��7m�-�%���Oʬ�-�j���	���J�I��]c�c<ogo���97�XY[��qtJ�
#����7������kX�2
&;�IA� aZZ�UO}�C^�!��b�����f�a��B�[A^��9�г�j��ŅUd�Ӌ��.�ۘiU^�h�݉p|z��-̵d���Q��4GG��%��hP�7��,��S�.�!��*�?���/����KW\Z9����kh1޽h/_>���i�t���P��΃+��1�P`0�4��Z�X�E�5NN�AG�`�]��)ʥ��
� j��Cg��A��#2�}��*Xƃ�L��}o7x̣H�a򬲪���y���]��F���9e�|�;�._��l~�$w^��z�^a\�ƿ������?�}���p ���D��r[w;�i�҆|	��i�\��g�%��3��^w�}� 5��>ubg��f2�e���:$���#[���q7�R|��(��<H9b���:�ϝ>�\Ȇ&�M�[����v}c�}���v���ɬ��R��p��m?y֞�|��W�k�\[��[X͛_�H[泰�L�N���g�R�z�}1�u�:�=
�-U�ֳ���#�J���r>��e����x+��e��kn����]������͑�Q9�^m��#�x��u�'�C�g�����,.����?�z�����4�=7��w���\�gn�W^�W���G����*�S3Z�sҡ<�q�W��(sS����^��L���w����Y����e�@�^�	��x�FN�(V��i%M
d�x�p_P>�H����w������r4KEfA�����g9O�/���M{Ƴ�v����*_�UD�+�jyz	OB�o����\�p5���!_���˼#��+^zCno�=�~{�x����HOЅs1,��u� � a���n�w��Ƃ��԰�Y�;�~��@��;�c���߸��6P�W��*�V4�P"�=������������0�mG ��Z���(+Kd�P)��%��*}�ՠX���2��a�~�qt�����E�k���=7�p1,~��S�3�l?	]y&�[�bT��x>��щs�	��pTõ�*b��{���A e�:^=(a�VZ�U�W��i�8�.�k���Z��}���	Ң`Ԣ���߳5�S"�4~�0�ή���|�<�.�'�������s7��sP�Cb���G<�e����?p)�D}�W��5����0��h�ʍ�@T�(c:M��)��^mF�t%����~�?*��²�t���l��EƎ�cٸ��yk�� ����*��f�R`�$����� �ۖ�Q���&G��v�P#�-~��/�	�߱G,ds��ls|p@�"���L�Y�˷�`��T�U�7�k�K��y������V I	۸��ׅ���RE4��M?� A�a�H�|v�]�,G��M�hY��:�݇�~�|�i���΃��Ɲ{m���5��֦	;�Q��6���P�R�Ge��:	��[-#�I������P�:1�۹�j�͕1��tCK�:�q��A�s���'?k�������=��s`���qd��	wƝ�j�V+r*�P�ze�=ޒ(��$�8�h�Ƹ�<�i�u����j���p�]�U�w]xO��K#�x���cK~2|�#߉�wGw��M��0Ң�81q��'rN�쌝-T#��q�iOCFM��J'���U<
��zVgp���)��/�%*\~n}W8����k�囊l�Mǁ�}�N�c��m�hKK���]�*ۆb��i�/f���asw�~�ݷ�7���}���َٝhq{U)��"��E��RТy�Pe�r��C����4�[X���8�.�u"~v��GQ́�h���U���zȬI��;���r����tB �̴8�9zZ�瑻�O>ƹ��:t꿻uR���S�1ϱt�*�����*b�=>�?���Q d��vf��V���M%���2��eG�	�|�.@x�a�G���S�����UWq4OmK�;���h�=�H'ue�\q�ݲ�;�q=eK�q~��.s�{�QZ��ΈE��!�R��U:��`�g�������v��^8�M��q
-:V���_����Qxڐ��t6�p�,��|�S���/,��U7|>���?~|�����Rё�V�*��xGx6O!5\z鈗Q�S�܌�-�߾����S�G���O��ׯ�d݌��~yR ^��[�����r)I�W��f�8G�fѻ� 9�W�pQq��r���]O�V�cS4�Q-� �tlHI�+���.�����[��~�-�m�����.Z���
{
?�F}o�� �n,1kϩS
��]�T����ɩ6�-�η�9�5G�0�V�Zw}-S�s�,k�kZ�J��i�<;BQ�(�\_gcⴂ���T���i�&�cx�ц���=h`gg?~o��6��j�@a�z��t|���ܖa�X\�ZL]f�UwlT��a5�rr{�Y1�d�"���K�ݺ
�wW�7�x�sh�7ý��i(4����y��؎xl.²Q#C�r�O�1�Χ(�d�)�鉣�:-�rfwC�F]�P���QC`�-�49���N����e�'���),�F5\��(@�b~��@?�B��3%��r(�G>ǥ�������
͊����ȬiK�;�����"��-�O*4vDi�BRJW~��2��C�����b�L^����/G�	�1�n��y��cҷ��V7p�ΝbR�x���"��;�C�H���z�����}.��F�c�tz��8C����=�%�/9
���{^����L��Kv.9J��Lr����buz�Gz���m\o�>��}�����~�>�z�O��;�����6���!3�e�� vX��ï��ѹP�.Ȓn4��p�������.}�M�dN"���77��U��Q��g������>����އ�����x��AoS��8�6���f0�ww�}��M��ݎ�%�L��Ѥ���|zP�xѐ#�Z���*������j��?�Ǔdx9���w���#���4�(!��=�N#�K.g:Ʀt#�s��F6|��90�QP�r<���wҘ~��7�W#I�z}c)^ʐ�x�n��o�oyi=�u�}��k�� *k�|�ѳ���G���ӟ��=|���W���s�C�Z�h���#]�"��I\�Z-��ZZ�D�'��f�2�rmM��H�w�"Ũz���������� ��=>�م#���*���Y��f$F�-����9�v*9ҙͰ��%�EƑՄG# �G������킗w[���ֻ���C{��~v)%�d�<t�.��%T84�  ��IDATqlzn�_}�-�!?����w�IO�+p׶콽�tF9i���_����6<��X�O��9��!^��j'�0s%�ZrK�:ǩ�����e�t��⦾H�c�����U�ߣ���v��~,�{��X���W�$~�g���q�{_.�?�ų:�m���U�ը��ͦ����G�Q�<�Uz�ͨ|9I�*"@cjp�x�w�WE���p��]�h�?ËT�A��P��u:V���9�N-� b�ʠ"�-�3��}�=��Q��+{r�k�0�j)dEZ�*1t�vv�˫a�s���G9q9���_�7_G��#���v��m��4�ͨ� T*�J[ao/���.w��)�=p*��.��n�w�sʤʁ��MO׎U��A}���4<����Q;��S��5�4����W�2uqu��.��:�НH���9h��ϝ!s�(vm`�4F����rS7ژ�:3���nZ0I�'��1���|��C��r�=66�x ����F���J��``�4A��,�
:gݹ�2��G�
a|jp)�:�� (@׿*����ZN}Kb��f5FT�*o��Ե�#{�a���2��[�В�ar#O�����U�2e��X��?��pvV�h5H���%5�2]}��O9��J��eY.�v����,s�-�������[�o)#��IEhP�ڡ%{J퉌�BL�}�Gvx�R� 1�K�R���_e��.�#*41�xo�{{�;�>h/{���w�y[Nm�fʧQ��U�v�ቋ6��83��Pp����a?�a�*:3V>w����v��|��Q�
��?ěa�v��
�hT$
*A�k�нV��g&����(���y�_PQ�8����VF�Ww�;F�r
�S9U�����4=�˵US�?w��7�g�֝�W�ۭ{��Ï>n~�)F�G�ƝY���f � R���ȕ�����W���X�g�_��q�5�b\9�`xF��vyu����ep��N1d���/n����mf�f[�q�ݺ�1� ����� �u�ö܋kmc��}w���x��=�*�v*�`éG�R#�����Nc]#��aT;������3��u?r���]�@/?j�ȏ������@G��㧃�!�w
���G{��~�8��8ks�����|C巉����E��(T�t
�B��ŷ̊ ��:��'��r���5��_x�jq]�m\��w��1ʈ/ck�+<���ҾƠ�?x��}��'K�?D�l"��{X_|�Y��O�hc��v
캳LV����ǲ;�;��'�|�>�^�y#k�2H^�*p]��h�ޑ~��%�(Ep�b�/]}W��S��6�6z%��'��%�=�u��� n4J�ugGȵ�t,�i`q�Զ!��
����-�����.A-��X'�͛������������[����SE�D����i��`[^�t歄{yG�x_R�zU�UR��羦
*���5�2�ԫ�U�B�E��#�^G��&=p^�1̜�t��:J?^��W����.����M��:����/��r_�H�AO<��;fĝ���\eݐ}`�ƣ-]���7y�|n�H���8�yN�hp�VH#h��b��x����zA��D�)憋����5�H;|�?�����l�G��d�w����D������rõ2�BZ���(�FE�� ��Xgh���9�!�����L��.E���I�WG5�*Ѻ�K��t��U�-���t��� .ar�ӡTJ�ϲ��.
���k���U]��d�2EI����+��;7W�d�������Gޅ�(^1f�!i��y���:�m��v�2�[/vpF؃7^�q+�C��(d0�A�4~�W���:�*\�:&���}��(D��!+�Du�+��}�SOc�`
�嫸��)�H��lݚ�\5Ν'��E���
�5��~~��	
,i�A��aY����+����w͊�6i\x�50SO�M����� ��1��0؎ ��'d��	�y�sk��/��`���*lUvK�j�f��k݇�X�僐 �4�4�e�ԕ�>�|��.*xOh��\bD��lRC�i���]����b���<�@�~�Pa.��G�����Cۖ	�����t��U���ǹ�. wj�d6�pm�
�<�m�3��z���NM���a�������;
\�������q��.���L�y��eF����o �֙�G��{#Z��"��St���-Ͷ��X��ܺ�];;�����z7F�r&
0������bhR٩ˆ��o�)M4&�eX�U�z]��`�������0�H��YiC�)�ᆰ@���j1�4)���������������v��C�"�i7,�mnt��v�h\ihy���w۝�;�>l��=n)
���1�4���)�GXe>���-�pR��8��F�Ѱ¿�Q���ÔK���k�ِ��U?�S}O[�,��SVR��'x��Ņ��N���޼l���Y�j��4O�*x���-,䬌�Σ����6�XWe���P�mĽ7�2�2R|�'������������v��vU��o�d�%��J:�-�m�<�N�zv�#�%��iH��k�|�d�s+FEw0*ޭ��j�r��qy��\�o������I}�EB١ ����s�>���?F�,�P)��s���Hս���Q��w߷�������_��EF�n޺��uҞ�'���3u������숪����]d��G��H۔]:��5Y��;:�t����Кt;��1@S_�����U]�YH�߮Ê���B�Y�A��a�+ω�K�^�kT9�C=�"79��}��dbd��wn�����}�كv��z����1���n�����_~�~�������� ��-���A۶�3h /�b�^S��-�z�@�u(������B[��<�w�2#�ґ������b��6��4H���%ZCI}���W��L�c|��_�NL�d��U�5�l���q@��v��
Q�!�K�t1�I_/.�Q�<;	lk���h��W�ګ����9��\�&��VEn�Q��:��/�V���{G��Y�RM��e��ޚ����mai����Bn��=tD;�]7�17�⻼�QuP�����ǿ�sw`{��F��	id�<��K1�"�9Yx�y��5��ڧ���
=EPVl*&L
"��.�T!�bk/��ѵ� �J�kl�3����'De˳d�rP����찵��� H���.�&$.Eh�F��~�3�v��Y�X�`Y���������r	��%a��⨻0�_�^����C��4��a2Laj��r@�"9~
E��ŏ����0)�'}Q�h&$a���껼��#<�\�xI�^����W�#z�����?_���D����r^E � ;�5�0�|�T��R�]��1̢��[���Fɱ����Uc�ú��*l�X��}p:�1q]����`�C��OL���<\�C�@���@¼<8X�d$(����q����JU�B���D0<u��jgFz_)dM�{*��E<O�:�l8�ȟE�O�P*���+e��/ �{���������ˀ#wy_�*0t�R�������é.Yu4�yA:��S�B�0�F���i���N�4�6��k�t�2��tp ����\�\��skӨ�bT���s��7�_���=����f���==�M�2#�"?��R�hT!����c�g��/M�1�����c�XGm�r#"Q\�S���D.��<��
No��$Zq�8�<�_�2s�:a��\����X7��GO:|�l�R��~ޗ�!U��kf�f�v���W��K���Y���"�id����h^�T�=��39�j㺻��o�Z>O�.B3(r1�,������0*�0=��>��5�0����2�<Uf�,�.���Ub�_�*������4mO(�r��y_�Ig�J�#ȓ��:"C%I��N �er7B;y�P�b(Xf�xŢ�Z$���mX�Y����`���B��ߋ��
G�,TB���ݝ�(�/���+x�-b08�-�?�TF�AZRQ�'��5���Z�!�|p�^��?8rc�9|ސ�v|alEP��3��������L��t�+#݁Y��ȉ�>�V7 �*�7��/�`�0j`!�ҡb'��
���&�Q�l�
:�ϳ�T��~�o��ۓ��e}u�X�Ћ8s�����v���X�o�?9'���'Y��4�Uz�����N�s��`�˳��ұ0�Iͅ����%Ҭ���������*����-�Kg�Xnha��}ڰ3o��@n�%|k��o���u��fڽ�w��������(����5F��߿h_~�=��c�w��zlh�B��N�/� wS�����RՍX�@��/x�)�y�d�S�O�1����x��D�i%�KK�)�T<���Q)G���2��3���^#��*,u:�
��J����YR���I�i����_�9'�5�N�d�8l�ď��N�|�h��&��2s�=�r-Y��7d�+����^��0q�`��e�y�����+���M�,q�}}Ww�;�">'��r���������� �����t�{w���R=!=b������/�z����m�È���ҋ.�̊J�F�FS����@z�$��K�B�"S����L�C�]o,S�E O�
����?�p��^�8��i�햱k�򭶾����8ٓgx���D�1�#�lﹽ{� r��(b���j�:,]	.��s�=߹y�Ȫu�_.y.���U�;|��N|p�1\�%nƖA����I���=�2�:�+D�s:5b�����{)�~�@u����h�9��&$
`�N�3-�Y�`�@A�"�
f�hQ��2h<E/ՈV��H&�Ռ����\����g{z31�r�M5�S0�pQa�,���յF�7��V�X`TaQ�S����>�۴���X��k,���T<<ߦf�g$ht�h~��g,�Oy�p���'t�/��1螪}ӫ��S1����W�W|�6%�s��/|��IOw��4c���w�K�W�Y�h��*?����[/k�����H�Y�6ZY%��'ԩ(6BF�r����0���rZ��rgG�\�ptP��$)�l<�8��8����$�o��4C<GI=�hmu5�qT�����O0����Q�Ĩ�R�� �H+g�z@܈�7|����"�4��S�N��n˓mmq�-�Ҡ"��sW-�`<M*�\����\�(�x����&+�L}��ț����7���� ��p�UIܺ�5�t/6#ϹZz��*$�%Q�e�po��{��h(��oQL��o�e��!7����(���+���������{my�F��_�/g�چP�#�S~䎰��U@�E�Q"�L��ӓ�J���w�,�'$�ʫ׍��:<�2��x*��xGz)\�lGʫwٝ5��H���HE�xEM�r,c�n�!�'�5 �[]���s?��w��g]�J�����N��~Ӷ�^��rZ�2�Q�sq��t�(-��J��{)�v�z���'�,�}t�Q��S��xW�-��jsT���LV���P��V�p#��<UNX_I��@�e���}��a�
�h���YUg K������~�$�mw�?�?�6[�����)��{�i�t�.���n�r���[+��d6{��Q{��qvBu�e��4�	���;��vZ��]�F|�����Ա��;�Q'mKw�G,�vy��	:�9z���N��]hw��"ݞ���#�����K�iM�p����������{�?����=Hک����>������#y;Ќg˩ש��L�,(CKޢĔ�db�_n�⡰¢��h���6I�r�P��S0V[+R���M�2��A:���y�Ε��o�*�V�2�WF�	��(y��S#�<��,��ʔ�-5Hqgg�cػ�3BLKK#V��,f�Xm��@F����u��<[ש/�u7<��
���:���M��;x�����ܡ��@�߼NFḦޣ�\T{��0I�F��M��Ъ#9������M��t�ކ5���7\�P'���M#+#Y�1�<��	E�{YD��P�ޑ�o�tA�� ؅�O�~�0)\sߟ�����J���Y!V��#���Uo�I�C؄䡁e�ʰ�QV�r���׳����7P����>�	��g:"���5O�ߦ�[��mg�Z�?��,{�F��֍,�-dRB�5���檑c���Ί����ﵫ��䭟�gaW�fx�J�W�O���(����4B�R"��'^܋C�ʌ=Y��ѬA���rӮ�F`h����\ݥ��Iu��V{�)�V��W8	�� ��C�2c��*�5�<E&����UZr�@�~a~�-iPa�,h`���id�>��B\\��7{c���a�t�۱�9P�n䠢u~1�|}��;�1V��@!�	B��iP#����R�X#�`�	��I���T�XVY�Ey��Z���2�����z���C�+����OOd6��]��E؏���0��2���=�Vq�5�DHã��4p*���
��_�z�CW��gY���/̟Gmc-ߙ�q�(nM���W��d��4(����Э��]ҝH�R�ćN���:�� d�_y���1��,�t�����(�N�y��i�:��<�M��)�;�t�[���#y�W/e������t�bsm}q�-�S.���vz�Ă��*#+���ف�;��u�Q��;; l09 e�H��un/ݨ�.]x���է��5'>��*W����S�f쵽�����s�W�p�:E%F�N	Þ�)�xq�FsJ�����ZX�/�pq{�񴄤�ڤh���rk�Dq��FlV��G�Sq:�ɵ�yx֍��/��Η���l��r��t'��. w��uh(��`�N�WG�R��Pae���d�g0��ݦ=�B6;���C����i�os���vt{��K���P@��c\��i���k���eƨU;a�4��z���q�C��C�'�>���;5��ed���.���(w�qv�Ca�I;k9BɈ�e�uT���,%L�]+Y�g�K��v�?�t}�s�;�i�購!�ʹ����߼~���|��F�i<mom�;��C�� �ۣ�*��y���k�|�mF�mÝ�!�Y�~���*��˱�v��'���4�AN���x#��S� N���Y�
V/�'�s���EY��7,c��(q�T73q��8��C���n�������<�w�}��'���ն�<�v�5�[ۇ�����/ڳ���Ӹ�܍i4�\[)�A����2`���Sg�-H�<2)u���[*=hXe�ᣮˠ1��Ĥ?iJ2m�1�}����F�P�@NE�%�*%�$Z|^��d��#�齭�i�0�ŕ��[w�{��Ҳ�Б�m��G�	Io�Ȏ��.�l�Zm �B͹��&{�,<#��׳�q&�Bvw���[^����b�>(0�	>��j�A����mk�t`mH�,d����������M���lT�8�}�F�{�v�X[�D1���Y/�l^Yc�d �Dp	��F�h����]G�D,�FR����}1��x�qW�S"�<N�G�(�����W��@!׊V���<����j�~}�ݼ�$K��{*%��6�)����`DX�-����:��R�������x���2�pidU�r��kc���g7�$���_z����p��%��BOC:���I���q2�:bV���4�����(��ΎC�x~���޽�F��"��i�7�����Z�tp(�+���1���ᷞRvJ'��/�pB/G�{�S�(:���,w#�/̹+�|F쭳w��j37��m>ȡn�r�S���(7�r<� ���j��l�>G@TR��<>#X�Y1.��T�0+��X� ��H/��9W8[����w�\�y`���ױ���n��$ʬ�#J�H$G�ǣ��f; ��w�95��ۙoչ �5h�.�[Q�vǎm�
�����(q��ףXM��7q�S|��P��m�U�
@M�_�h��`0��턁r���,\�N��x�M�*�Jy�r�#���45M���_�_cLW?�*c��W)(�����GɚT���%8�MeC!4w�A�T��h�葳Y�Xըu	U���Me�aU�'u��:���x�.��¥^����f�ݝ�9�!�����L�ҭ�������;ajC�#�7�����miq�-N��IT��[r�Ǻ��-�o.3R�!��9�(�V))<�i�d�$�������LڢS���m�C���W5c���K�U�
���d�&~v|��w�
���.msF�J����v�L���"�����mq����'�VJ�N�΍Q#辰�nj�~�)�~��)b��Ifzkm����Jo���v�6�i�7t���yR:���wڋ����˨��)#峭�����4���#�Y=޹$VW������n{��U{��U�e�ʚK3ؖ�U�n�����}��I;�>�a�ussM۟�dy�N;?;L?P�2�
N�Nw+�UZS��ヤW0�O�w,�.�ٻ��  `tp���e��w2�^#q��	�f&C<��e�����qxY-3��e�\�-�m�l��a�	%�Q���9ҧ�^Nk> %o/@��r�hX����
����G�ly)�>
�����y�&@�`}��/۳�O�Y����GWoxR�i�6ү,{��o��ԡ�[�Ħ���e�y]�F�3A���q�`9�%�U�S�*��r&�TP�_�w�=���tV�.N�\YPE�UL[[�������R�&Fiڑvpt�^��mϞ�i�^�k�G���y��hG/T,;Q�Q!]����mS �?�Vy��սlOgs��k�E[���=��N���E�q?τm`_%7��k��\�#��i�,q��J+�]�]��Y�*�V<ҹ�<��}�C�zp�a���h�ŷ��^�K��7����C�*��O3,_���z�Y�_c+d�z�L�������Z_�	�~�*�c�z�b|�<w�&��p�]���8�A�Q�&}�V�.�A�'p����N�#��hӓ=���
JVs/50��_���^�F����|���s%�a���Rnj��8 ��ܷr|�Ř 7^�nx;u �`c��F+�׌� L����� �B����$���:f�+-7?�Xmm������e��iײ�BI�O�pc��ݐ ��9]@̼��Ģ�KDj��ųؚ)�S���:]u0���¦���	XNBf�
�"�D-_��7Ó�#"9!q�:� ��G'Z��=�._�D-�+ґ${V�$P^���D�VY�� �K2����}xt��!ԇ9��ݻ}H�e���
؎��!a���r$��,�*8Zf�\¹��N�:*y
/֟��� R�S�Y	-�v��{�fg�9Xlk�뙾��[F�BaF�rI�#�rg��Q��r�	Kۨ�y��.q<�a�׵{�.' �n�d��J"�uqZJ���:�>"�'Zި�O��,�B��t�Q��9�G�P�:�OK{XW@�f�ZF&ൂ���U��Vݾ.^y�K�g�	�������۾&�%@lօ;��Nz��_�H��U�e��WJ�?���#(�S~�����K9}��5`�c���!���[^|�~Mdu��(}�}x�ɛ�ӎ�n�>1=�;�.�^CG�7�%5�<�z��hn.N�O�s��
�xb�x��^���兲�cgs���ڻ�}�=�a!N��ٔ�_�dMLg(_�Ķ&�(x?2L�/���man�m�-��9�J��Y�q���5F� �B��R��f�Ą�{G�et�[f2�^6l)%8�Y�e�,�i�x(�M��_<=)]����l�DT��R�e�
��3���2"85����vs~��Q�޽~����T~�d���,�ɥ�s+me�A{��{mq�Q�_jC��짠�I����0�� �Q&G�UT���L2�Fr�ρ:m��2��`U�R�l1hӷ�w�~�Ͽå�8}���۞�O)2x�~�Re�08�ʠ�����JHf7N�o��㣜ty?<@X�N�dϺgu��y5 Yy���_���{��>4�:��Y�z򯏭_��{]P�C��7�q{�vv_�\���ACi�h��:�oHq?&4>�1���w�R�v�w��ʲ?�/.Nr����>*�dǙe�ە���6�@%��I��K��yK+RW<�wy���Q��/�Z[P!ܥ��x�_ɻ�4�#ǧ�&�s�9}�P��9*���1��
�m�+�,L���O��y�޾~�^<ڞ?��橄��7
y蘃V.Ǉ��-x�7U�
�K�a����ʒ}�3�;�J�;0������,�p'+U�QgD|]RN"\E��QT�k.���<����b�s�!�CF�JhJpD���05�i/P������V���|���Z�<�Cm��)��A{�z���/n�Y��\x"�P,�I)$��0�0-=�����:�mΙHK��Q�R���=��7���vO�7���Dz*���B��\nS�q&�� ��Z�|ܽ����(��笙K��=O78����_x`��U��9� �����{����e�'/�6 ��aF�6�H�4U�	_P�A�S���QT�O5G}�-��H� ��O����^���+�<c�R;�OT��k��w�#gԒ{c���4]��"56�Y���2��7�߆���I�e�{(�0�w�?���ե%t���;??C�B�љB�
��<�����~�O�V�t����4zqAl��${d�/£�"d�W"fX�4�Dւ�>��OFX��$���� ����܁��`�I�����n��/�{�߯����>Xy��pz����Wl~�L9"���5��r�2ӘJb �T+]Kr�bMW"�@�+���(\�����OB�vQ������;�#��6�v s<j�(_*`{�._���<�a�Q��w�������E��m��:�s"R��g�������\�_�7ć��A4����	�g���,R�)e�*�BbW���q�W<;S�$h��+�ClL$݌l8z��dү�^[흶
���w>��M{��_Ol���>�d��3��z��
����c��i�$b:]b!bb�[���џ��+ߪ���>4�1L�v%xk��$�Ѓ�Y�F�j��X�2���;����{p?��Q���ˊ?������c�9☰�U�����Y3�'/�ב��r�y�m=��Q�h�D<�	�tI���<My��3Q�,�'j�w�����&�����ni�z�_nx��e{��ut��.a����'s�����?�N��V�f��e��n~J��zQ��t�rJ��S�*�5����;�ȫ������#D"\y��ji�3of�q�Qۼ���/odi�����t���.�^Q(��K��[C���%^e|�k�>��|�~h��7&�+�zT�nDyusV��.�͟�r��se�-/��ٙ���~Fd _<ms:��Y���$~'�;Ęn��]e	��q?}�W�QHZ{v�Eڧ��.7o=��2K�\f7�V)�|�ï:a����Ƿ1��C��S���*h��Y���y�d�����GB+L�Bj�m=˿_y�+����~���~ݤ�.u�@��^7��Q{��!�2���:��Q��y�iۖ���9��Aȵյ����ʖS��|g�=��NmVѓ�L&��o6�6��a�w���O���%��r�G��¨R�p���`]��m�`�Up'��A>�n��ɣU<��U7��$���B�k�/����/�
|B�|���5t�K�=IU\��|���[\ms�
ӣ��N�L�7Jv0=� �>]�*���'t�մo�-*rgA��Q����@z��S��
�N� 0�Ȼ�G��<�G�Q�qŁ�ce#�)+G��o��k����AP�.�Q�:q�*!�`���rr��<M��%̴T���C>*��x����Z��k�ٓ�[-������r�/P�u��y�[���-��7���6o��=0���k
'z�ŉ���>x���<�������*?�9�s}G�v��Kii`�`��ZZ����\a��k����<�/�տ��W��^�k/ߠ�;��%O�06z���I�B�Qe9�0�4�D����p�5��	7�0bC�F���o�;���2��&�@P��9׋f�?�+��I����J���\�92`�JQ�5Z�hXJ]�5D�S�\.x�����Y����N�S�X�S!4ZuWӬ�(��ٗ��g�c�����>�#F�S�Ѵ��gm!�^�p�R0���(u�fqOڱ��"S��CйH<��Ҕ51�A;���+��H��'��8]��K7�g�*K�TX�|s_@����Y!ʣ��F@�2]i�l2�c�)��b��s\6B�,�,��B�:�֓���e#=`KL<㦊�1}�7�7g�N��{��]v�~2�Z��2�LP��LV�rN�l����Q~�@m�u�m-���u�R���LS�sqX|�i耖2Kq�}���#��z��u���&�r�_�"nߗL��R)ui&������ix���;�E�O7A>4��w���bwO���&���0}z�P���R�d�Wf�,֔��
��B���t��QX"qGLk�'�AN%:�$=��#�&.����4~sًiz�����Ks�'�4����^{��M���%]��΄K �W��9
�;�±�������k���8?Ֆ���uEP�/3�T������*hK��޺�+�/�Ii�-_���!�����>�fq
��ӵK�O�I�Z��z���x���"�d���RWg���]��no3�2���9�G�:Jtfrie�m�\m���-�n�Q��^�l�k�͡�����H����vſc�� "�W�i~���"&ƯĊ�lG��v�����=5.#3��
gf2���������;�^	**�Bo�KFw̷��)aK��˪�:�ү�}��)��T�}���y���77~a�. �\2�R8+�g9���|����#{(b]���M�ǯ���P;9��{?��(����
� >�SKl�\�T�QQ^��/���GaD?��<74Fz���Gy,~�{E���qx��m�Q��{(:[��Q�<�}�;�_Aף�=�]�h�vT9[_['�V����Ͷ]Zvڔ�IO%�i蚆ߥ_ƹw�^�޾�=��}��'E�<� -�?[�'픎b������0�o�i�(
����b}Q��?�n��̏o�K�1�
�=�����S.�+�K����US�_*9/�/ ��`�{����a{��u{��eہVG��>⦴�-�,�;�fȑD#1���������C(+����[:?n�g����֕9�S)�h}���j���7O�U���S�����UW���_d�Vpo]�ϭZ��!�p���Q�錯qTv3�H=l?��6��,�s���0�O�קg^�L�Չ0�-8N[d@�Ft���;L��m�kf��+ۻl"
v�1�����V�
w7DL<��SiT��ٸ|��]Q0|�.�P�BB�|��F�'��)9�{N*�)#{5D.��O<������m����/2���F���Z�>{��^�l����� C4K�P.��)�JV	��=Ha;��RS���A�g2�3���h��vl�f$i����X9 �۽`����y:��ʽXވ����/&��X�\�xp�d��ߓ��up�WɺF�h
Ht�R��Ni]�� ���Ue��ړ� �G����"c>&���0�|I����HB�<+dEh7/:`�(Ȝ<*TEK%�N�h.��� �%ZI�KW���Hk��W�B�:��K^r���� ��eNuh��xB���{"<�W|sͷqLG���SB,�_�M��`�i�<5�Tkm���1Z?a%V�@�^巃�l�ˋ8�����㺔��D�(G|\&hy�_��2���̻4"����!�*Xl]�ggT���.�2�a)]������c��M��MQm�O3x�&�{$��0��}`*�Z�R�B�Sޒm���{|/k��wM��>Ĥ~�������=Z>�Hy�q����ζ1�*Қz�����w��K�>QJ��sQ�dVtp�t�X4��J��	f�d�|r!"
~^:&W����O�)����*��(Y{{�{fg�yȤ-?5�5�B���W�"q�tGpʲS��k����N��-δ����4� ߩO�I���Kc6´Hĺ���~.|�'�	l�Zª�kcĵ,·ڸ�0��Z�����)���G����-\Fj�����:Mn�Uf�NO�i#g1����l�}REam}�m?��m���-��k�3K�Be�־��Y�^�
�H��i��Bv~�����܅�o�\;�箼e�g��ђ���~Y"�2 :�;0t�3mye^x�-AK�f��i��}'?�`��n��o��fSe�ME{W���JsD�����z�޼~�N���o�	��{��G�������৸K���d�*��t٩�O��O���C��
J��AB�����O�F��	#ϡ��o[[��;ߥ��H�Yf!MR� =�-���C��n�k�����O?B���l�o�Qz�5�۾��B�^�Н�� �a�q�o�?�R��G�I���6w��9�k�~���Խ{�!�c*g�>�����'��������G�'��X��`���:��̓�ۈ�3�G�/OBQ� �8��M�t +�G'�}�eW��L�)YE�_���
��zLL�U.�+s��'!���˹'ka�\ADl;�P�P���l�v�FƬ�%�@��W�T*�N*6*��o�f���U���T��2H���G�����@��2=�G��L���:�S�\��l��HY���]�����%����]�P��,+2N�#]@6
<�~17?�����Oc�Bcs:�몌�ͭ���;�LO�O88pzz���'��ԓ�Ѷ��\
����c�����6-���Mx�3q�U<M�F<��{o�~]>�%�|K��V�q}���A� )������5�s� |�K�y!?hm�`�ॺAn�&����N}��m����Nɺ�K�NU�^�Q�d`$eǑ8Q� 6_H�(�3Y%4��#��:�;�i^G��PQ ��j�
D�?Lӌ1�7���KAgg3ra^.-���_J�DGb���AbKgZ
<v��Ʒ��v&%�v&��#���%�(�8��ӎ@k9uSO��!�ޤ�WB�i��y�ȉ\�9`�T�p
R�g ��ˤ����� ٭{~Q���_	�N!������{e�o"K��PuZ^�y�9y�UB�)����3���!��/G���0�4�2�N���A��������<QP�ʣ��#Ўg\<�HW���t���p̲�9LB�����D�T��q����#�S4�3g�b}/Ƣu�K|�t*g�\��:��1�3��awo�wV�d���Hǋ�+��JV���e�7�M?a�s���F��&�cӮi ^y.�!��5��4�b_����I���2&F����5a�s8�\���X�mcϫ�~��{ؖ�ֻ0��XO�]r� ����%sc0ZQ �~�T�7�Eɂ�m�P���a��d�7ΐg)y�K����ʇ�>�,G"K{d�G�rG֫W0�w�2�k��������*X����.K���1�E7�O���8�z�ٶ�0[�^ ���âdQ!�Z	��.�r�xc?���ܩ䠈�O�d��<���]fb��l�G�(����c���U+U��ߥ�abX�SG|�i��+���'=/���[&���woP�N�0^��n�|������mikj����4��=�6,�q���fr�
��0�1T�Jt��:�ߗ�N�[M������1}��rY�J潎��*�Pw�vw�禢������C�Zj㝂e~����>u�������l�O�*��|�x�7q̯�R��kϋ��Ľ�<�_;������������4�N�v[��-~���۶�F�i'��#���./T�6���v}!&�7KqS�p6X��>\�0I��`��V!:3^�3��eπ
m:�����H[\�C��h�|�%��)[��+뛙IX�\ok؍R�����c*2��(d�Z�M���1������ %�!��KU���}���V�G��b��Ҷ����#i���Y���v�@��9�0�N �:Kۄ���_�!���
7ɑ
V���d�]�N+��jFC��&����g���+�^���
�ɩ� ,�0�*X��:=3�>ޤ�mie>x����s�^���@T�.�9��rYNZ�t�0ȋ���u��BQ�O9�_*XC�**H
�|U<9�:�%�յBQ��c(6��"F��'b�d��;�bY�x�0E���Ҡ`#ܢd��@�y�o�]���&������p���\&��5����,��qԮΎ,L�*GE����Μ�'���
����vp����(�KT�Ϩ`Y1�Eᄼۗ��۵{�#X�o�y�I�ʻ������[lf���w�� ��?h�����_�]�3j�@x���
����"��J�;�W�qRמ��а� �!��'φX]qE�6J�F����3c����_�o����r��C4j��1����C�3��;(Y=8�J�̂e3.
B���]A�����anHB��@�%�(f�S3�B���N]v�Itn6s��ʖڹ�4 !@޿%Db*��NɢO��J���{�$.v���
��? (��T}���s	ߒ/�z���[�^������D������PH��%�#�,q���Ze��)�UQ�A|��5M^S,-j��
Pi�]x�D�=a|�7�Z�9��w��X�8*:��:*�8���q)���K9��t��e.��V�"0̫�FW��'
"q��raYd��VxF��Q�*Z��xx܎O��:E��jO�^%�����wf�<�½ c(���R���ɮ��`������۔��V-_��i檫σ����I������^���l�X�.����˴���{�I��W����[;x��e~e�ʿ�ݴՐWe��@��A?�K��/���L�������94pu�Q����)Pa�"���v��1⎩���0�ٙ3\��y(�)�����~ƣ��`���.������a�	��������i�\h�T��(��!)_��m�i�2M�
#���ё�631Җ槢d-���`�Tg� jO�L�����\��%���#8����7$u���wyeI0��E���J�7�D�N�C�);�h����ǂ��Pa:U6��9�[��x��!Ԝ����ɗ����{@������at���ǟ~�=��{miu��NΓ�D调~����RA[
�~��>�P#lw8E=��������2��'�w�Τ߉ ��.�D�oB־�W�z�@���^����vN��ia~����3��>����R>��k����M�+L�h՟�	� ��KE��=q��y��e[lr�;�<�ަ�~���E�*�h�y6X͢�d]���EW]�7gf����9�W͐�Pҷ�)��w��Ƣ@_�����	���rAK!�U$����^'㩡�^�?z����#y�{���fg� 
iM���,.,e)��B�]v	�{���<iR�w�1����"����Q�����h�4p���s�R|�A�p: ���d�Hz� zD�N{�"�_ZU�ͷ��5���`U�T�Ɋ!ܤ��Ƈ��<k�T�;�^�,��k�LP���U���禨̩\ -R���s�ˏQWQ����>>�ho޼�f�n��7�\877]_�.������<���3X��q����Qk�FPV�Z^�n�o���C�{봩�#i�E�͓��kЀ|�Qb�g����1�V�w&��{ѧ�W!r�}V���߫ +y���Zi�{�,�C��Qؿ���Ľw����b8��EX��~�+ҝp���<t£�=��af=�I��̖ף�=h�˻w�#4��6��=��~ܠ-hC�+���~�7�.&oXc�|7�A8���}R��@�0�4�A����+\�qŽ����盳X���V-�����Bu�y�tE�||qIa7��א��,-�F��d��=�����f�2�Rip
�+Yޑ5%b7P�
�2�{Y�D�"��R��q��T�\t%H��2�D����$��)b	�B@?zquMg@�ZX�o� ���f[[[Ɍ����^{tvl��r&�%�
�"����%�V�����z鉎0�HD���g��<]����g!�������:Bb�ʕ��ǷdG�j�A�:}�y�K�,l��W�88�Vǖ�U&35�i�M�v�J�}W���o^Ͼ-��(`��%6�(w�^�K�03ӗ�!�T�I���kZ�8	�����2\x����])Y�u��I�-�	�3[�},�'N�N�������`��RA�p$�%�W޽����4���������^�0L�m���_׶2��'�����3ɳ�!��ZW�֯����"��e�.	��t�e=����Y�A~�&�q{c�����ܥI���aSK7T�J���*) ��������W9LHEIa'�=�*әɂ�X ˩Pz�e� �����ʇ���
'^l���U�f%n*ԩ<�=}�M.
u�Oޒ��N&?ae�*�"�B�z*h8Z�R��鱶���87	��i���r�2#��4�_��`O�������tap����<�����2aa=s������F��Gy��)da��M�!�w�
�
 ��)��!��ŵ��Ҧ�J��/�}	�~�O�5mt�)���\�������wۣ����7i�iJ�@�R��i)���W�Xe�����30����~�OS��[��R���e��h��x��(v�`�l+��pf�Ã��Km�*��=�q6=av7�$������ٸ����3���>("h�L�
|x��y{��v���]_�L���]z�� ٗ�o9֥�Y	��r97�^K��U���c ��s�A��*L���~���.}�5JF(z��l��~a�6@WV�ؾ��E蕬�Y�U�Y�����ݔ��k)�'Ε_][�����=˴�Q
IC���5r����NA��HA�ԍrG� �U�ʻ�����w�C��yL8��Ŀ��Dq˄��/�Ox�	�� +Z�f_W�l5��Ds���K��r��N�MƀJ�4�4 ����ce�1`����>��پ5�RhuwE�����'�y"���2aTv�Ǐ�,m������,4�l�К��h�K3(OS(.����J�����O����q��w�O?�~��=r��6�bc���.�U��������{�y����e���+��5����2Q�����F��A	tu�4
�3M��Ӌ(gK|_��ѣ�?�~��O�~�G?n���w�ý,7uCE�=~�����⽼�Զ��2{��%��>����l�����~t��)߾{�vQ����۶�r]i�5��O�����S_i|������חp4�1�$�.M�|�{�IӇ7���'��Ɂ�y���Ꟶ)�9Q��F^22�tk*����~d�]��8�ׯ�ˊ%�����(����P�6���?�^���Bi��%�3Yo\.��,�Wg� HQ��+�X��d�X?��'0��dYx�`�4�V\ �4�]S�
�dM���7<�Wcn>#}5f�HOL��V�N!"O�w爘N���N�9+�P��e�͚d��|���X��zp��ux���պ].(�U�*D�`���HT�/���<tt�{���������	��tJ��v��mf21������@�n��ݯ����XmHgW$�5B^%K�UT�A�)�aL�aU�F@�\��!�t`�ĕhz�E�##(>x:f���o��B_1�����Na�%,�Y�jG.A�\��1�$k}�I`e��'(Ϲ\���yr�'/e�Ru��f ��,G��X����y�f�\��i�t�"B>�{%���w������f�^ԯ{L;�K=����?L૵m�ug�o���n9�3�"z�i����|�MA�w��Q`����燦�'�/G��������Q54�%��CF����;y��j���Փ��H�����J���2�d�B�e�߃��f��C�P���\ �������8b�h�gOړ'O��W/s����0<�O���V�x��:��_\w�Jf��MN����,�EB�C���d934�R�@B��;� ��3\��~#,�_�ղh�� v�]�ę��aҰ)ܫ�Θ6�
�ǰe�X�D�,ɇ����zAd��z����+�(��2���d�2@<�v�2U-�����?����'�i+��tf�W�-�[	Z��
�4NĞ�m)�<��C��]{���ml�o3��m	~Cy�$M��ԕ?d�6s����|,,G �rP`����Hb�7�����o6�~��*��?�-�\��<?�i�Ϟ~�^�|�������9��A���f�`���kh�}���K�lR����Vr����Z��|Jس3���Q�
�.��?��	��_�la�˙ES~��	By�]#푾.?"Q��B�ַr/(��]�P����iٕv��6B����P�#�e���� -6��f��S{���*�� �3��<@��R�Β)��yw�����^��Ʉ�
�TO�+.�ȒC�I�+Z����!�TfU��_�`B.���w�:�`:�����v�NE��8ٖ��=��O�a����(��Y�%�Q�F�ؚW�8�����{��ݯv���Ї����ڦg��##ȏȓ�(Û�k(4�Q���ݏb?��~u����E��\Xg1=D!��g����}����q�����p�'�
�}��x����3Q+k+(V+Q�<��JZ���;� =�^~�E����滲�'3{o�'�.,����0݊��{�<P��(�IM�e���b��,�E��]��xᩯ�N�J>�t�8�\�@��(X�Vg
S
��=؅�s�-q�*���~q�I��[o����nq���Jl�$�_)��{��r��{��#T�@RD֒�x��,g��h�X��v�����"k�.������6zs�F���d�3Yov��A-�$�,1�aA�.��/ۉ�0@h�,`��a�#h(�� B�p�C$�'g'��4�!04I	P�HqI/#�����<��\��0��u��B�r����v�d�Z�~
[�PJ�M-<Tk����J�nM9�M��QZ�lc�k�V�'�PW �		����o ���2� �c�D���fy�
c���/>���b�DX�:�3���Z^Gp�(�B��i�z��IL҈HL ��4�׭� #4-GK�A�Y΁�hD`H��U��~֣]�(���d�+�--�0��Xf��/3��P<QQ��^��¾��m^��RS����)��5tI���B,�(xC���i:�U�?e��W!IԵf/��J��L�\p������F�Z�Իi�n}������A��o	���������\�w�RY�f�%L�c��O���m��(}��6$љ��Y�`1��ͤA$��x��6t�-i��&�ry~L�:z�]@�Q�<��Y��Sg*���E��刲x���#nk����&8�`]lH�b~Μ/..E�r����2�{�6}>��y�|�^\>��a� �M�z:s��Z!�B��P�96VvL%�٬	��Ge��*ʈ�<��d>u��i�H��@8�Kr�-���x]�V���\J;��΂��f�\����~D�!Ţ9
���v�;���=䌂ʛK4����N�}���}�M8��}M>�mve�N�݇�DyߖVڃ�?o�>�N��z�F&h�R��p([ʣ��+Y�=���2�}�l������X-p�;mW��9�Z�
]�;1���ԅ�n;��e�.s��7�f�#��?[���;�6�[����l�3�O�X�v�+���ଷI�+*X{��+��'�|�vw^�����dA�����%���g�`	���:xWKt������d��C��u/�|���V�_�zdg���p�����?4���y���pES�!9܀���#�L ��<��N.���uJ��kF\�J�R���H�����5G�­	��ʬ<e���,J�/�����z����8|l�$߼���[d�W/r�������%�PMҵ�W��K��G~.�~��f���S}7߰���C�"���W�2�����˃�D�lk����e����WG*�u��{�֐�T�~�	Y@�R�R>r�a��1�3M8g��m���D����V�2���<%�٣�%�����1
ѣG�(4��S��?q��K��t΢�Ͷ����ų�8y���{�y��}����G@��B����y:�3Xmg�Ӱ=!ғ$P��3a`�:��q*��?VI{�&(xpBT��f��S�QI�.�$�u�E�_��<G��1���������u�Z�����W����w%�`O%��>W���,��R�ݐ|�[��y�� _����ޝ����5_x�@���0��/Qz7O�&�KSy�����c5��<�e��]��S�R�\�:pE2N�v8��+k\򼶲�D�By]�Eƾ��d���/w�\p��!f&���BQ�y!G�{��d_.�P�)�������.]ɚZG��}f��cT�Ѥ /�X�8�q��͞�/�s�h�N�������w�W�(1.�k����v;��u�=�rAg�r2a2�%���q��UV��!��n!E���K	p�7�3@=�H]�a|�[!��2�k[�d%|Ӥ�wg���e��6�l�Y&��hRʎ�"�.fKz�����[l~!���;��V&���B�$!�P��DȜg�H{ɞ*�շ�ئ.��~bT�Y1�~6���K�j[��H�3�#(��;9�m�c���d&��� ����:3v�LA�Q��iO�ry��ݓ�j+
VXz1g���ő��j�� C�Q�j�b�bBwM��`^�$N=��j���=��*#L�O��[����c@�ͣ�40����aꑼ�E�nX��Ԡ>�i�o���O��E��"�'n�Ѧ*=�����Jn��p����3(@�t^���N%���ER;.gu��
���� N�J!�A1*�*Ys��0�����<M���g��ӧ�5ω���i`��c�#�T����+�*%˓�܋239��1֦�xy??=��^Fy���-�SЫ#\�%� ����0���d�?4�7˗����6�^����+`S���0%�ɥ�0��=�W(��6�0W(��g��M��;������'��ӯ����=��S�:��S�����<x�m�Y[ۺO�["OͳN.�P�W�����D0��+@*����x`��C���~?���o7U>��WU5��G��|���N�������r*���#C�]�{���z�K���pwMo̐����&���N�B�&'G{�����o�_���]�愠���Rރ�J���d����6��`���D�,�
��Q��&�3&�pA�3x��X���"ցNQ� �W����3�=�6BKᬉ�Y��YTs�֦/�7������V���wg����U�Zn���sƕq��iV���[��׬��z�U���	�)C�Ѹ�g�h����>�z)?a�c�HZF�*��:x��իv��x	�}�M��2e�>���Ӵ�S�<Q�C�Ci�f��Jds�4��gy/i�R��_�<���}h~�,,4O��y]��S�tҋ���7�ǟ>n�����,ҡ�� �ř�Qh���B[_F1Z�Ef��1�"D����6�_Di�B�@r	��&vK�l���K�G�9���Z%zjj,{�T�VQ�6i���,M"�N'm�c͢��}�fjf&���Ч��\O>���Le,K
7����ʠW�,G�zx��_�(�8���ԑ|T=R|�˚�%�8�5ܵ������� g�����C�ߢ`��{%K� ���"�Sa��$�2q����?6��X_���7�q�����J��1�|o`+n}�_|W��v��>�;��M�6��.�d]:�V�q`~�앴(#w�7P�F�ۺ�ݷ����4%K�9�?{���d�x�^�ڍ�H�1%-��3:ͤ�%D|:� ��rA�{�����}��#�R��E����GK ��Y��!(dT�J�@�w㹄������IB���i`kb../�I��% �D���P  �H`TҤ��b�;����Al޷S�H��aݮAl=��1����<�SƮ�wt����3I0(��!��q!dWC�@��/#Y��Y�A���<��  ����ڬ�3�A�a��pW EY���l4�̀�F$���BU�Q~�',
F��v�X����b{C�a)ʨ j6.S�
G��%��]���x�H�A4O¼��@.ݏ23A��!$�P�so��"]{Ӷ��v��1��Z1�b$,O`Z���m�~x���yD#DB�Sa��0�||j�Yj��ޱ��&'y��ύ���K�"��p���������N��X}��F뗻�(]&G{�w*Nt-!��jZ�Ho�y�������/y�&J�i�ZU�����7��' �f�쿝��Ym�w����Kб~�uL��-��*�i1��f��N�F}��X�g��;Ȓ�8�I�h7�B���{~n!�M2xw8�}d
^�d�����["_q�&aE}�r����IO�`L����Q&^!��/���7�ٌm���081��'M*d�I]�H-s�_ӟ�my�zL�'�i�8=���a��e�����\9��/��d�8�B��-m��FǉJ5�H�w�}��=*Y����^��d��~�޼l��^����v,c�O��A�k�Q������n;=�){��"������}��gl�l�_��<�'2cm	��/,������eim�=��;���|��}ʁ�\��F���Cπ����4������V��Y���g����B��6+��٥�'�{a�QH�L?}�x��>t�M0ٞ�BR'�"`�tS�	�]�_K-o�H]qT^ �0�)O��
V?���W|6O5t_��p�W�޾@�/Ώ�/;�͋'�
֛W���J7x5t}��h7(���'�ÔG�G\"���L@�5>I{�K�V�p�]��Z�o�0哧�e`���Q�/���Q(�.m����O::JV39�	�C�5�l�*}��*[��v��X``��4KA�\AYayv�>K^�e肶�/:�&xl�CtA�;����k��!��E���8�@H�r�*a��6�6a=�f��v`��hC�< !*g�����k��s�#�S���612z�8���x-���5y��J��T���F_!�;����xr��Ma��5��=f(��JJ�q0ڡW�ʽ����1�`ۧ��ʣ��_�YW�q���{��?�n{�`���̵i�{�&�p�84���6���e���4�9��0�A��kc��s�/�������� �E���Y�.��[Q#聅D��/��?�*��XBʆ�n$�݋U�A֤�F��R茡\��2X�9kGǞxN�&�t	f_8�r��g.�r�g,83,];^�q�\���N{��E.����
��}��rI�xV]�AcE��z(WJ�l<랈Xy�4E� �&Mx�7,V� ����5r�{���R�{�xZ)]M2`-;ux�ހ7�!�"#dq���e�����(�zl�+��6Q�	Ҩ�-t�<>9�VV������6J��,�����d���.�������G�#��<
�K���733�;�J���K���HK�!�e�
�X�m�n` �� 6�R�)�a)~��j2��,%˽X��h�K9�2G��X�@�
�uǌMP�=YǗ(X^.zڝ.�L��(�c�-WU�l8�7�,3H�a�F$� E~����w�N�w���]\�I�V����S�lh�BZFD�J�{6|�����֤6qK	쐼K;��[ߪ+���-Aư�W�m]|5i[N����0X����X���8�S-D��%�m0 ;�K�$��Iqs�EsT/��R����:!	sԦ�9q�wpz��B(�Oe`�����i��l�	-�j_��c<�P�X��l~iFp"��u�_��O�wO�FXD�	�4� �J�+,6��Glq_����@T��?�f���%��?���?����� ӿ���Hz��'K_&E.���fo,��X@W�btk4�`U��i͂���ވ\�6�3���)�Q��!�Dɂs�� �����H�LZx*T�W�&<�ǿ�����y��K-��
��8�S�L��˗mw�]�{��moS��[ES����y�B��i�knz��O��	�]�A��i�4=�<���|j?�H�ߥFvY����;���7ue,@P�FN�����x��Q�R�B�U����������{��z�B�|�^�|
�}
��W(��\����U�:;=���Ƹ�ăD����DF����ټuvaNS���"~
��w\�+�QP̳*�xSѭ��=���IѰ�����6#2�Gؾ?ؾ%l��'տ*�JS?�9����,��T��{|��z�4ė�g��-�0Ho��)#�$�;vN���w���M{����~vD��* )����C\=bjz�M;p�!�9DII�zz�G��s�y� wt1u��Fp��@���*'�n)�ʾ��v��u#}��Z��80h�$�~� �����L�����I���2��j�>ଆ�#!A?h�
�K�=^��{�xv9�K�<�Y�9@d�n�s�
(3�>w�0q�� ��Z��J�qϱ��`�)��5����g��}���~��6?�D�'�7Ti��{��Q*���_�,�u�S>q�%���(���/{݈)h�ל;''�.U�%h�{2%�W��ߛ�m#��..h۹
&��ٜ�������ͥ�8��m-�7
hc��������P�EH(��������~����{Z E��+�]^�+�Y\�,a�\�?0Ӗ��+`�zz֎��%RA*��K��A9��>��XB�rK���e=���6�?m�˴)�(�93�}��}?́_�����;;��^0�`�8/LhKp
s��3�yN������2xHeͿVpPa�� ҄��mu+��_	,����v���� ��oE�1��䳦FH��><���ޱx5+��=��A/v���ٓ�e��0��(�x�UYw9���;��\[n��m�dm�����)!���������n{�L�k�Q��L����ܽPb>�d9�Iwiߣ`���L��g��J��=����]�ۆK�2��"�VV��S�\heu�md*��,� F�2U㘌��=Y��ߥdvJV�ZA���F��e4�/'�n	�zjcH\;g����P?��!�V�2c�b[oчƕ	���}�,$�����w�f�U���WI{���¸�%+�X�i�KFF�%*ߖ�p�D��y�W�KA7��ӑe��.v����<��+Jy�dM:��2�U��d�y�F��e'#)����$@�LV	���^NLz��#;���NUǲ�XM.���y�gP���-����I�Sfl��d@%;��i�o�i�w����m�|��s^㙮�[��Uam��� ?�Jk{%���J�K|���σp:w��w��o3BBL<�)�/���	bX�|ފ�NA��<'	܁R B�sh���bb��u��ޖ�`O��`���Y��W������b����a�.�p]�'/��B�.>�{��ޕ� �GS��K�D�(�)�ͪbԆ/# �����Q�fƢdMR|o�wv�Y:��q�ж�-?�5�>)���0��t0��?��������u�l�{�L��JP;� ,��RL/�<<D����1��޽��/���K��7([ox��!�pg��(W�J�e���kK�+ٌ�~��K�1�����=��F'�j&�'m�;ۂgg��b:џ�o돭~����X��_z����t��XS럥`!<l��Q�U��/��4
���{�C��Z�4y���J����2V
�{�y���T������ڳ�_�7(�'�$q�.�Z)X**�g��'��6;��+^�/!�8�/�@X����h��s�c9»H'�4ԡ�C#ӡ�����9­�Y�7.̩�D]'�Q}�j�)`P0���;�ib���4C�2��4m��e�^�wI�w1E9��^�������s�r�+��y��S���l�n�6�@�V<�ޖ�:P��U&��
��t{�]��{����h�gQ�vw�S��E�Xm3�DT�\�vA~(W9�:3P*F*45��!�6�I�(�S(ɓ�^��9r�
���t�~.s��Uu�ǵ'K�f^��"#R�Ș�(��S�m}e�=z��6�������p*�B}vz�b�+{ः�^��q�Ί�� ��G{�)�Q����I����^z�EP9x�le
g�<����<O�^���܅F�W�޶7ov��0
���~��']4�1��:;u��b?����*Vo߼n/�?k/h�ׯ_g 9�f@��Ba��Y���G����}�A2Os}���gO��J�_4����'���{���C珑�
ߤ��tq���>BᤢV}����O?�Ӿ �_b`�M��V!+T�eL�+l��/y�3��)�w��1�}[�]+���}��#��5�n4�Y��R��硪s	.N�d�Fɺ����C��	������W������+A�����(8 ��z%K�O �W�P�.�c��N!��5��V��Fu ��8/I��Ց�bB�i��������r��F?��9��H��G1���%r5��h���{%-%��Ζr�y�t+�� y )���L�|(8�h5�e�*o����h=Ƹ&\�l���JW�� �D�[	&��%l☪�Q@�Qi����VX��ȳ_�E�R$$��	�@�K���Lx�c\��*ֺ2��K/�����L�±�����I���� OOx�k�Ap������j�B��x�+���¦� H�a(oa"B!s9���{�:��J����F$�!*� �@��pl��}�h���ʍ�c��6������u��?a���%�k!̵o�<�&3����Q�ܖ���<�����lͯ������pĜ��s^��}	�����]�K0$�I�n�%�8[�xp#q���*Y�bɠ���`�d�}�}�U�R8UX�>
��p�c���V��+kmk��7s��eR��.��o`Z0��#��	@i�x��C����\�_*XCm"3Ycm%kJ�:�����R�����W��V{�m������;��t��FG��JK8��ܥ�eMIÑQa�r��$N�| 4��x��;�;��.B�~���a��N���4Ʃ���KK�#Xˁ���M��7/�]_�n�K�h�r�ĤGN˻XcA;�����I���
*�#X�f����/��M���n7#~�>>���XWG+l]�j����V��OS��oY�I�a�+�� ��pL�(t���g���*�ǽ�G������_��O~�<�B\��Y`"/Oޫd���P����i��,�h���qg�����Y�ߚ�N˾��G�G���qV��k޳�ŢQ��N���Y��^ H������d���^����E�8�r(�ySO ��kƮ�,�'����'�ȲW`l�@Eڨ-W�\��oA��S'�^��}~J:b� �{�s�3)��Px�<��N��ha�౳�A��Q������ꎮ�Sy��w���0z��7�/���|��z��4)�CK���;������K�]��^h�wW�w�%�+9la%m8Ш�YGW�(#~�=�����(QBͲ�*Y*�����m��,i�']/��e���,t�9SHX������������(��+���}��>��(��('�Lz�m7A`+���I�J�	��3DQ�T�����ur|����n_}�}��7훯pxK�*8��[��#��kevv(
�����q�.~�_�i�P|���)
��x����n_}�5��������4n�B>:q�J�+���k�E�O��ϩ��(i�����`dx<¾��/e/q���\���ի���<���x�W�v���IlSZ/����0:��j���j���t�>�{/eL�����5}C�g)�*
�����T?��Ի|%��$�D���u֒Pf����`"=1j�0fmz���Uܞ�G�_i�7۽͵ܑ֮NT�������ʙ�~�����3jA�"�%���\P%�����,K\�Əp@!���|��6
���R�M>�L�P�26���{��|2�Qh��/�dmR���e:�L�x؝�nT�Lֲ�x�<�}g�s�Q�U�(~�Z'L��Y.�ZQ����H^Z�g3T�����3l��d�H����׿��<d��!l� �ߓ�
�I`c��:�C{�2e4���F��s�#����"�H�n$k'*$��&�����&O	b���J���^�O?�K�(~��e]�%����i�I�k�M�m���M��m.\n���(���H���W�ê�pF�x� Az��N!���F�R��\��Xh��s���5t:�{�T�=�F<��0��|��`�y����f`�~�.J�t�+A Im������"}�6L!����a|���á�2���x�F��ǿ�J�{���W&n}�w\q�7��{uF���g�,WB�0����P�/�к�C%����\o4	��j�`E{�����U@���Y��;�e1���v����F��5�wp93�����.E�2�ů�V=nDv��ik�#(�T�3Y�ӣmaf<k���I���y�~Q�R(��8�*��:Y\F�I��[O�A��Q(��[��0i�0�׺ڧU�\�9L�,%�d8�*��Gםs9�)I�f^,���S㔝6�� Q��ff=-k�-�hy��\�s[C��D [A�D�������c#����R�pP��[o���&�y�ʣt��j?Ʋ�.&�:8ܕ���E�9K���T�gΏ�>�oЕf�_+=Ɍ�
S��*�< �~w0Ke(���oT���K��㶿�H���?��2��D�R_��V���>��;(�ĘJ�Wg�e�{��8�d�"�<�Q�����P�lI�c}�\�6:1�;��c��༳ԎN�����.�rf�W�cE�J�Q贏�
�P`n����(�WW�խG�K]T��?�n������B��A�Ύ��L��F'��g}��PP��2}����s&���!<�3��Pd)��aM�.�;1���I3�<y:	�B���HN���x�������5�"�S`���s`v�TA�^C*E(X.�B����V3�(;�[���ǹ{i�:�$ʧ]�vN��/Xg�(߆�_�^�J�(�
p�����g�8.l�����\:�!lK�mc}����!����$
�a��˧���e���:���=�z���}�����<I����� mC��PH�Q��vp�P������}P.�����^���E��/�l���~��/��_?��J�^޷���^;DY��n�@����=�U�}���ѓ��/�j_|�e��7o(�K��g�	ʗ��1
Y�3r���t��]f�^��y�b�������K��[Ξ�e;�cKq6f<q�MX�~�E�M;;9ρ?�!�p00<���:ϴVZ��hWM�>�k���o{�+f������D���q�V�u��_e�����6(�/�Y���ț�c�+�"(�����uZ*-��~i��ijb<w����h�Q��Kɂ�����_��3XO_�=Yu����Y��dn\j��y9��+YE� ���UɊ�E8��a�l��iXv,���HD��h��*cu�'�؁�9�� /^__ɽ�k(Y�i��B�!C�T��ɲx���A0��l�*Yg����24��E�Vp��D�L����:�!V&��9M���'C���IP�[��]:�p��U����H)5�$h5�Q�g�W��L&]��t� !e42�H|��'��+�҉�&?9�$e��'P�����~�~�d	���C, N�����I�M�_a31:�f��@Z��:��f��h��FY��wy����d�+�w
"��Bw!|^���H�ȅǱ�Lp	�j	b?�/ˁ�6i�dW�‶����B w���=��X�Qo5��A\�m��ꄴ/u}�x~���
�6��3qK��1�yN�	��Vz���:?�R����=�7��������㧠ЇI���]B�`��]%~nx�������BhxT{JɊ��Tu&��Y�(/�騰��_O-\��ޕ�,T ��*V客%��2�o��#�}E��2G�FP�L�E�g�~�i���d�UT����p�<���i	�B�JmM|���u�=���YD��+_�i�ٵ���L��p��S�k
��=���8F�G.$�Y�ѣ���7���j�F�rfؚ��cqy�������dI鷩pU��W�X>�ŝ�E��0��p+��}�������&}޶�98
�#@�F,ķ�I���/�G\K��Ǔ�t���^���%`x���4���஗����G���ܙ̽����z���/�^>��7���Eh��8������ʞ>J���y�QR��ֻ�\��B\�M�(f�g���s}�0]�o��Ik>�w���i;9s&��9He�sU�~��Xo�ܥ}��8� ���	R�+��y��bv�OΔ�v�����,�=X����>�{�r	?|�*g�J�)YGw�ƽ�ac���٦AE�� n�G�2�(XIg*��� &@ٿ���d*�����3Y�p�x�����e��Ņ[&��ߙ��@�p�i\Gj���(�]ў�/�z���~�=x����f���u �_"wA����/�	�"����"Z�>�Ҩҁ�v���T���{\���Q�� �����5��n����E����Qx~ٞ���ؼF�����M{��5��׳���)��k�%��7�y��y��o�W_~Ӿ��I����훧/H�E{Fz/_Vz/뷿������˟����s�+`�l���n��E�:@�}�Ӟ�4�$�w�vPjH��/�n��嗙�zA�v	�O�����!޻��w|��a�F�x�"J�W_|վ������-��y���e;(a�ڝ]���P��<��RWk̢h9�vA{�z�����Q�N�2��<-��6�hI���VF�?j«t��ٷ]~�4nϟ�m�G|y{���>O���N�e|�{��X�	E/�wЯ�g�~|�!���p󀼙%��>��;P�>����t4�8�L�V��`y:��=#7�W��?�d9���/ߢd!��d�Lx��;b�L�S����NX�������y����SIʚ]���h0BB�J�#��ųF�¸�jjf:�;���	��,����z�����P�� {%K C�T�FǊIџA��[%k��Nuڎݤ����5�Wx�����,�"w\(k+�%to�h�j�J�}?}�J�g��+bd�� I�Ũ�4	c�"`��s��d�%�Ѩ��>[_K��vɃi�h�Q�6V'�� ����2���Hp �aiSG����KG��a\�ܓ&�!-TLcr����"6�̔6J����E*�H���T	��N��.ڻ���V�@<�\�5M��P�a�󄟥a��?��1��Uf�p��- &BV��7xw�4�r������#���;�
V<Ò+iu�B�q,�Oio�M��'9��N��������)9Tz��w�L�oɣ{O�}�:땷z�p(=���_�7!�SW��g�'qm�=���xa:fn��<T�k�%�!��Ib~�	'5�U#�9Ō�Cs��ZF��]Y�>����@�e3���~,�e�d]ed�bP���!��� �t0�5t-�A`�b�47����%���5��������^P0V*<��opBJ�)�P��$KC�S�'e���Z���Y�;ဍ�0e�i�oG��Q=�$t$�̘g)@�c��%��+[��E�d)X�_ns+9d&!����.�/M%E�B��M���?�W�6H�K�����7��M��;��� O��
V����q�J��lqB��O�,K��I����.];�>*�K�U��o�Y�k��{��ɋ���(P���Ϋ�������/�\}��_#�~�v߽lg'���	x�����D�̌+xf)4�8�+�rKӳD��+@��t.p T��G"YZ��aj&��.nfF`E��P|����Ke �=G�{��U;7�$)�E�A>��)\��8{ws�373���z�'�3r�/��o7q;9��d��Oʳ<���`�#Ɂ���%肃�*0��K��ߑ1q���c.�dͥ�*����,/�7��M8��������[I�!*Y��߾~�<��=G���^��O��A����r����=m����(�����G�ǖ�s�.�����C�(z=D)Y�i��0��v�Y�����<KǤw�~e��=�����>y��_k�s��y/����/�b��2�~'�R�;;��i.�S��y�}H;;{mo����ӗ(;ߴ/Pz���7훯��oPJ�y�,��K��i_�A�z՞�|}�R�����Ȕ-G�#�"+����9�����x�7�g�*9��Lԛ7oQ�������Ǧ+�+��`6����8:<F��m��I�q���0�2p��(&�}�CO�MTn��8s�����(Y(������(�o^y�ӛvB����v8� e@����4�$&8�D_����w���Q�����t�0�w����_G���(@���ʲ��/���8�}�߄Z&~͂���8tp��e�I��r�� s�ə|�u��c��6��6vq~�������J���G059�MS��2N+���!A3p����� "`(�Ȃ�
��U���y�A�S��Lq]�`#i$6"��:��"��<�]�����6�=��ե����Uv(ˍ�r�2��!����d�흃�*Y�'K��g����)�m�G'�q&�=������k�W����N~4����O�<Q�^�2��T=�>��PywÊ4a��_˻#\O��5��q���J/��n{w_?��̀�M%�Q�N�'/�S�F�(ɬo���H{�ɪd�z:�
����$8��f�<GQ�&FU�&r�P�@�ȑ��E�$=h	G���:���0W#��m����d���LG7=�}�٫�aɱ��#�uC��+ <�?A��hm���v�{�G=+ؖ����Ŋ"N���%T�H0[�L�?����/i�jɰKO�x�G�:ǫ�u�0�"�o����Q��e�Y�r��>����񑷾������)�(��M�T��2�̻�[2	�H�:���+q8�dX�S�+���S���*Yκ�h�cX� ;����MY�}�4`�g'9���ힴwp�ŝfO�Eܷ�(���0{�,�yf�����ei%kZ�,� �T١���hKgUd
>�L�j��PIg�[Yaj�Fya�/JX�M!R2R�̓O<3��5��uy���v�ݴDk�(�T|���wi���B[Zބ����Q𛚋�55���r�L�΁g�7f@A����go�χ��cL���/~o��GF��^�{��s�P&mK�;�n�Kp���Նso�~�B�+����p�]x��^;@�:�y�w߶ݷ���WO���b���7(Y_��/��,֛�O���N�0��%��w�A�U��}.�MZ�]�ec���,�q)`'p��BPhCx��]�����*T��3d�#���3��si�o^)3��
���u�N&���;:173�Kl?z|�=|x/�ЎO��
���2�����d:��vI%��<nb������{�b�mm�ϒ?k�"��{��I�+��|��Yf���4����i>{��y�|��|��H��3�NbU�<>,%�M�,W�\E��4F����l�_�xǪd98b���N��
%ke�=�?˥V�#���1�5
�{7�v��'��*<J�.��	q���o&�B��N���.m$z�&R�(Y�}�}rx���Y@�K��e��S��nD	w���|/��<�gg�\���N{��x�*���ۃ��C�}��ew����{�^{�A.+<:.e>WH/�keVz�lq�^:�c��#��q����&
V�c��1+���o��uP�v�� ��z����c^-�ɷ�k�qݳ̣���ӏ=h�܏����������7_���]���(XY6/s0N�,�M��]�ݽ�P�����G��-;[�,P���d�.>o���m~-S��)�vI�/%?Y8�9��O�LVR��V���m�Q�x�b�Q��0r��%'����K�����-hXFqK%kya�M��o�/��L����R�����)@�.��
�J��0n>�9�YT�T��)����5�W����p�(���.���U~�+ŋ#�ٷ%�]��(��U�-�|N��L��a���4��������O��﮿�v��|'������O*�G��Q�X�#����T�FF=I���vV贫mr;�1]�&�66��3I�	���.	u�IB���ע�zX�K�� T��q�.��CS�8=j�'��Ü�tqr�f���,�Ť0��K��%��bx�^<��6���57��.�rHZ�l��;;`�������àIo����"t�,��9�T;R
V�+��lbH�������%��[m'm��������ۛ�s*��f������K�2��$X��z�c����NA�l܊��l_��N��O��P��?��x��\o�d߅�c�����
�=���G #�݉>Ȼ^ʯ��b�Oi�4F�(y(�]����r��
AJ���T�h��7�ԓ�5_
��'iFX�7:�ER&�2;����h��P]��H�LF�-�e����b>ab�}�Ͳk���)XM��{\�����W�̽�EPHG�)��I�F
������ɪ���T�C�i�C6�RAA!�Fb's�Y.����"�S�F��~�J��4�i���3�V�l����F�[��~�@���?�!m��k�/�+9H�"�uO���^��yٞ?��}���3#��?��������/��������������=���[����W�������ӿmo�>������:6
������,L��[|K�:��L	���h�AA�{�N��`��I�
���{p<E����ٹ��F�k��Ġ���wf����^���M(g�/y$}�|�+;�$-��@?~����?h���O�?���Y��?�����~�6Q,��"��Ea���M8���3N��T�G���_/��ŭ���I������?�Fg��/����W_����"�S���!��U�䛺d��:��rd�r�L��W�� ��+.#�JW��(pૢ�+=0�%�s�ee������L:%XZ	�{��i⏂�
�S����.��Odt�v퀶{�Qt�E��J_v�Kf�?�<�{C�B��)a��'�y���h�*Q�֦��Йi��M����e�V�؃U����c��z��5��k��w(*���x�Lq��G*����{(\�<�}U^�NYk��h�p�V�ZD���mCF	RyRq>�q��<�7<��JY�8�@�>���Q�rB!�y(t��;�VƑ�v�*Yh��kmmm-8�~fWh<��+d���`o��.'����%9����$?sʊ������R�z�i���}�m3@�s�+��6��E?�d�tq��?��W��db-�������I�:�,� ǡcWgm�⤍ ӎ�!玡p���cīi#i]G�,i�*ʀO��k���]0<X��9�t���
�}���ď���ȧȣ�i��1b�T���.����D'��t#�7���+XvL�1�.�T/�=noSB�,f>���j�V�W�9FV 5~a|��߭�g�<�Q�Vr����txN�>%J�;��qa:����P00��d�}���q�ã3�9���=�X6@, k��,�r:gK�J��;��4�
��mm�w���T������~�e�(Rg�����^:�)� ��������zm/���qC�J���������^��?�	G痈�K�R�� W��Ns�=0������(�W(gg�P�`p�tnh
�;��ng��O�=p�� ��<ǫ�40}�%Lg��ޖ!d߿���w͠�C�	+`�h�_W�D�S�;��������WfP���{ʂ��-�>X���fV�OU#��a��C�~YĹ"��
Ƞ�]D�k�摸��D�p22i��J������˚���ΐ����}Y
8
몱< ��"4~
��	����q����x ��ϻ���2��'�� (YV�|6��MK�0_���Q+�����F�����������LV�5�U��
��Z.谌޺	3�RA��Zi9V��m3I9U��[��%��{4�h;BO]�@ұ>i�V�-��4����t�LB�����,Rk����5���A�w㧯I�l�r]yp
m��s�������V�m���~�l?��?o�����o�������/P���=��o��'_6�F;�{�?��G��c��ٓl��ρұ���s�Qx�B�|�YLy�Qi�~
��y��� .����uO�m��,��ҷn�r��۔E��Qz��jpF㌘�F�.m��a�
/㯭���>�����?i�����O�񟶟��O��}ֶ�6�_�S�R>���/u�WW?]/���/�V障�C�Y��/Q���B�_��g����h��~�?oO�=�^P�+;㱻�v;<���S0P\������pGڣD�u]�� i�W˯Q��mY��o��F��~�� ��a��p����4{�+�oϋ�݃'�wO��\�}Z^z�^���7�]x�iL�;���v�(�B���ʒQ���e��:��4�:�
˝�>=�����A箍I��QX@��gҬ�㥑��D�sвQ�aN��D�X%%����#���mkƏ��ܾņz(=�LI��������>����2y�t�S��ѓ6�����W��*�D������tF���ţ�'P(��4�.Q������ÆF2��i�(����H�����#�����������W��10�����+��۾(ZE��}4�qg�tІ=�����:��a�w�֝8�0�I����}���*~�y+�,�ֳ�ʯҒ���h��aVa�������6}�:mC��!g�Q4G�/�̖*���R�,�m����Ң�o��?{��ߞ�|�^��;k��������!H"H4=��8	` ���D�9lÊ�;
�)�xZ�G�*�d���ҧ3�D8O�q�AD�v(��A~1?7�6����Ѷ�����|��� @'���R&Ҵ������t��~��h{����^�k�O#]�Ը`�0U��#4�6ǐ[W-a�6i2��]���Z�W�͐� )�9p�D0��,7�Fд3`klH� #sB)����T�X>�eG%ގ�ĚY��q|���� *A�Ӎ:�]k�% v�!�	� C0R�(%U5G��0}sμG��bG�|R�⎽zO�]�Χ|;�����Gą ��7oX'���8��2@0F'Q'�)�X� /6?��,�i�c��j��]�����B�]�w��m�Y2�G���e�4�)/p�_%���+:PN��=6��-���v�2p/��:�6��36���!%y�`�ix�!�[�C@^��ܑ��tDIk?�����Ć4L���ԫ�����}'R�,-Ԓ�u"x_L�H!��1�K�D��D���G"a;�}�ߋk��>�����X���Y�c�.�.������F�f��#�c�kl�=Y��ֱƎ�jd�:�"Ky.�_t��'0㌌Cj������_E������#ܽ��=����,?{�t�B�1�RH��VuB����PV�q 5��1\G�{����T[�������v��r�D)R%=�#�p���L�z�>Agr��������z��0x.=󰗣��r([�\Bܥ�2n�6�x)]uͽCxH�3�E�TQS��(iO0s��r��?���u�ba~���fg�k	����r�]��MS�
�_�`�OD(�>�sz#^���� �6�^��������&���p��Kg�_u��>�M��M��>��lL{��'e�/�i;>|�@�e��r�!��j��Sů��#�p!گ_��"Ot��
�ff�R\Jӵ]hV�(���_gK�Ք��Z����
�E?����M�c��^�8y���G�3:�)|%��s���/���wH�����O%e!�+?(|��Ӄ'�D��n������1J��x����}����w3C3����,!�����ޟC��}I멢��8;v����%
����?F�����=/��kGأ�f�z����{�R>�!S����J���a�D�r?Ե���I�N�޵�Ͽ&���8�U�,�����F���*}v�vF�>>�錞0���VeJ�q�qy��p�=xp�--{"�r��Q������/�|��A/o�s��t-
�B�#�Q>�˔C9�?0'���3�F��1;r��Q�����r��\jK����ty�d$@�x���z�zx�%s���'x%�8Uh�K�Pn%�g�,��{�X��wPfP�܂�����3b
�p2x��8��r*���*�.��P��*����8X9I"A���s����6kE�6�  �y�U�0��v�����gdO3<��d=r|{k��./�C��/޾��_g��%�'G���3+@��B�*u��{4&y�ߔ�(���uU�cu�F�
C�K&�'~���?r�.�v��+�
��� ��]�}lZ��D� 
�6r��W���O߿V�G��bW�9�Q��]'�a�4����x�,ε{�#6W���b��h�2��Jֻ���z����`o�HT��Z�(M6��?�[���)_��[a^zeK�	W ���N'TI�U,�JD.�J�h|���Ph�e:�!b5Ⲷ��0��6q�f"��ᴖ	R�C�L:��� ��=��U,�p�9�ĪPڦ�<.���(1�ՙx��-<��}|ԕ�$%#a���|0~�R��$���>����>t-k�`i�._1�S�yэ�l�8T�>�g	Eg��~�d^̇64A�~`���gQ�-+L�9�Ar��Ԟ,���oa� \�ꦸ�;hk��S��z��| ��?t��U����e�G��?@���'$yܪG�:�������fy �P1�35�����p��S�`A~���&y�_}/\	���G���$��gT���	<�G?J�r�5)�Xij�|O6=�a̪\�5ܭIY�����#��}�1��zw� ��{TX�?�Տ���A��~;
pY����L��ޝ���S�ro��0�
���G�;J%]�Byn��Kk��i�E[,�����C�AhXZZl�[mee5����P�|����}�-�;�����T��#��(��Бt��U�p_����jEd��*|l������ ,�ON�ПiGdQ��W(��$o��Ս��P4���&Qh<��A�v�U��Ȩ.0O���]{�4�� GtNp\ԅ0�R�9��,2}zL�5-�&. p/P�������N�x��lLjy`����p���[�0�������o���������|�=���Ë���C�~����wP��hX�Ӿ�X�8^�����P�����?�h���p)"	��m�
����G`�s4�>�l'�ӇhmlO?,k��A�����H5ًO���v��~ �r`�=B?�~�u��z8|�䘚����u���s�8}��f{�h�ml/�o����"�{��kޏ3�����)�Q࠲s��Kɑ�'�IC�f=.����l����b����I��J�L�e�G�G�/��g��{��{*b�u|t����Q����m�����s�o��������87gI�Q��3�e�c�ey�%�`_�K�v@-�BIvoڃ�[�G�/�%2�(Y�^<o_|�u{���EY�m����]q�5mm(���hN�����I�'`���^�)�������:eX%g�]�܀�E{��y��c�_�@n8	��RJ��O<W8�-��Lf�����ٳ,�vF�%���h�wݿȋ(|	��!u�"m蚶�͙@|��߉+�Ê�=��ř�~%��Vt�\��zՌ�ư)�/q���|��6K=� ���Q���o^�h^ ��\��)����t��%��d��x���n���wJ�+t^���:t���?�?I���b��Z��96Q�8X]�TJ�T����]�s@����";Pn�Q(릙��C�q�nΞ���������:9�bQx���������~����c��O�ʻ g��{�$	�G��, �@�s铈"Q����i�d4�S�Q�x6#���S%+��{Y��;AI�\$�:���l��򎬵Ŷ0����oe�"�,% m@�����d��up辠�t�T��A]��e �4%����!�UC�(Y��w�@�J������������ ��<�1�?"h��2�2�VL\¥-�e���o��Ю�D�qYO�Q�ud�� �H����#XG�*���9�܈�(]�Y¢�Dx�_[3H�z"�p�wx�B��wY�V�*
֡
���+����'+ʳm�if�d]�:b��j\�s6�2�kz���?� ��U[�ޙq����=���c�����$�[K�o,B�<�D��3�����'y.k^1&��T��6�R��t���^��C=u��$���_��a�G���'?�U�.dOC���A��:���x�U2&j���>�M��x|���+䉳���d>���?Җ����%���~�2UK$��!�]"dLovf�-.������2[� �7�{\�w��v�r'� ��z��v���A^������6?7A�c�g�k$��0�.�-���w�侜5���v۾w�ݿ��ݻ��=|�	���ֽ���ݖU������J��_���u9I��@�rӿR\iRhe3��Fc��Ŕ�F	^Ja�%�~�1N�ʙ�����^���P��&�D��b�/�^���I�CSa����|���?�_k�E�� ��K�m�m{��
��vt�K�8py�m�O�K��hhg9'���ҭ �e�Pl���5�VEƙ 	�
�r����CY;�Y�K�7C�RVs���O{���.3C��Z5��W�,)��ܢ��*Y�'�ӽDipf��6W�A+(/¨i���.���-L�gfsz���J[]�O=Dn���ѝ�^wp����Q�¡̤ ����	_��9Ь�L���5��ϳL��q�^{�R����k�S�D*`�(P���~g��{y����T�q�v����U����|��6}p|b�-,����{�;��/�
��J�J��]R�L�Օ��b}��>tm>��T�%뫯�Β�s�D�v�q]E"ŗ�k�Miq�\ז�KD�O����d����\{���ѣ����J[Z��|zy1�⺗���)��	M��q���p�й~v�2���A"���G�r��S�v�S>si|q'�ŀ�Y��4����50���G�e���/^�͂�X}L�_6)��W���s)@ʹ�:�˳2�M��S?]���p�4Y���x�M{������s�q7[;�UH�`���� �2H���gJ�	m
C|��2�%<J�!n�w�/Sy<�3L��3=l�I�տ�3N��\m'���}FI3�g~��'<����r�mn[�CC�,��:!䄁����|��������Q��0;%˙��9]p��f��>��
 Y����3:lxZ�9rz,b�ĥ��"l�(5��@�".{Ґ�ϻ��	Ai1�� V���:J���
�mnv*3Y��žb:*[��k�$Cg�i��ɺ��,o�w�V��B��EҘ�*���v ,� �yDKJc�0�-"�TJ<$ZRK� l����s�5y�4{3��+�fL�_�&�:!�Ncq�R�	r�\AX$�Y� ��PF(��R�\
pQ~^�rF�,�Oe�r�R����QY�(&��/��X�I�3�O��3��ӳk�νWg(R0̓+��R�Q�h�c���3G(=�e�j4�	��#�{t/i]�h���;�%Q�ٖ�ԣ`%\��r�`���]U4�<u�~@�4�紋8����,J@��Ã�K�@������}*�y����g�>�v�j�v��q%\�wg����{�c*+l�c�~���!L����g�I�g�z2X}Uft�����2��	o�wy�#p��+@9ڔӷN���I�#��Bk���Rz��2���)c�n9��W!k�M�x̲3Y�n����PN ]vb���KuI���Ͳ?j���s����L����(:U]�T8	���i��u�6�\mn�o�(V�P���=l[��\��Q�K�ŕu�F[���I�cVX�~su1��'���p(����0�d�F�
*��� ���,�ZXt)�bf�T�z%k�r8�UW�t}JZ�s���mc�����|���?�_kP�k�R	rP�,z��Y���|}A?�����r�r*�j���٫�pO�´K�T�@؁K��ӫ�^Kϵ����4�����Q�F~"='y�z�萅��(�x��%� ��X�ڧE���7�pk9���(Y�$쀛�e]^9�k�@������QP��T7r�K�6�����0�������^{��%��[�K�j)�{�3�'���չ˶�d{Y�}�(Y�H`i�Ch�I��m/�N	t�^><)���٭���n�J
��xt��	�Ωd��p��B���rWf���*N��Km�����w�O?^ ��Q���q�Sx<aB��.�o�v������,�\D�Q���N���+�6��<qOz=y���s���t��ј�؆qh�H��LY�#���ڧ?h=�h���E�
-=���>y�~���l���i"S�f�h�l"|:��>I��I��0�z�3}���r��Nz�*�Q����X���I�ف�^ȷ]�
^�7k���fѼ�?�M�X�k�S�
����p˩ݔ+{�cӊ�Uʝ<I����x�F�}��]ZHoߵ�ƗgG_ 6�E���R��!�n�ۂV�zk����j�[c;�K�$��_iu�y��X��ESi&ݮN��`ߗ/yw6�iCy�4��T�7JA$��`�<�,�ʕ��Q�Q��G�9鳺�����/T��jOV7���BI|n���d�W#��tk��o�Q1$ ��i�4
qtk��G�|<"R�O��Ī���D������� ����Ņ�6;�"@��N���¨d�?��LV�d9�� b-T�$b���?��cT���.���6��,GWq���_�����`�K����j���ĭ��HBo�eL����7�|7	[g�D�~r�(���q����c0]5��At���2�!�S%,K�HC¬���l���12��.krM~��ʾ0�������*g�h7�c)X��:�=8�i^$�Г�!�wR�D�T]_���'�yf�$�./�dG� ��.�����Y���`�c���Tm�Q*O�I��oL��	S��$ʿ���P�^�LV�$V���~�#`�(m�wm
]����|��{�u;#������!ytf�o�7?�"Q��k�nT�g���!��ݗz��z�0BŸ{8]�1K�	/�J�#Ď�[Vg�=��E�}����^���#���D!̐x��Ɉ�.Oa,��Σ4�)؋�v�loo7�ΏU�H/3�(s�Jk��0�3Y�.�"{J��h[���R��i�?"MQC�D�3��U���Խv���(X��[mYe
�i&Ǡ/��)=�1����L�.���e���(^+�KK�N�����uי����)Zo:mV/�l�L?2��l�f6�05�ቈY*���Q�S��d�R>O.u�$�)�}��>U8���]Sa����|���?�_k��Є/����o���˃��=G�C�= a2�X^<WO�p��&
ܞ��B���K=5=]��n�k[(�+��z[ �\���������=ti&�C�[]�Mh��ۣ���AA��J�(��tz��/��4������R�.��ė/ ����]9Ga�Dt��e������fy����ʌJ�Q��7o_ei���̮af���Y�=�do
Bҥl�aw�J�+�)t[+�����f�O��`�U:����^�~�"�*3b.���]���,�K���!��13��8e)XX]�l�����_�Ӷ���p�ేmwo{XpL��.7(��So����L�I��^o�3��8�曷o2����d�_��Jd��� ����7?۳_���?e�Jr��fۣ��w?��=~�޶6�
����s���~���ŗ_��(�U�C:$����e����8H�aA�d9����S��g.iƺ��Rf���/iC����\(_(��ԓ8����F4�.�q���Zf[�e^����oB1�<�>�7��bU;%K�My��r`R�8=���
��W�P�Z�Q��n���+>t
����D=B'�:�q�cy��m߬~L��U�g�)�z.kHٻ��e"���0z��I�~ӯ���������ƙHfb��cd/�$�Ak�cz�)�^j~=���D鿷��6V��-Ҹ��R�z����� x��LJ�*Y|�I����e�B�VԺP۵�"��aX�O%��d^�E��,��B�x�07���P����|�
� �L;=�1���9ђV��c�u:�{�ԝwTdA�pyM]�v��!16���*`�9��/����Cb�!�D�\+j�z�9�__㙠I�6.�q���|�����B3KW G��li-�%Q�q�!U���B��2$�Q��t��D7�3��0�1���q��{el*�\*�r�1�yW�#���6�5O5�����x�,x��S �KuL�x���G�c������,�8��v�Q�l3N�Ǿ��z�6�?
m��7�֩������-�4��*l�϶
�� �tp�3&R^����|�������'m���Y��;��3�4NGXͫڴ�S��'����ߚV���J�m,_��s�K���^����@�/�Yc�o��*E-��A��ds;J��xrJz�	����
r��>�½�����1�Q�::#�'�]9��d���\?0Q�H�s�u��������Df��"4�}��yyI���/��.��M�*��o5|٦Q��m������>�:==��������r�vc{��!�N�L���mأ�Q� ���!6�.}v�>G3���|[[]�m��Y�IaS�y;k[�o���3��� b��GE�D�'Z�G��۶ɨ�#
�� �d�8�E�c(XC��o2�hxh��!�����m�aG�n��w��~���u��&�m;�G@3��F� �{��9�P�`��m�hi3&x����
����
 �
nn?l�}�<��=x�Yۼ��ݻ�|�X��������,k�l�J8�q*uѭ��8�*��^P��H�Gܯ�~q$�����O���t�=Y�L���3g.uD�.�D�~���>JEk�2����f��`�g"q�~ģ�U�^�~�N�T�;J��w�s&��w�!p@c
!�e��T���D��e,�{��A��U_X�)y�8˷\ʷ������;�TҔyh�([
�*[�WU.�tC������\۾�����?m�_���ㅶo޹�J

�V
->x����{�t��ۧ�1�mӋ�yv`L�Q>|��]`���i��{ld�B;f���K�93L��P���O/W9�'���J�����>F�Z#��6;-�0~�ճ�{��Y�S�!�^w�^e���2�\��{G��\8ئ�%~:��	�'�N�p���+e6-OXߐ�
?;���c�]~�pOٗ��֊%����n);F���e�V��C	|�P�W���C�LE���+�<�����cڣ��VE��߲���|�������g��.i�,?�#��ҩt�͋�J�䪚ݪ�Y4]^}����{���L��}���x}�P���E�P�F��G�S9r
%˺K7��G2ذ��6�c��r����56�v�S���1�>����0��ڬ��+�8�"���i�C��Z��� �t@*��V*��u�+����p� �@�ՠ]��+��O��ֵ���|��ԮKDW�[jq�~��bWļ�92� |ѯBr�5R����Yު_��g��=gƐ:�H�:��ȈDۑb�d8�|�<Th�}O�a7!O#�!ԍ͠��g��z���R��YiSskmz�Q��6��]�js��mv�^���j3s[|Ǎ�;���ʳvnްX���]�x��&�������vz9�OZ�=�n;(ƻ��a�C��|;C��^D���`���w.g�.�T�Br�e�۰8A Rx�J(=������B�o��]$��I+���wk��H�%�^��U�`�5�7�{��,IGB�bq�O�p)���7.��c�*	f��p���l����t!�-0�����㧟�W���|�Ť���z��@�S��ݸ5��C�RJ���0���^Q��{ �{�B��=f������<mO?�����rU�5�U)Y�y2O�<k�P=Fwsk;{��<��n��:	Յ���(Y#���1�.ɚ��$w��5�{�`�;�5��ٶ~�>��������?j�>����
�{�
4U� ��	�>Ҍ��K�I����4X��V����eY�uEHB8A8��.��c�I�fN��h����0��L�MC�:�9���T����Y����.o&��V˄��C�
�(��O��~�'����?�o���?i��'��������{�u��X�m=l��ڊ
vy�~[��n����ܾ�=p��'�o������j�@Q�n ���jH�5_��.����##P�*��Q�Ը��P,QR�3���LA�c�V`r��=��Ƹ|� @�e���$�BW�'�E��|PP&�i�N��YZ0n�UЂ��g�OA�K_r��r��������G���㌔Ku=|&�A�<��=WO�<i�^��저�x��eG��XS�.g\YYF8�h��k��#��	�����8r+�z�3�Cj���9�̣�3K&}�z�K����ia�s��x:�=qQ@mE�,������Х�J	y�
�.�vyy?�i�¡R��R0��(i8�G;K���+l�����g��`���9e��U2�2�tS�P����>����4�3��^=�I9,[�?�.�kT�\*��hc�ZEL\(<'*�[�J����K�%Ζ"\�v*xI�������ڦ��*�R%�g{<�/���6�v�=��;��������ִ	���>�@n�˭o�_�F�n��*�Efx�F^�y'� �����m`o����l-���(�ao����נ�tŸ%��KS-A�
�Z8�L�~��;f����80�Q@.e�N����Z"�%,񺆰\��@ά8"�2����m�t������6�t��YӵN�#B��ֹ����3I�6�a�a�V�%ԯ����ۗ���<e	������Nw-�
���r���/.����2gT��2.�X�WVњDQ�C���5�kd|��E�Zl�Kmrf�M͢t�x��n����6=�q��}��E�B��C�ªh��e�o���֮���E�#�X�d�Ӌ�\.|r6�NqU�T�.ޏ�Xi�Q�bG����}X������ՙ*�´L�b���s2^��V�(I<Ӊj����3�A�1n����+	
?�Jnu�����ט�Q��U�A ���}��o6�j�i�[8�on�߼�����V���GJ�1@���y��g[Q���op��|�v"	G�aN�f ��wgxL:�+���KBڂmO����$���!�3@�L�Ѻ��t,o��ٶ��k:i*\�0Q�Vf��j���W�G��wߙ��y^Z�/��g��#�t@��ʂ�O�RW�+ff(�$}vf�%�`ml�Ixg�gV�����;��q���i����(K���$/�T�ʀ��bf��'Է`���[��锑�=
�w�(����R����,xw����Hmz�¿�8;�e�(X�Khzڋ�<���TQKџ�/
hkk[���B����������)
֏ۃG��<=l������?��g�(���B��_n�Kkm���P��h}��ڧ���}�����gmk�q[]����(�Bf�_�|��BExTiP�)�P|ͧ>�=gX\j���� ���]�Ժ��VNE@���Rgg���A:LJ��/N�����{�+9֞B)�؇���.��>�i���z����bF̭���9W��4
�;uui�C4R;9<n�;{��˙��s��(LEg��}�� ���ն���V�����aK	� tK������*G��ϴ����A��Z��`�c�Ɠ�D��`&V v �CGt��i�r��9�,�r���a;<:Ȁ��I3GV����<:����T��J�r�d�,�䪄�/Pf����+�
�y��Qrp�˥;I��SJɷ�X�`��yu�"u�H��)t.uWѪYaqQ:_����2D�`!�K�U��'/*^�ۢ�5��}Q��L�<��8Kꅌ0� �;4?��ʩ�����S ���[�ϲ�1��VL�ڶ>�V�3D�+��%����G���g|�怈˖��Y]�րF��P���+ʞ<5U���A?���}�k|��&��c��ĭ�Y�.��g��+�U����+�^qfb���m Zn��J��\c�����[g,?i�~,&#0ߺ��v��C�DK�B
�^1���H��npwc����-D��1U��r�w�����;J��}�5=�L'��Q̌��Y#�������4�ɾ�#a��+$੃O�<���Ql�٢�'�HH\;0I�U�we�l�G�*!M���U
W�.�u]�kx�=XS!E�
�Dxs)��$J��
.LU;Q���ױ|ӝ�NM���>5U���ƖH{�η ܧa��
��ߐk��)�k�]
�bU����p,t��X�g�%JX�|@�� �Q:��g*Q���+Te��h�@(���F$�ó~�;�D<@+�4}���H4�H�2���=�K����nӿu?�7]�fx����_�A|���w��D+����M�����+o֡�K8 �G�f�*C��oU�rS#x
����:����.������Щ�eX,g�L�8���@�z5Y��)��@�ZL��pi�B���@�|���I{��1B�6B�J����r�٢�+��̜>
��,.�����k�Ƚ�I�����@@�a��69��ֶ�O>�N��{?@����om�h����>=�FG�;xG���KP�D�)�WX� tq>��B�@,�&�X�0��&p�_ᾏ�8�@_\(��Vұ�)
}�Bɡ�����f�������N��ࣶ�q��-�Tͯ�T-���9h9<c�k�!�jB>㳼dbj�M�̷���6�R6���V�dYჇ���}N���y�f�ye��l�h�V�e葸�~��	p�&�ǳ�X�6�^�i*Z-Z�	�Y�Ї��1�����[���{mED8e�!��efo<U0p5=��,@��?Ҕ	e��C�+�6����-���<J��B�CX\��3�px��BE�AU�P=��I��~��H~�����Sn.�ז�v/Z�n���ŔM8N #�����[?C'LUU��Q	��e��+ZT������Iϧ�QЄ�)�l*�Q�H7·������K�*9��rɝ��2cO��������T.�*����RH�q�s�l���=oz�S�X���&�2ρ�Rp#�-U�U�-u��+��%��%�**X�U<?��/�NZ�_\�>:���#�5p�;�`�k�~��U���2]�D1����YG��5@mG�o�,��Zi�L����`������5��4�K>i]���T�#�Y;՝�������TfU Z/����s�A\�(<��n`�H�WY�{���Z/��3�?�S'l��8!��I�s93JV.$�eEʠiX�D���-I��f�=��~��灏���DM;㷤QĮ�S�cQ�x�?e"����I$"�mCU�7S��h�2cG
��1+��y`�JI��X ˯�Ʋ�XK���<�XFC�L����5����_!���`�~$!��3O��;bV�7&~<K@|�M��"|���h�%z�g�+Z
X��΂:�H�]��0�:�B942A��qv�KǼ���ɢ���y$l١(O��`<���D�B�������t�:��߻�.�b��K)���!�g�6� ^��¶��8t8lx�@�N���:T���l_�oq=��{�6{p�҅����$=��,��r�[��j��$M����&(���>H����nl�M��:���ѩ�h��d��!��o�NUC�<R��>���*�'���ʔt�l�r`�M~�����Q��;_K+L%aT8�+�I[�f��!�Q3	�E�e
�W�`��Kz$m�
�p���A79wi����p��{���R��XG�|�>�����G#�=l���mr�}���W 0_�7	�|a�}+/�ӺY'i�ʐ�)���3�O�Q�xA����Ʌ?��}��wrז�#��@W����c5�jy�բA�#�]�j@*����kϧ-S&�R��C�����'1��v��L�:�wF�>!�p��%hu)��G������[��:����}����>n�Kk��D��x�\�a)i��Sy�RR/���E��<?�5��'�~rv	ek�~�1���([��{��ou�̀���A�f� h7 p������(�;���_xH)��#�02^Y�ME�t��J��-,�'�J�˺j��i�:����viT�㌍�F�%��s����977ۖW<%y=V�@eGE�7��=*rQ�p��,�5����A�p_�
��?�KY >(�a7W(EO�l(��,.-d�N#�����{�$�P��7�F�p@}0�������=��l+2V �0ox���
���l����⩶W5]|yʫ~��gf�j�����9��f���5�@t��!I����+.uF.�M�o�T
%�k�=���-x&-�>�l��_����, G<����"�-�A9VEL|Մ���jW��OTYY�� qR�۠�EY�,�H��ȏL,u�]�(�y����W�8��Q�q�_g��lL0�ct�/�QF��,�\�r�<I�vA<��9��\��/����������I���}o+}dqi1ʚ|�`H�����><[6뒲��W�Ѥ����cR���oeKy��_J�k��I<����5snBa��F�Qos��b�Y�����Dk��p U�1�vLzTC{�&��iP��-X�!���b���Hĸ#QS t�i����IFM�/>���<xE%ɹ'�OH[���rr	���s���ݜ�.qb�2z$�D��'�ySN	��x���c�z]3��*a$a�)�!ғ�xL��b�G8wٌ���o��a:b,�o�)�^3�F���JOR4��@��i�.<qqM���WD�|��V�x�@�(8�}��D�Bi�������=��eZ��u��a��w3I�Y\��\ ���~d�]�q�m�0���q��	�*lCѺ�!�L���G�\jmb��]&�"��)
�8J��K߷n
VEO5�%M�9;G<Uц؞S^�]��Y�$�2s�
Xd$���.!�?a�jvJ�`$��C��M�����%��l�!���u;; 2�:��=�i+/]�9�(�j� >m��3�}���W�#��5]�3ܭ��X�"��7Km;��5�!��d��#��	7�#�8��Hbt˔O<,%S{�����G�I�Qʪ�}�WJS���J�(�]FI�O��p�Ha6�"�X"���/� p�#��>�;92(���$����\b!�U����f)脞�}g��c�D�f_��0�G-�]�t�I\G����+h������
�,�nȖ���]��1�?N_>��Д#�%��l{��~�����}�����O���7��=�R��ҷ���I��>a���&#�2�Kq^00\��Z�G?h�RUK{
�;��̂���ѹնL>���>�Ώ���i���3����ơ%F2�径Kp�Z�M�8c�"���I�c�sT�:�M��&���J�|�_����5����`����ρ�ӈ0����{7��k�[G�Oѷ����{yt�.OQ ������ӯ&hS�V=����g?l�����r�ڐ'��o
�-�҇B+n���(�\�d<��=��t���z�����Ǣi����6����=��=�����'�kK��A/x�<;�pϫ> (�q�x� �4al<��߃�c�*iˈ������-J1�=�;>9�|��Ig��Yi���z�8?>n7�!�e�*5]�ݠ 9KC��kmu�}�����|�}�?l�G?i�'?m�~�i[�XoK(rk�Ѕ{m��6��3���=Fڵ'� G����3h���D�r��B��R��uO���]���C˨�(e� �c�]��#�/ ^ًI_���}+A���9�4�ڧ�rt>K.��ې�.����A�GhX�=��4���+�FN�:�U�3�Z��2��e<�i'�oIkBG:��Ix���u��#�gq���|ߺ"�hi�^�	�HQ��B|���!i(��4�Jm$��*�a���$���R�ZXj���{��UdiW�-��	����V��x݋��S�s9*������"	��CH ����ʳ'3�Jγ-�9tֱ�Wj����u�YZL����� b,���ax�@�J�KNQ^T���TB��"�iNx&��v9�)O(��X_�m'c(i�%��ن��3�C�2�b��|;{<���Kmkۻ������ͭ�����Y���iᄻ�K�﷏?����'?h?�����G�?�n{��;W���|�����ɣ�b|��@} `_�1v��z��r�(}\7'�c���T��ocȠ^j.�r��dC�Vi��a	v�k�W�O�Z���6B�?�˫�k�k��)�K��re�O��xԌ�3Y"K4l�n\z�I
��խ�I��"d����	�I]A���ru.���-�4�]��G��r��9��(�:kIM�M9�pR��s_f_�u�;{WN�2��I[6�;��無�k�۹2��W���&B�6�r�B���#�>�W��3��{��L�d�:]f��B�{��K�I
sh����X�X�&���m}��9���U�d
�fvʻ̴uK��)��ն�/����>w�3�o����t�wR�c�Kg1��N���'~WlS1�i�X������~�Я7�����q�~�/�}�>$
�χ�yvi�W�N�����%N�ߚۼn�f�� n!�~�-/I�����)���RQ.%�]��������^���1�c��G��%Ͻ[0Z?(�8�숴��0i�4����{��Oד6�T�k��w��Ç0��msk���/BgƉO�oT�K�>���&�)�-��ˁG�^����O	��~��������K�mck&x�-���A;3�p��4	�4�q�7K��!�e��Hp�� �%s3�}���׿W�[s����`�۬��^��}�٪��\��Q���}Y[G@z����~�W�[h�<����d�f?�	��M��
�����4|��J{��b��zb�b��_I�˙��L��E�A�X��ѹ����n+V�O��򚝴��T�.�=`�m	���K�(p6�!gP��$����w�z����?~��{���������m�������G�=}q;ta:�h�Ԍ305 �}9YbU�:-C�0�ʒ�j��1e�*:$����^
� �iy�OauD�^�yӞ=ٱ�n�,��B��Ni�4׺9��2"�e��⌶�
�]0�ty����;��~�au��図>(ig�Ǥy������hGi0X\��IW=e��Zr�#��V�	��|�AFi�t�	��+qk�CM���ڜ�Rѯ%�X\�8|F�B�ŕPd��Q'3:���K�TS�FHwR8 ��\��HZ"���APʤJd�����x'�|%K��1�mC>u~�-��$���ƕT��|��Ň+�2w;������n���`�x�I�,�|`�����ֺvss�ݿ���ۃ�Cl�ߋ�����ѣ�駟��~��������?�A�����>�������h9�᭡�/�з�a�Q��;E�F�E���9r�a�<��a�����ZiW�dIw�c����ѧK��x�lUػ1°�{�6^�t� �N�"ZIl��P`�y@c�E`�)t�8"��i�mL7�f���K�\z��:M�Η2Z>lF��4�֝�F�rV��s��[�X�Լ�A0�ʿ�z�B�sv�yF� J;���a�)I��m[�
�h��_x�vL�,��.S+{�h9åruk��b�ܧ��ޟ[�=e��В��0�4���y֒o�0ଫ�%�@]S�~�׵6eu?�u�(�#�*Z��9�q�`*^����q���u�NqǦ}:��x�U�|���ڴL��mR�m�t�_j9W��̝8���t��΍��2� �;��&��M��b���>�{~�1�*�����B����t�~�T޷e�t��f{�+WN��M�o�O���]�"vQx���Ǫ��pw����0�M��K�.lN:�c�p �ש'F���e<~���� �Q� a�2��c��-y�-I_I����D-��{�m��g�]�b��=�o��.F/�X�T4ץTu
���v�m!D{��_f	�F�u6���`���o*z�^W���<�e\ۅ���t�����myۉv�	çy��T�Tr<��y��
������{��| =yN�f���n���f;|����;�A�g,�=��r���3�K��/
��t��[j�ݝ[�@���i��'��)G٠p޴L��c	�r�z��=����M?��y�[�&`�-7H��>�w;z�Ӡ�_i���]aqq�}��G�G?r����?�Q���?���1B����ʲD�)g/"8�L�
����J��-t�^*��-3P��!��N�Rʹ��*j������|����/ri�G�{,��9xa�������|��F��?��lI���({��{h���4����@8v6+<P�<(��篮�I%+�_���el���r�:K�%���@�5��Ҷ�)����4�4�Y;gpU�C�T��<-�"��n��
gt� _��JĳlR�� 3(}�[�{�����G�o=��,����e��U�Omg��f��g��*��Y�b�(ȿ�O��I�Hk���Q��SDЯ�፸�r��gk��Mx'���:���}(����(���S�_�3.C3VW<8f-|�A��͍���ݏ\�C�z��G30����G�O�U�������C3���lR%����*bBܱ�zglqY�X_l�cCğ;m �kif)�E��ȳ��ｩ,Vʖ���؃Px�ူ��B�5{u�`iEx��b�+�i0=��n��lN}�,	��I!L"�M�H��J)�I��Y��!��Ͳ*\�/`�Se�Jܰ�%n����K]
>e����Y��S����Q�]�|�	��X߉չ��QUj>��{�\�&�� e�q��{����^����i�R�����Ehk����*X.Y���u	B��;�\B�٧�X�k3+F��@����	�^?�df�Fr��K]��~`��L�g�F�Kb>������g�e�� R�?0g�+�����?~ɛ���G�U�,���`�I<�͟np���L��Eۻ�T�K7Ow���S�B���wO��6�_M�3]����;��bsk�Y�
��I~�gO��X'�2��pT?=��z�Wi�n<�i���c�M�Y�nt�������>�׋>U����C@!��VyЎ���y���D�4kT��j��25�8\/U��G�;ף;C-��⎂�Ǧ�
��K�@�҂�J�����?!([m��|�2��O�ґᡱ\�� 댁��E�"/s �
#5`�x.w�)p�`�������*����,Z����E�|����Vi.�_��}�=z�Q��3��(J���2f-��IQ<����x�8�Y���τ��s�cP���ĳ��[f��3�s���C0ּ�����ɧ�Q�+
�q� �)X��ػ{��C����*P����\M���-S��p��wp�h�{�gD�������[47&����a�|yy�MM�	�(�I!�N���*Dk����*�J�}q�����sY���'���-��n�O�\	���߾����W�W�/��˿m�^��~'��%�Ԭ�H_.٭��r��
���8g�<@cB:!<�<?/e��~k�G̿w%�ʕJT)5�;����]d��	�gi�hW�*��Y`�j���*,�o�%����U*�Z�t��� �m�=���M��xa�S��LG�p+#g��#�U.����r������?������������m{s��P`��;	/2]�nʚʗ�K}�g*W����;-@���Q�����|�d�
�z���T��xc�ս�?ϑ��?�4��ا������x���-�}u����5��Y��Ԭ���j�.��B���(\��R�Ƴ�o�_���(c^x��&=(P����2h5�1�l�c�����>�c�W�W:Ƴ��B[����Z����%'h��>�&������&<h�dY��a�Vq��V��a���#B����&���ق�,*N�c���F�" �p	�k�ʼ;@P�[�����:Y~B��D,,�H���pu���:�1M��G�1����f�����!������Փ����+����w���{b�V�����~�o�v`vI'�U�j&�6R���^)+�QFWFX�|��(e�T�la/��#W���:�e�.#t�k;	g _�,#a�c}ע`�������X]M�-<#<|��-�5�;ﺱ��w�A�ō ��L��;�)n������� �v%�ӆ�5]�|�p	4x.�t+�_1��w�h��r�^x���k��Rr�M>&������_�mE��҄�x���iCo�����* ��h6�>��I���~�_͈Y��n~�+��p�O^��q�>::i�߼mo^�E 9�޶��q(�w�P�]�߯3��cQ�R��N,q7=vp"�w�o+Z{�����]X�̬�]�[��Q��FM�G%@�����L[Z�l��e�ݦм�X�ꆺ{ߕ6˓�h. ,��#�
-.YQ��L�>e9c�nK�%�e����7}�	o�ip�6J_�kd<������=x�>��Ǫ��7��(�,	���D�%3$��mւ����p�8����E��Zv(~�д�?��Pd��(��F[Zv��88MYƨ�dE�e�������uÇ�5}�5"_�0��d�`GG����0��~��a��a+�tE����d�tjff��"p.ʹ�Yp f�sSAs��@]\Bl�H�����~���,�k5�g���]SIU��RaObt	��L�,���� �6�=L_�����f�]�����o�������o?��ߴW�_eF�ڨ9��,�V9L�Ijiq��!8{i�G�;���)�CQ��H8]��JJ�5�W	н�[ʕʖ
�������{v�.N��B�	o.9T&3[A6���L�S��*/�a��>���6����9Ț*(�[p"�F�S4��W1,H���]2	<R���e�6����O�������(Y�]��?�	J��j�����~��}N�OPHX�@�ԕ��_
\͢:8hI��2h�V)e���.z������D�%�#�ۂ����CL���Й>Ϛ�1�m|�j�#(x���˸=B�-<���'=�Be��x$�J�kcC�j�����΄��ݻwo�"�g��S1�LNR4�h��S�X�K�u?�Û�n�Ao��w�ԇ���W�)Y�>�)�(X��u��.����_�HR�[S�;��]�`&�|��N���OONC�\�-��ְv�C���~eaE�>�ȣ�l�f�zA,�5"z�*�t����ܖ�L��VF������Pl�̨u����f��{��_n��Y7�u6�Zr����p���ގ�6U��q���/�	�ō��d������z�����)��w��Nr���{
�Z���:�����u��t~y����?�R��8g�<z=���0g+qI�-*~H<kA!�%��aӲ�^g�ӭՏ�I�2TK�t���3�e+
��5+p�\�޵�����}��&�r|������~�P���b��L���ꕤ��p�t����(1����ܝIYI3���A��� Z�W�.O�Vr`FҨ|�W*�Ў�F�k����6D3�d�bD��M��=ES�Y�[���Z�z�Pj��{�'�S��!��S��M[\�k��ˈ��駪�	Nd�ʃZď��O�km��:ʊ��6wM�C���[�����$�X	X2�k�c(ZK�mu�~[D���8c�0�ؑ�	G��ݪYjk�LV�gQq�#�&����iS��V���0�І�[ԯ�Sp@~f�~��9\XZl���٣��������=X(?
�If:N�X�iOåy�w��̅�߶��*G������)g�)Sּ�?ze%�aiEk�M�R	��e ��i�w�o��es
�"����R���@X=>i{{{mgg�e�����i��Ǟ��������)�7�+��2d��)�'y#�^!�S��L�J��w�B�'x�{�T������ laE���y��������ܶ��>�ޏۏ~�'�'��O?o�[��w��|������ߵ�%����?��{��eY��i�p��ZG����,��%�fM��g�^�L�����)��͛���õV�}?����+��X�M766�0̠�7_ݶ67�@x��
����O���"��~��K?|�֖���*��ˮr�fA�l���V�c��cx�篢p�f��܋4P���O��R��(`�Jܖw�U��((f�#Y�^�RiJ9��$\��6���<�ի(W��$#A3�ʃ��8v��-�rX�'#�tD�*P*X?�����G�������������O���j��(u�!�����	����Y[Qɖt��3nY\`,F��u	��gp�8F�-�Y�rVc����p��KY�b�KZ�Ų�� �igg�F�a^�����J�״{N��	����J���^۾����@w�x�{��������^̕��k~K�pwP8�#�U�!��S�ɛrNl͕�'b
��T=�N]��'��:/5'�9��h+k���J0��$��tąސ#|���X1�CcA�cÓ�Te�U�:� AU���?���/�v����a�]����,n���)�0�9~Ñ��#x�H��4No;� �Y}Iƺ({��WJ���M��P��f�~P�{v���vA��恅��+�6��'��	�g�P�&�)�&̜�W��{��v+\����S~l�NQ��f�ݛ����k��bU(Ƒ�������;���{�ȐK�*���ꄿ���!��7��_l�k�a@�oe����0jxC7��mY8��mp�˿�T'���տ��@K�0,f��0�����ř��_���CR�?4Ҹ������[��i���,�`��Y��.K\��?�Wy�~�����*i��
�̸�l9cW�/�K��o9,�t��p���N2Hy&"
���q�(n��g�T�g�aϊ0�,�u%���ɓ�MM�OI���?zx�}�����w����Hn���:�&�"��]xi
S!��8�Rv�Iww�fhk�Q����ߙ�̒K�^#��v��㶸�'<+	~�WT*-ǂ��6]�&]I� ����qن�����?�I��|'}�\a<���-�g@�fv�Y�{wۭ;w�<�Q�XzT��~N�@I���J���u��Y�ڳ�<�γ��,��Fqh���@�%�|�K?�1���2.ĸW��b]�ڦ�����aW��㒓�����4�~��U�+H����v'y��s�:��p���oY��G�7��M���b*��;\�:F��7Ȃ�G"���������oLH^��g���㼸fޛ�����k�P���g�|ޞ�?kw�?l�?������g���?����į߾n�~�M��o�epow��sVQxNȒ�Pvo�{p�^�w�N&��^;V|<��-�~Ēx��N����v��(cK;g�|���]������bf8�8��m��:�I�Z��-ziQ}h�Z�Ү�-�>����ͳㅓ��M������L*����U��'���=kO�>D�:��X��;�y©�KGʀƽ���.Ǭ��A�F�3�Ez%����M�g���e�xu,'c0��N���|���3q�gF�����ʄ���*��R�T�J����4�J���Zu���
ai/�ϕ��
��ظ���5��>�v���"�2kU��Ï����>D�T�,g�aj�z�A�E/ҍzN�%4�:2��+�ſ�i�'VxV��	21U ��� 3��B�� F�!5���g�Ux?�8n���m�j��hG�Y�(Y��hGm�߼3���2>�d��=�%<D�Oc>���ɇ6�E�)�JK��6����aN��J�Wf^ݞ���9e�9c�py�������Y�FAܸ����+ L E���:*�U-��S�rx�oN�`���2C�ʚ
O���T�a�tLڇ��zV����V'#�@���N�a*?��(qӖ
�]Ƚ:��v���s�l���|�=6�_���	$��r���_�%t����1�3��2�ŉ�z4o=����*U���a:��w(9��7����rϣ���?3w_���,��|����+p�q/���L����@$?j ��,�x�冔��d�g����fA�F�Q��O	=�u�t0��_2�\kw��l�<{ܾ��||���2߃.���>�fJpU�,�ǢV�T���_��7�\������*Lzӛ�ϻBp���|Ck��OU�Ey�v�*�3�#��p�W���D��K�	D W�*�j0�G����=o�-k�������e+�+Y*[�����杁M��$~�����k���o�J_EiE�����]�['�L(Q��ǭ��h��"׍��6J֭�w���ګ���\v� �4�G6�Zgt���Bj$�j0|pR�~~�<b߭s'?�������w{���MM���ecE�.�+��8W���J����'�� %k�`EL~b\>��x���R�q��D|�vN'B���g�}�~��_�Ͽ��ݻ���PW���{��'(\_|ў}�)J�=��zV>v�wQ�vs[�[�"�[n�.�eSu���N¤ �mx/��tow��Q����2�&ar�J� ��B]�ȓ|�j�
��a|{J���#o/��Є�x�V��(�^��呆��Rl����^���b��ब:!͒��n�(+n~2��<ݺ��� ~I�z���r�T��۠?��T�\�R�T�NUN�'�KR6r�A��	�ɘ}�bU+W�j���5&��c�L�b�3��1����[;K��t��3T��W B������&�9����1��Ī�	�0 ����Jښ�<�կi%+H�#����?�9)��$pA�U�-Y������F׶�]R�QI�9����LV�B�ᦡ�H C�v���s��8��kv�<7�@6�D5��p���,4�Zb��T�� ۇ��_�%`QRV��V
ئ5���Ì���\e*��Oj=�@�n-u� 3�`�$��@W����|L��� Ć!�� 4��vy#��pk�ľ���G�� �L������C�����%�<����|�Gei@c)Z�I^��̰�b={��fpd02��4A�c�~j-4��3i��+�,�4�h8ۥ��7`:��d��e���w0�����ٍ�p����5 ��6n7I߲tg�w�/�,�X^�E7��GLp�����;����ҫ�W��L�5�\a�{aG�^)#�iLg�%�{��b�v?��s1�1�V�M=?�3�r��G���*���5g��r���3�0Q��#ظ��m�*}
=���%]gKߌ K���;9��٧��p�N�b�򆪿�0���X%k�(ci����P��_l<&�Z�z��ϵ�X㷮�~u�����v#+W�����ݨp�`��.@!���wœv��˴/9[?��.|����y���bS���J�d�M�������!V��s�nf�gc� ���P`Hs��T~�r��,;JV�����I�(�+�_ƨ�n:�gBB�š�q�x���/Ws<���  ��IDATt��l��Aiz�V�*�o�Ӓ\����'E��5C�IH�O@���sʣ�ð,�|!��<-���,N��k�N(�w��Sס�dt^K*���`����R����G�������>�sI(*(��7J�Vp�/[��9
�]�����{�)�u*C���4]���$hvwv�>J��r~p���NV�wM�Z*U��*���;��fL�n1����~D�2Nx�[Z5'Oy�gb�/���! +���峾5�}���,Zu2V�,3�.܌I����*S�n����C�󂎛kk(���%���\��+�=��h��N���n�yYPff��v��_n��g�>���`����g��m��j��)(�*�����>U� 'TP� @c>ֵ}��>2ƪ�Q�X�C N����-���ʭ��&f�^�^=�Ŭ��π	\6����is�6u$�Q�E[?�g;1meU)��~��J�(ibF�?bDb
|�4��a�]Ă�P�i�0˨��3��B��E��K-Iτ��Ҫi��_Y g3�I�� �8�7��*L��J%��P�h;ރ�S�~L�Vn�Jx��������[�N�(%.].>%]�6�py	�>"������]pP�������l����>~�7@�k6�TW�b�b��8��7x�"�#�L@E�-��ˇ !@޿������ϼ�U0���+\}GÁEz�m�bd�r����P�-=����r��E��4�x_�YM�ÄV�]��t:�v�0���	H�8�G��\�awz�ψ؝/Č<t���*H=Nlʹ���(?�&�'=��lO��&ܓG��ʿч�7�{��T�=ωM��/�o����l5�Q�Y��:X��bԴN��.�*�0)C~ݘ�9ڟ�1v> T_wp-0}�o�ZZ�@��ik����\]���������G��W�V���Oc�$ 2r���o7����� S�ZmF}�<�� ocK�n���W6�f#~~3�����2� E�
y���H���u��?�f��������z����̨��U������oΗVVr)�[��B�so/¾ۏj{��BC��?0��Ǡ�wC��'M��θ�N�C���_�)�l#�F�Z�!?��[��#�&������jK�����O	�����1xC ���ا3�K�>_
����HY�Ȏģ¥Ʊ�t�R�c��Ii��F�dL�]W� @�Y����67i�3ș�[�g��Ӻ��4�G��"k���\e.<I�L3�,�dk�T�
��c/�k~������)����ʜr?�\^ޠ ��%�\fd���&�n^��&��Y/�ݭd+��
vq7�31�ʎ�� ��N��V"����M0���T�7�몓g���.�R�U�틤I��B�b��w�*�����%��ݻw'�:ܾ{;�����)Yǳx~kѳn��W�N�R�-�#Z� ��z�I�lC�K��d������ƪK+,?�6�в@��#�0����X���e��o�U[:%�ׄ��깶߂M��ʈ�;\\=�~NĚNd��=��d%�3�F:���mVQ���S�-�BhEq��KqJ^P�u��z5ސi3#���@U��^���0�A�
	NW/b	 l�=�f~vqbnmq�Z[]BXqv���y�f(��\�|{�#���������z6(�<����R{.��bW��]$9����8��s���p��Ն�r�g%dg�p��8��!8����vt|֎�;;����o������o��j�J�5�9{zH��EŁy�rs��Z`�͜n�v�}8�h�����F�8^G�pG��v��������N�✞�ig�����vqB� i��%] ���-
�:�g������D/�_���wg�t�	���7i � i�w;���m3'�)�W�����H�������URf���^�8�%]��f�<B9<�o3gm%q�q�b�6ic�g�T������A�vvخS����m�p�����a�����8�<����ͣP^s��V�\�AΪ��G�����qv�R�o�3ma��f��sܮ��q�;O��%�k��5h����E�]��S�������R�A��,	�a�>#���]B��������7�d�8�5�:�U�|��2�!J�,��S�M���!�b?#%�q�M����2:��)�gm��7���K���`Z��z�.�k��L[�W,/�\�|�AK>�p}!}��������kfs!�ٙ��f�]����2Re�^]8��LyH���|i�����9���.'q����k���Q�_�{(V�~�U{��(+w�(1}Bϗ|@@�[p9�N�&�0�d�n]I����H���ԣ��n�m��)��_�r���&���u��n�|��V�_��<@�0� ;���tU�-�s��x�,�fH���S+oMj< �荏���U�x[gB�3`�����Ԁ^����QS�?u,���<�-�ɇ �B�m%k��J�j�x���kیy�tx%	��;�a�r��w��t�=��-�>��G��V�J��|h��,�W�V�?�����7���fx����5�#,����@{��Nc�r���ɫ#�"�[��	�||v�N�5��4x:]��8J�Sx�홓����l�R�F ����k��v�sӝQ&B�'���ݶ��ٶ����<�>�<�-�.�����*�<�򇀇��S�N�#����݃���z��o�m�|��m����Q{��N��ԧ��v|>û�m��SW����m�~�$�o���~��,|��D9�����8�m[��	���k��L=�,��ԇ�v(�g�SV���.�;���~��%tH��6%�<�v�5?�΁BY�墽�Ņ��|z���gɓ��'������\��9h�{�iK�1�z;��3��"H�Ƨ������1�[3�{¶S�TFp��d�:��h�9v��0&-Ck���������v��KrlA���lyk�'�r���[m�zP1=w2��lk@��}sV���o��ݥ�֭��}�e؆֕�)2��9D,m�Ȭ��`��Ӗn��,���5r��<߱<J�uI��z���D=�P�ζ��kre��Td����w�*s�|���J��G�'�,�H�WYH�U��%I��xd��<�G\��pBȉ�����D�_�|$c�,r�g7�iw����6�*RN_��O���[J���n'e�/��w�8{���=�<���2�/�g8��M���'F~�	�P�J��������Z^�BPg>�$��Z�gè�Gk]ZL��#L�a�4Gyb깿I^��q*�?qT��,Vf��娙g�2���4��^.a�i*��l����O�g~��(�9��	x5)0���'�<�>C�9G�p�t�����N;��v�t
N��w*=�Z`�(��v��g��Mx��Ļzw� FDZq���3�p��,�}/��!�����dE.���}��aH'��
�r�����	��U���/�x?�e��=����3 glל��-���0V+�J	-L��mr,�&6�:����y��I�n�]a�ք�?
>m�4�?A��]ӻʵ�y7SΉ鈤	Kzѷ�?�I�2%�T�(r�s���ղϻU@�n����x]������a�+�<$��Kw���j2�F�♺£�M����0i�g���a�����v<�-��q޽u�J�i�H9�128�D��)�B�+S8��Gn/�� �h>�7E�#�����+�a��.���X�#��1�b�[c���ɛn�v������3��0�_���:��Bc�hs�"��"�"<9�9B����5�z5�'ɑU�����h}�H��[��ʏ��(��V�u�m;W,�g_O��ת���L�d�?�B_}S��;�q\睫}��L��o���O�#�{���
�u�d�,�1����w~~�����
�ֻ���P^|��"W��k"*�F�u�!����~��Hxp�b���^�y�~�w�����߶�o������/����ߴ��w�ŋ��M�l�Ɋ<u�`�*�Z���"�h�Y��Y���l~��ܕ�ms����9�վ���9m�T>�	h�	��}�I,��v�}/~���֒߄��M�m�1F�:���a��ۧN��N�����u��c�N�[���S�爛
MAx?
�%p��W�{�Ql��[7n�r?�{���!V�`��*������
4�2nP�\o7r<�Ye���<���a�2�<l)���5c�{���E�g�9�`}+3���U����i�gz�btO�J7�M���J��?��@{:���yd<���C�ů�T�aFL�z�NnX��U�ZA�����f�fb@�*٘Q�
;JX�/�M�`�_ppc�n���E7�=�R��4	0���ͺ��KK������2�o��2R-�i��qE�
�n|'�Jg]�8>�%v��S�ĭF)? �]=�e��:����DFB'�>�I��z=YH��^�ƀ{CM8ߓ8=F���u N�}��t�"r���b!��EA��Ob�v@:�p�[p�=���ӣM�]��>o����Te+�2��K{(bS~�Gݭ������o��C�v�}���v� �9x�	��;~�y�}���wqZp������ �^��2���^�<�M�K�q��@a�����{�aw��ፃ[��U���ϭ�*o��:�-r��,�QFv��$�Ц65�ۡLޤ'�6&Aď�c��K�#_�9�2����s9?2�O���1��U�0�#�'}*�ÍbL3Nk͊�bu������}Ӳ���C�V�!y�8Ka���̣7"93-�R`�M�*Z�y5(Z�Q�J�A��7Q��aӿ��&�6=,�'f��_I�桍w�CMҘ0���g�}^[g<Y6��Bwxn�Z�m���,�s/�PacRV�����j3h:�d;���}�(��mMf�?��~�س>�sо)(D8֨ D��8[�i�������^��#/i���2<#T�W��IF���8�o�� �0�z�q���c>��:���)�7&�+}'x�]�%�����W|!g~F�c+#��ho^>^��ׯ��c�a��QThZ�͸�pN^n�D&�>w���*�Ӭ:��m\]Z_�����_��_��]%�/�m���վ�����wߵ���v
?���юn����,���:��Y�Q��__x"U��{��n߹���y*��O=�Ÿ>f.P���vF�Ð�*���V�� W\�ۭ���*
*�����u�E�m�*U�;�8^�fƋО�_w2�������|�旗QFyW��#��<yâ��
�I��IG։7���G�;�u��<����A�~X�6&}[��Ҧ����@nƷ��ߧˌG֥�J ~��n�G�;�f�W
 Ҽ� 
&#�d2�ӑiF�0�A�3�{�G:�+(�"�I��V`~=�eL�x*VN���.�G��uQ�q�T������U2��Y�ζPyH��z3���N볩D+!7�*��i�siv���� YM�����T��l�f��%H�6�H���c
Y��3}�4i����4���4��Õw�����s��լ�d�
��e��􄸂s�����f���w�2u�"u�:("�(NJә
�
����W�*���dU
���P���Pbʯ�/	s�CWf��P[Ŧ��jek�c��1y>���@�OH��h��0oc��o��v���ΰ�֧��Nߴ��5� �xwv$���p���6?@��+�)���r~����&�	`_���M�{���/�c����F�;���wJ��D���[V���嶸(XCْ�;���t,B���d�Ğ9�1��5�:��dd^�z�~w�>?Ô��Ǧ�0�!�A���g�����L�GA����^wg����?����	Ye��T���PZc����GZ������L�����X�3o~d�׽r���@�J^���z��\C�ZBɢ�HDq�vGW��W�ˠ�@h�*���X��
��?�^)��Z_����Oܭ/ߧ�(g�o�U���wNj��=��v��|���߷����g6���1�+����޺���߀�2䂘�o�i!f�6�v�O�a��MѨ�]M�����\�ZXXwԔ��4��3άX.�w�Ne�~�ė��C'w��;w�׫���&��x��������w���O�{����N���V{��E{�����Ջ�����0���D���v��*�����<�V� l���S��㶿��R����µ���p��z��}�ݯ�wϿio�_�|��������I�C�U_^���P�����.�̠���@>�tE�����{�Px�
���{w�M?T���p3N�aW��E��AeJ�*�y�� ����^~����> |r�-����~Ol��`���dyK"mO�"�Q�M�t�c����s�l(���V�e�$kW���i��"�{�{v@X�Y�X��骼���O�Uł�W~(/�S��v
���e]m#bO��_'��W��;�Ɔ��X�O�+��k���w|�= c]�z��5���!�Y�,\V?Q�8�d�j��_m��g�d�#�id�q�>U�Nh+wӮ�O��I��cR��X�}t�7��L� 2��W�lfV��h+,��U[M#��mm�T��W��Z,33�Ǧ*�CԳ,<��"�mEv*+�FW�Q�����F�#�lc �`���a-S�Gi�I")
����ʤ�V��Z���zD&qM����N��A�Am� ��%�d]x=�[��־l��-}移�c���sJ���}��w�g�խv\�l]����Ļ<�}�*OW"��P �KP�:A���j��8��.e@a��)~'�J�	ʏ�(Q��H]�D��4����W(`(V�/�d�� ����#��{>>�Rf�
���8;|8M�;���u8?A�;~C=��KϮ�g�S�e;����p��Ͻ�{���m9�&�]���և����:���Z0�b���V+mBI�E���+h2P!���7է���0�*��m|�0DH����s��@E���s�p�q���Q��T�����'�U-��Q]=)%����I��H �����)W|E��g�T��%.�פJVȒ>��|��y��������0Y�w庠�f/0��{˫m��E�P�D0�:�t�1ևѵ����6!y����+<�K�@��ق�RG�W�H�y��j=uE��1�'��g"�8���
�4�fR�ғ�O? mlG�F�XA2���Q ��l�l�t���t����џ<��C�
��(|M�4~h�[��72�#|eA�=�r�L�K��Q�vU�ӯ2�]H�.ʣ
�A��`nߺ�Bo�\C�I�|4���P!���O���+��E	�|c�Yaw�m�}�޾|�6޼�6���ҟf�jFĝ�Pր]�3��N��2SϮ��d��a;9���gԔB���~c� pǌ8>k�G�m{�lg�4u�Oe �Y��FG=�Հ� {�R��eU�|�k�����V�T�Qd�C�Q [X^�w�T�n�h�����*��?�^PL���67x�<t~� J�j��>��o�<�<*UY�-��o�y��7-���K{�(�I���*Wچ��x�U�U:�.*� N,�9!g�;?�-�(qԭ�D$�z��7�.����fI;Q�}�W��샅J'��ȸ��
�9g��#��6�I�M��(�U��:A�t�jTQ�-w��h��~����
e*rs��A�B����F�
W����Lj�W�/T�o�:������'�
��(��	Nɧ�x��vU/�����1�}�-�g�����KEZ%��L?&^�_o+����¬�L��&�'�U�W�5UIU��0"��J�r�7k5q+Pa��BU�KT"6��k�~'~#\n/�c��*���r��3�������w>ޓO��U�"�Gݖ�%�#|�����W��@т��,օ篎a�����_3��V�u��V=�'��	v������9��ClW�	�9�Jw�@��ֶ��:Ômr(tn��]�T�P�P��P��\�>?.��-�n�l��i���Z5Si)��(4G�('�(9�(<����������T�@܄E�:?^�4	*P/�P�P�����d%��2
��6ʖ�M\H_씼���D�
�s��)�#^��ݼ?�|*d�n��mӞ�Ќ��\*Y3*Yϴr%�qc�~����͛
Z�e�Q����3�����V3��1C�I��1�q��<���w�$R6�@���<S758�?�7}ۉ����ɧ�)c�AƸ�;�.�whx38_��}�0�Ŕ�t~�H�K5��7W)���Ǹ���-�zо�k�A@e�³n]g�%�!�C�E�p-���������4i7�!�����X�U���W=�vM��c��D+��81�u@�1شA���-�?���:�j�j��N���-㭊	t=;c,M����7�C��+�>O���8[�g����5I�t�11������P:RȮ�}��s}0\�3�t��hO+�a?�W9��ǤJ�#M��b�*�Z�V�sŋ��T)Y�^'�/�)���+�+�q�w�=o�����w�>o������~�P'K�Ve6��G
��8�y�Z�0�r�����N]���s58�g���w�޵7份�ӎ�~y�96�T(W����~�A}GY]�A�w�j���ԟ�)�����2��v�������B���r���*l�ŕ5�ڛĹٖ��P���9���3t8w]�l9J���Sw�
��͉���/���{3���E�iW�|�PZ��*5J��R�dy�&�eM�b(�y	���.�G{xE��[��!?��D�W�5�ll���0��S�����S7g��L�g2_�ٱ�6�Z���O��r���=V{j�,���)-�P�K��z�w�z��3l�%r;v�_��YFy��Cv�a�qrj���72v�F��w��T������C���~L���g
��B�d@*Sc`��wU��j�tBx�42���!OD�����
���BiItR��8Zd��Fo����Q1���G�-�����4�h�N�n��$����j�ئbC�� �G�`�Г ;n���������� z�V+�t���g��8U�\Ͳ�B�Y�
a�X%|��aC!ę���*G*>(NB]�pu�B�Q���@�-]u��7�xU:��n9�S�FN��n�<w �~A��?���{FA��E��v?�]
ڕ¦��0nH�+@���
��)�p���	�\��>x�an2�>��|8}Kqޔ}�&��3�������{�ҕ���T%���a=_A���U�3�� a��(�c[b�VՊU)ZQ'+a��x�����ug}b�z�++Y�I��b�ݴ�5��Pg���B�� "@T�@����Lh���W�tz>WfʝN���Q��&�)I\�̢�$Wi�����d`y �I���He�/�r�o�w�#������<G~���+Ԓ���A�+��O�!�Yg��r�|>B�-s �w��Td�浰��*�<H�,??�G~��+4�����h��˔�8�b]X�v�����:˖��<�U�������v.�H�.���!F�m�c�*��IF��`��_�4�f���_˷ }Q�w�����ɹE�ڛ23a��j���.���#��ϧ�Z5qr��~7L����}���u�P\��wҘ4���.@F��.�@�e4Y��v̺G�DP��
�cAVe_89����f�VX�"�i��D���1=�X���B�َ���p�E�������5�0�\t��8'�*g���էs� ��.!��f��U�ʭ��<;�� ?[jK��m����B�{wo����j�([��{��i�Q%TUm�S�*�QvW��	W�t��q;C�����oa��J�x\V�\1#�	πW ��`ρ�|-G��}�'���U �-�PVl? �U��{؇(��n�'�p�a��_^I]���9i�s;6$���v�SW�T��M��q+���s����f���|K{!{��v'e*�[��n+e�Kd���'㊞���R���m�ʶ�o�3J�8yֿ+d�z	�n_��u`^�Y��h��x�Xm�U,iS�ֶ�P/8�0��0�t�	��1N@�
��1�"�GnF�T,�[񙬬Ev��9�SVF�ů�/�@�ΠSW���AV��]tl�5&��t";��{�3�=܁�(�AF�d+A�|��%��ۯ��Z��9�qv%k�i 52��t���ww��Pd��T� j+˥�,�)�P1Ư��*���E0"e��#5Vl�M7ۈ
�t����?�$� �0��."�?e ��~�u��QY��k��2b:ʎW�P��w�����8�U�K�w�l�	Բt�<�f�R'�2U�t���y@��D1�(=~P��04���������r�$[PqD���!�Qn��.��v���m�������}PA;�½���V6��0��*��?�sU9[���9*��u�7��Mάen�I��snMw�ܾs��Lﲭ����̳�H#� �]�U�z�ޝ1���0!V�4�r�ӿ����Zɂ.�a�T��j����a�����s Q�+�ŀJ7<"aG2%�t*ĄYiʮxq�K�EG�������飕o�f1�b��껤#���0�)�OIZ�-�������nQg m�L��IQ�@��!�o����k���ic�+H�G3x�O�j#�$�M��j7�s�N���8�;�>n��-�3���v�f1x�v�~�"�f�=ߏ��:�1e�G�}Sm�CStT�+̠-`�/��ޗT
��_x�Ԣ����:=�d��*(��{���.��13흠ڝ�ƖT��������Bӆ)���A��y�_�K�0��Q�)<�ϞE���DpJ}���Q.�@KI�~�r%?�E]8<:���M)����B�� -.�����K,� ̴c�<<>N�NE����e���붍µ+&�@xʚ
�
�+Bˤ�����䷲���$�Xo޼m�_�A��D�r�R��6DW���-�^����h+(�n�hk7V���\�����>\�:��6�Q&�ޡ��?r����P�AmQ�>@_*[*U^񎌎2��b}�m)+J���Ҳg����0���aß��#�poH�q�&8ތLi[��a���e-��K�C!`\l_����O?}־������||�>������>��O�~��~l�|T�&K�C�N�Lz��A����ӧOR���pe�ݹ{�ݻ�ݽ{�����&-A�����&i�V�)Gq��N�X���(���ca���1�z�>l_ʞ~���U�߈G*$�*S������t2Rp�{�+�WAe�>l����N��.�+bԗ�{��8#��Iz�G.q����^��+[�e<M���n���,�6ka��W�]X�����d��q�q2O�V�U�dHȑ�@��+d�D�8޸]d@Čp[�^���T����ސ@�'�QP7�ǥA?h׉f7%�dMWR���2��U������h���|ǊC#�y�	G�� � RJL���Lc�)gu�Ą�rE6�
Zۜu�.9�� ����VX��*�F ��7J�[ژo?�7����!8��#~�Qlù�&��Zqs%nfF�ū�t	���1̠�ͼ? �!�v�-�;����r��$���v�3l���F�vy������Z�X7
�E�so�����sp��L������{�v#-���0��)?�Q�\�7i��5>wg�Y�z��4h�����C�4;����^Oc�]�*\��O=�ob���7�z���)�v�H�	�sh;�k�#���è�%$X~��ɖbnu��DM˨�	�%�HC�j~%D���@Si�2���ۑ��ళ����߶�w�mwo�Ӽˊ=a����"n�q ��[�*����a�L߇����������qcY֑��U�\!pPBi�-��2�E҆�]��:П�3��&�{8L��߫}F{���&ѯ�𷽥7�\�IQ/|pf=��y����ل^{��g��/x=�7��`�0�(�ڕ/�_�A�Ͼ+��g��+!M����1�2�	4�����u��c��p8�/FY
��2�w�W����}s��q�heai�mq^
������o���	n�s�HE�sr�h9�8��Q��P�VVn�`�n7oz]������2x�Jv1�2����l]T��GY�>\ɷ���bLd��o/xP1P���@W�6�P��'���7�o�˗/ڻ͍L�ge�2��a����(��JZ},�>$�Y*�W�Jw���U.��>
�{ԫ���q�7Sx�\��g4�_ϛY6�#��&��i�Kz�ta�٦7���3��?���������/��?o��_������?k���W������?�3�O۟��������C9r�N��U���c�(��Q�~�G�h�����O����}��t�x}����/U�>��s���e�OI���2����<(�yK�ҝeJ�Γ/�Ըd��^�V��
j�~1�O�+<�H#�L*��j����$G�W�}�/��)P�T��������R���>m;v��_!��(Z�b���˕����$>٭��mFi��o��Ҽ~���C�;�����M%jT�v�~�go� 1�L��gz1&/!���v��T��>"B!�m��ԉo�02�qЭ�?=,�@Tq>������e��B��mS���N8��u��B��E>�s�w��.���|�.�I)7c��4JG�����#��Z�����S�j!���1��
��!V>pJ�9"�2Pi�bW�n����m��-��B�Im��S�r�J��9��f�1�+@�g�g���=�r�%�a+L����
\m�<��
�ͫl��� �T�FI����;�)�i�ô���!���Q�-�u�;����2��h#��ؖX��B����.S���64�#����)�wy��=��O%�/���T��+J�6Sa�j��C�|x���è���^��]g��+\��?~���
T	;N�$~����HǺ/�-��M��e����%4�&���[������LW�\N�O���c ���W�[��5n�>��L?���פ����2������I�Lꢔ�RH�-�������^���Q�~6É������o:���0��߇���j��ض��o��q�e�T m��|�`y�V?h�Ԁ�A�/������J�~������J�'3��C��B�����1Ɵ�		Gȕ~�u/|�ޥ<�燹'�u��#̒�B�+Yn	t�²��=g�D���"�j���:�M�
ԹL�4�¶������^���w�=G��(~J"@�l'�G(e�'�KT<��gp� e������}�!P%j���]�GO����<n�n�AH_���EW���`��7�i_������S�� ҏ�����UM�{�o���n�;���ݠ�Їx!lZW��+)����Wٖ(�t�D�Rh&�9P�Ǻ�&x�|�W.W��W�-�k�ܹb����2�n�*X�\ri؛]�P�R�·�������	�����6J�'�>m�'�D��������_�������������K��O���W���F�RY��OJ�?"ϕt/��\��ٶ���>��(f��_���/��?o���G(]���_�?�s������O�/���ӟ��}������G��K�Tjݞf9�1-CA)�
�~�XeF%DMze�,	A$-�~e*l���]�>R���x�c�V��7q(Hy݉	W���V(��@�}l�d�.�x����P��o�1�)��16@9G���8N�G��Ǻ	?*���+����|�C��q�i��(�╱�W�)�G��������������fc�mmYH��*� �6����b\J��U���2Pq^�k��� �d���y���S�8���[ƵbFA���N(r0+�ٛs:[:��
�8{��=WW��oB��ۓ�ڃ��J��@�l���B�];�h��[��m��m���ݽ,k�R��&5?+\�¶���as���:8������.ʽm�%g/��r�[�e@�
�#�Y��l�v��E�u�陹 O~�y�<*J���
l'�]��r�s�1�v-[�+�%Pp@雥����_;hIȸX�(4*�G|��e�eV��L����~��f`��qK��ZeqP��e>!������to2������ؒg�I�-۾�����|�.(�yg=���u��?��$t���y�jO�66^:囟��7������o�ڙ��C�ֲ� (o��jG�K��)�\VA��� �������ܼ�6Q��2V�H��3�8�L�EQ!�RX*Ӽ�bU|�\'��\�H}�M�_@N�E0���g��2����Ҁ�IG])Jܼ� ��V�Z��(��KQx�����q��J�Y��>�yL���pU����\}�rƠe��/����B[������|�[���ʫ׮dm1`8p\�S���mA�a�'�у��'��gO��Ϟ=C[��}� ~0��eJ��ؼ��=���&��Sg"�*���ʲ~�@?�oi�Oh�:�����Pe?�ͥ���ö��m�{Վ�w`c�r��3-�.[��zmAƃ�����5��O��)Ϡ9�����-��),Uc�z�I'�U�[�6?�i����nc�q�8�îv�F�㷚1�>Ȗ�)���=�]3"����ҏ>d����0}�[�fs	�B���}��v�~����{�|Pޕɍ�%��<Q ��6c�:�mۖ��(m���é�أ4�7}\39?����� Wul��Y�����2����v���+�ٶ�����6wQp�.橣;��%��+&Ҭ;O�5s��u(j����ZnwnηG�o k o<��Ak"��x�춭W�m�[���
�*
��ʻ���e�p�޾�m�_m���������y���­��x����㶍vp��A���axwr��߇9/�Xn3�m��^����{������]���vc�>9�Ґs�)mrL��?:���m�oI�zD1�_����.���tD�gʃs�p��~l��@�!_��%��b�k5�U�N�˷��o~�M{�қ��<��:q��nbó�]�x�xS��m/��Y�����xf߈�ğ�q�f.��Kp�'W�V���Ezsm}��}�z��Y�5'�#�HZ�lǃs�ZhI��X;s�nޞo?��S�(W�~���O>i���������n绉Һ�n����Ɖ�<ߺ��퓋K�����xA}�ƽ�Xp��]Һ�V�^2����v������|پ������������c,���QV�/�O���V;<�oeeJ>��u�2e�b��!���9��P��D�En�E�UιF�9ҙ��g����3����F�[+'�SZ6��R#hܺ����9+����E'nS��U|�*e_��J�zAX	���<'{�!L>�M�Gf�S;�[m{s��}�ʝ1L����+ɦ,��-�7HS<r��b(��d�3��'���2F�{\����Z[X����niu�0��?�o�m�h�e����VƩm�i�'ã#gaS����a�_4j���	8���I Pڧ(�[1�
F.Rq����= S5�0���z&I�K��~��X0~��B��0W��Z�Q�e]L��nI���) �U� ��	�b��aF:Bt(���3�#�yW������>���)?�a<K�jR�@ZCa��>�4k���i�RP�ś�-%�[�&�nW���3a��	�<���)0]�)p&���"B'"��PeP2Z����{��z.��*~�ɘF���uw���U�k����=0ލ� Bv��FL��ߏ�%(o{���/^�����ȥ�Ǟ����TB���I���iw/����EJ9���}f�U��K���`l�)��ضc�3��Ui��:3� ���*�}@�H�?3�������Jǁ�v<�i��[��&���w�A��;������B3ң|&��4�+i�p�G�Rt�=�u߀q8H8p�3'|9����DJR�����DP�/v#����B[g��_D�u2��s�ى0�ejf3��
��)&o��8��#���1��k~&���MOf�^�N�:��t�!L�#l�d?ȹ����~j5�(,-�h��nA��Z�0G9*S�L)�}�����*�Gf�'ܧy�t�+�c��!�8�C�j�׆Ogр����4�mR��V;�4A��Q>`�cۏi�2�n��A��"�z^�s4������bGxg؝�q�X!�sX^2��w�ۿ��n��/�}���U���o�w�_�/ߴ��^o��7m��6����|���k�Oځ����9*�:/�W��@Q����PL�,���i;pUl��nEoE�m{�݋����������*���Q���m��[�����'�}8	2O���"�v��>�����?S�����kmE��+^�P�P��������M�#���{��-�ax�<I���� 휶O���R=|t����z}y���o߮�w��~�$�;��_g�O3�;���1����VI����(;�'Ϟ�g�ﴇ����;�n��7��m�r������w��{w��ڭ(N��gIo.��X��N�����-/"�{������������s^�d��_~�~����?��_�?��?j_}�E{��~�J����W�PfvQ�q���������9�C;X��@������*L7��COLT_r��m]��߸:e����@�^��mllDYz��m�
�m7�m���l������ݬ|y��-��w�5Oth,�w �%T�q�$����� '@ؿ+{�աw�N�zw����# �w��s��@8Q�z�?f���� �'�i�l���0r��n��GD��	��y/J��as�ݎ�Y�������cA��&9�S���x=b�J��(�(�NBF���p��'�0�L�ſ*���`Yi�ExO�D�I�K@E𽃈����=�A��31�&�KeXO�S�?�U�m��u��f�K��a�5��`ԟ���b��6�+;f����u��Ý�_���j�Cg>W���IsV��r��LwI��R��V�j�3J�[���(X?j[�X��:��tuM%�!��դo�~�V}��g�k��\��gEV
� ?4���Fu�=}�r�k wB`����-�J�L^M�����E����	3qkWԬn��k勾0�e*�.�p��q�LVf��jғ��4y�s�x:��}�����d-/�0.1X*8��*�g�r&�$��HϾ�L�)I�;�o�C�qƔ�5���^�XRP�=�^A��ꇏ������aJ���2�}>��`?�O�Jn�:=�ʜ���۷kpG(W	sP���Y�m_#�H�zTQ�4��S|��0W��;��=�i���nc�#�i<~����L��ְ,�I�Lj�0 ���X�u��}n��bn�s��<B�7ҍ��(YЦ4i������$��i��f�������p������t�y��+=���D���q׌ʕ�X�x�Fa��G���1�#�0#��U���gZ�����VV]����n�Ȭ����{�lx���^���DxT�\�٬}�N/�p7��7�([��h�]G��A�<v��=������(��5�G%x�|�
��V�g�n��آX�8ѳ�v�}�c��;��M$��v~�BC}кmA���C;��w�mk���Y��<��2��DQ��wQ�Y�ԇ�����
��<�K(��o�jO=EAx�V\!�~h6���[��6���:sp����\C��N�ύ�C�}I����׮ʹG��_���<���ݹ{�--^o'�������W����F;C�ۛ)?ʕyT>�IW%�eԞ�/Q���Eʰ�3m�XG.��B;�[`h0� ��a)B��,��
��"��B��5/O���)��6����гW�z�ʝkk�������v_��ΝvE��<e��=�����{i�q̱J�����u�n��w�z_�W�y�7;���1o�e��(X']��w2.��o�0mnnve����P���ׯ�+���W(`o�-⸣D�-��\�I��W�#�aj\���h�K�*�*P7?(gG��A�&w+��W�͟w���ъ��cT#Fh����B:#�E������#s�@���}6^f8�����w�4@���a
���ԋ����#�2�\~�d�E���� ;`gt`(� [E˯���Q��,s	0@a_ϔ��c��d>��2)�̤�S0����Y*��]�)���7層�r��RPaI������?��Ca/;�'�.�Sǽ���&�S&yO��i�?ӝ�F�sfn�t[�J�NY�We�26;��,�R�{0�n2�c�r��'`<qx�0L�����Ai�>�7����c��b��+%��$�O�7黕�~�̻鄇��q���F�2�+S���J_�ys�w�i8��%y�%�B�0㆟�xNŧ>�@I�hs���_/���s�Z���;�I��IeA���������j�ժ���lx��v�:V �E u����Nf�,O�9�"��U�� /_���a��gﷀ=s:d�T�F��J�1��Ӽ�M���$���v�D�	�G�B��t�>]Q��vns�&n[�ʞ?
��4�#^(�a�6u2�`�?��>�pe>~��3U]U�����<P�dl��@)/P1�솂��%w�{m�oY!Q��ѿ"FNR���#2��d�)��Lݝw����1�Hxp����SZ�vG��a�L91��%�QɲO'4��u�U�~B9S[ҡDȟ4e����/����B�+T*;����v�����ɣ��矵O>�4�gn���	?t�G~�o�m�����w���������(h�qtr���0��\��u�ޢ�8/YF���n޾����<zFne��=~�	�7��#�
<�J��%|��������0�<��}J�O}Ҟ>|���}J:O<nw�PRh�k��muke�=�w�}��?yܾ|��}��q{��~{�J��Ay��

��ʄۦP(֖���;ڧO�Ek%��>R�l1^A������9�t�mq��K�*j(��D*Z���D�u�mr^���'�۟��/�O�J��v��-��"m}� ��m�}��Qn�n��b��*s(a�н�q*P���|��t�������
��|�*��3�e�m�g���~��4�����MO�*������*��)e��2�y��@V��/')w�
�|2���o�I����i�xp�q�핎�Ҷ��[�Y�2���C�z����1v��8f\��]��~/��C)��ގR��⾵��I��i���*^���^�BQ~�^�K��&�}�sB(e%��g�.�>�x^:E/z!ڍ�0|�aJN�7#���C3&d��c��l۬����������[�����O'w���bNFn�Y AW��:w)9�)a�����~Fu�W�r�ك�.��JM�k��
!,��Si�������
�V5d�dݻw�=}�=}��ݻs�)S$��V{�R<�����{��y��;A+�B���re�ؤ�,G�C��4keD kHAC�JX�ؽl��i�`�ӟX�
Vfu� �a�~3bZ�� ���|�Gi�2�6��[p�͂��[�^0(�h�Ξ�3���x>kʿ���1�Jh�Q+z�'�Fw>��_���pO����C���{o�L��P��.�7��.;��(��I�4�"�ǆ姎gF�ڵ��vma��-���O^����Γh�W٧��P9�]�[�#9i�-�n����\����,�02�2=>Ʒ���Z"#�����/+f8�[W��6��a�z�'� ���T�����R�y�x��C��M��1��3�E��.�!�;��"gk���\���9{-_��:���:���p��
�c��>Ͼx� vF��n]pzwg;���)�K�7�Ҳxө��Y���c
?I!��[�GH %̴�U��{՗�yQ6 7�M&fd����
+��v�0�GB2ގ���9���}�������mo���1��w�x������C�ٗ�����mye-8\�S�c�s\�0U�x��O���L9?rO�ދ�������S���BK�;L������6Kzy�M?�[�*�n���B�=b�u�[]���x!��uM�qD$x
.�s�Ϻ��#����|m ��G��B�R�%t�D<3� q���L�Kl��pm��-�3����a{��߶��ϯ�~\�aa�o��\����wo`�Q����ٳ�����(I���&,�=} ~�����s��w��ju��2r�v{��a���O�����Y��/~޾��+��G�e�e�'CW�}�y�J�Ͷ����+A��?D1{�r�4�x�O�!����e�'�x.���{�IOQB���>�"��3W~��g�������[w����\�n���O��~־���ӯ�l?��O�O���=A9�����޼�߿�[��<y����1��W�e�{��J���AۥNQT�PE\U�l��4���r�3D��/�P1U�C���U��������Ϟ�o����i�W������7Q�PJ�Jl�������߶�/^g������5x��E�@��eu��AY���m7o,�G�����n���s5����/�"����m�� *K����Ev]��L�z�������vQ���ܗ����FG	K'ɑa��||����M����(�c@Ҏ�e�1�@�BzK++y��\��ToW"B�M�9��>�yW[�<]�?S���1�&#��0�2����%x��um���8V��
��v�]���`��v����{h�L��ynd;u&J�a�u�]{<�U;^���?���U����9d˹��D��� �U:Ztbam�ݧ�ݡϫ�g+���o�߹��՛���uyI�2Vu a�J���u���G�B[�(YR���4x�4��X����u�'`��g9��P�(�[��1� �td�U[�1��4�}�Q��<���E?��@�VH��!��s�o��;m�g��(Z��A:;��2�P����d�rA,
�V�`.��;�����Dq�w�l@������`@���u�΃���˾�N���B}O�6� ��E�s�'�!�<�~��?J��n�(@��n��!�\��z��{�����M#�K���O椌w����}0�<���@�7���Vx�?mOs�~!��+U
���������VY�UȲ#d4�c��\_js�k��R��Wh�nPϼ8U}�� ���1_D��ܕ�~EP �=ϵ�!e�b���x�i�_O#�I��`�|ޙf��LM��<����ʿ��5�_��{`�K��lz�ecq�Z0O>�8�C�t��g�H��\JG��?d�n�7��	�J�L�_x#��/��}��d� n����Ǐ�OT����\����Vf�6Jw`�de���T'�F]�sb��<xD:��z�]�nʲ��X�O9GQh���
�2�gm���<��z�&㢛�p������	��f�ټC�:��f�v��z��>x<<�����w�?j�������C���*������5������nH����Ol�u:�����׌�q��p0|�$�'�po��l����mm~ȫ��	�(@U|�Ǧ�h?4;�E���M�44��q�Ş7�����1���,~�D�Ӌe��8n�>;�k�[��_�}�!������?���,�x��c��' eR���6izˏ�/�l�p/JĳO������q�#yE�r�
�]䒻�/-x��Q&Y��җ_~�~�󟶟��'��3쟷�>��=x�0J���7oނo�J׭�^&㙣�����������y{�	�JГ���G(K�	s���n.�����}��O��_|���b���?o��s��g�����ͻ�U�����G�����'?%�Os���(Z_�O��t�yܿ{�=��w)��ݔѨL	�33׳���w���`�Q�oS���iZ�M��h�:��۷SE�:J{�o�{Wx�>����?���g�E[r�l1�q��G����mB�{9��֮sƉ\��r���$�m{W���-��������P8;}O?9o��nG\o���;�y�"�w@��c�dU�pl�+D� �S��#�^����Wm��f�R��D ��c��8Q&N��s����_�_���Y��#���vtEG:$2e��n]�-�x;�y)����HƗ(T��BW��焩�?e���8���G���T~f>d�1�Y�~M��������e�l�U�::��5�n�c׎�~�;��Qw>k�?���e��(
K��3�FW���ek��ƿ
sŻ�-"�ܼ��nݦƌg�G~������u� H��?����/^�E�6���Cv*L�`�!e����de%�6�,E%�0X�-b޲b<`_kE�Y�,)���ڬc�"Z�I�N��&�YMAj	%����0�G��v�J�|)Y2^�&<x�*e��K5��
A%kgW%�T�����Q:�l;B{/Oc	@�h�|�$yذ Un�A���|�P ��E���[l�f�L�\~�PpP�0�%��9�-5�'�+����*3��
�b�;+.��s�#��z73�k;�qc�<��`<w���I�C�1���J�JW)K�	T���چ�Q-Ϧ!�>�$�4HK�{��J$��<J�Q���]��H�a;�O�3\	���D��@!
���g]^[�*o��o�dݠ���g����LZR�y�HZE?y�,Yn
����ٲ����u~���o�H�����/���ۼ��7��S;r7yN.�/H�i����I���(�(w�u�f��G�Q�E��//�'�2�������:��Y)"�����V[f+/�����𨉒e���8�DX���SDVu���OO3�;P9p�R幊���|����kr�����_ԟ3��<3rVtmM����]�N���mHQ�����R�V��^W��^ �)NC�*<v�&�{Y!�:Q�p�,�w�oڛW߶���vz̀���d �����c$�(���Ö�n�vA�Zf���q�"8I�R*����t���� &e�*{x���0)۔}��i�s��[�z���:���� ��[�5[�h���ڎ>rz��ʶ77��m��YV^Vo�eB ���ȴer�?)8Υ}�?m�	���g�݌�Ӧ�ƄX;]&� 6<`�~��V&�{�c�m��˶��M���O�ϻB��N�7w����A�>�7\�m',�s'>��3�V�Z@ɚ_���A}���e���mem��ɂ�gW ��
������xО�l=}R�~+�m�7nx��M���+�,�����Eq���ժ'�>�R�����Bu��]�C~�v5J������̪�E�=���*��o�k7�Õ��'Wo�[�+in��A\����)y�����E��}��(?�c^8!_��P��;I��w���x�D�c���o�u/�@�qUKL>����CU��� F$^k(���7Ic�>���
b�,��Ǐ�?����_��iƎ�?'r�ۻw�ȴ;(*��9#�2�¾�����=K&�;e*���qF�	}[ן�y�ow�ml�|����ߵ_�����՛�J����p�:�!�s�������mm��Q���o�E�ʥ��Q�� ή���?��6a=���w/����ū�m��@h5���` /��,�M]u��[u?���ny8ϳc֕�?y��ӳ��[�"k���_��1�;�zE���+A\��$���Q ��\H���n*KN`�ݵ\8��Sw��8�8�*�n�(Y*p�JVp1w�M�O�U9&�����Y�Ū��=L�g��z��H���I��e��]���~�����5���?���x��JV_�:�XɪUR�T�P���u4R0[�(X8N*�έ0(V䕒���KI�JRr+�LNc��p;��Y��m�6��t�=zp�}�ɓ��	��6v��Ԧ��Q�@ޕ,�,�;��I�p��T��f_�����H�4Z����j��1��Y�ʲy�܇|m 
�W�^[��UW���)��@���wuU��V���_E�+a���i/љQȮ-*f�����V	��PiS�+[h��A�}��
?�5�-%�tM[?�gP���=a(&��x 3�=��<W�I�a�Dv%����rD���2ZJ�ϓ���խ�p�:G�Җ��Ce�Ҭ�Q�=�U,��+��e%�&EX�5�O�p�)2ԃ��;�O%K�;2���Q�B�Ҳ�:�Z���Tz�ˊɻ0��ބM[?��O�}���8��G̴]�kD�����5[$TX�R��$�����3 \\��� ��:�W�#D�3<>$?�?88֖���^�R�,�9�1��<�zt%���W�@ȼs�a��(L��Ԟ]�#�{��i3M�s��D�r��s!`��,�8ބ?�*�̬.�tV�b�ܭp�)i��NU��3ֹl���EB��0��0�Ơ� {v��b����/����U��
7�	��L�>�z�-,�e��v�.E� �hd�(@Ѿ|���[�!`���ģ��c��1���� cK�~���m���C��+W)Yp���X''Y���zǸ�G;\F8�1��A~g*V�")u~�{�;����/���X/��+j.(�jAn�Ռ��+x�Q�����
��].P��:�ʫ��;�m}k��d��d��(Y�/)S��9��-��[W��޿���=~���v[ZqR��c��n�T��H�J��	*[
^�
�����B��PT��귶�Bs�.J�]^1��P��d;�|	�lAo�vr�ƫ��I��,�8y�Ǜ�T��XR��N�Ƕ��:~ ���J��{��=4W��Pv��z�UN��b�\�	%��
/�r�\yG�^zNݺz���Ro�E�r%���Y��N��N� hn<ݲ�čc�+H�y���l"�l���j?���՗��kC���~]l�w���9щ�|7�R�ֶ��T�\�������s
��u��������|���:��/��"�bdxA�W��G�J1Cڊ'(jo�m�_�������ߴ��ߴ���v����B����|^��L��N�!�����qM~i9�k{�y�	P�6y��=���'��Oऌ�B%O�g`�V��:�'�ʧơn73���w|,y�W��?�����k#=�f�q�t�����;����?c���t�m���Օ,u��D���8�O��)W�<@٤t����������ϛ�[��m�nq}��!}�v[v�1�����dmA�~�A�����P������xj�]��.��Y���s���DtiɯV;���K�<$��\����U,�v�D� CS��bU�V�2#�ɳǵ]�=��*hUv�,����Q�]�����i���(Yh�S�]�r&K�DIˆ#%����!Ȭ�^D��<�x�S����)�%@%+@����`��U��<2��SJ�D!n���k*.���)�/ʚ� �坊 ��-����F�IP���XU������L�����PY�V�J�*b�3�����s�x�/�k(]�nCiK�R�\��?�gW�h��Y�eu�v���>3s�����	({=l�w��;�v�-8��u�V�X�$��wCɊr-	��
�ȉ2Pk������ĖQE �a�����'�����({��c-�W��V偻^T��e<����z��b��z���_y�2V9�>a�;��Y����PJ��U���MS9�'������'՟���:�e�.dx@�����yؙ��vA�)F���V_��<��ay�3�n�O�����>
���f��ߍr�q	���g�GW����W ��Z�c��9��ʡ�^w��������iB
 d��Wb�M����
H�R��v6�X��Wc#\��woۛW���f�Ï�_�]��3|�]����;�=p#J�+��g�Pa�Z�}�h�� )���jĹJ>e~��C���A�4��)���C0$�m�{�$�8�E�L��ZŲ��o�ǥdI�ҵ]�Y�%@�w�6][��'b�ln�u� �S�X��ҧ?�T�	���v/�U�Ye�t�/P�0�J�=���z��n#�n�i��ȏ~���G��F�	
�NVT�d].@��f��N� ��+LI3�X�ƾ��?��ʚ㭇�)�,��ʺ�l�F^��E��u���$u�Ƭ�D�W���:>�G�K�QH��d�(	�3���W���o��j2��v��ȕ���#/>��Aǅ�3�R�E�ZM0w�P�z�V��S�����&��3o�Ca��
_]�E�ŝ:9D�z����7�՛��|WȪ�N"p�C��� O��lp�?�R�I0"Y��v�o�k�?��I���O)+e�8#n���_�m�Y�ڷ[�]1[�]@��@@���ye���n�SU�t\��2���o�}�~��sܯۛ7��&J���.��A���\�z�YޅE�s�O��p{C�ۍw�o�u��_�]�{���`�([ ]�z�R�y�^����׽b�2�I��s�J!p�@k�����h[�B��Ң�Ndx92���*�
ִ���I�>k+̳CM.t������jy��s��.�;��GY�n�����W��\�R�m���{ߝ�?�f� �a>Ҹ&�?4�aR���I٨O�Y�b��VL���5�:���3�,���U�G����Fɲ>Q����dm�4�r?��\�N�2	㩕�R�l��/�0"�Ҵ�!�j�
a֔6W�F`��У�e
7�x���y�c͒�=ѭ���
���5?D�����Zm�*YԆ](�P�͖y���N��d�\M�d����|<d>t��k�#=ύ\X	�~���j��uP�@W[�uTT������U�\JW��vU��a0�R�T����@¡��O���y���h]G!B��?ʎ��G�m����~Q�H+�Ӎ���j���g�6��(M��I��]���<�E��9�qC�R�
�Lz*q��ʕ�/�Z`>��-�v�ճJ����b��Q�I�?gp�О(yY9�})Y�Q��H%�4��9dU�Ѹ3�HAV<CJ�-�����&Qʐb�7#S��{m���
Lc�&z�qC��7�n*e_��q��*@���_����>�1����
���u�y	��u�P����.{ =[�0�Gw��3��%<_0H:8:�U&�O�Zq�:s�#���#
Q��}'�\[�A'��noF�P�s��Ύ���k��Г�F�=x��U��3p���DP���Ǻ��?(����[��gU��U?�����tO��������kے�����9��7;��no_���M�S��3t�/����*�y��9u��=?��u�f�=�!�Ƒ"�*��t�R�Λأ�e&�i��a�N9�4�? C*����{FbH�Wi����&Al?g��
��h?J���ΎC��#\̍x�nW�1�m��*J(�f[*���Sm�Sȿ<����F*WiR:P��O(o�Th���gG�peq�m��y�0�V��x>��+"^w���^�=B��\Dɠ,�(Y����c�s�H�y��]�rwI>�J�=�V�&tzN�Տ��My�F�������r��O#ȗ�����+Xzݵ��}6�H�͋"v�� �b���k{��UQ�b��=#�~��+1�🀗J�Q��f�7�D�� �Ə����k�Ĩ�mn�{���z����.�s|zDwF��W2�eK�t�%c�PB^�zӾ}�FYأ<*�*�Ɵ<��S�uHs�l��+�$ø��+�����}�飶pݝ	�dM���]p��|�Qʌ�fPTI�]+�<s(Y��Oo��,4���#1^������W(�oS&�Ky����``�pk��Ǐ�2�WX:٨R;��d������_�~��7��~;�=iGȢ�A>���mn���Q��'����� _cv����W��0�B�ʰ��v�h���F�F%Zo=̇��<z0�de"��l���Yc^�����&��%L���vW_���U}�����М��|�s�2�V�,�|�r����.��-�U��O���U,y�����Q�nٲ�xv��؀1�b�Ņ�m���\Ls"��;'b�<~�o�-!_�A�d����M)Y�[������W��H�d��3κ�R`9�G�A���ْCWo�C�i��&�ӽ�
DU)
��D>΀�C4�ʖ���v��:4��3O h�c=~�H��]BEf���w��o�>���������s�vv��<2��"`�8����,Yd��k#T!)!Ė��OVC��g�!j�Q�/eC&���KV�n�J�s~%���{&��Ul�{ۄ��-jmN�������@޿��;yy���Θ�ƞ�o���n��7 �B�`v�w�(Kkmf	�b�.�3��,�;ps
n�k|�7�̈03���FG�E�j�\����[4-�'�O�$m��&�,��rcڕ��$�5�s�w�:ω�O���k�ױ��p�nk��n ���v��R�^.�G��!����e[���t�5h�3gC8�إ�*����YY�=�Ϟ��*���F����G �Tf[0q�vr��Mg����0#.�x�Nƨ�d$��M����e��1f��J�JZ:���8��,�Z>PA�6/�})3�Q�\a�?~@�DM!��c%��0�L�!`8�;�Ʉ��R0�,�o	*���,��e�X��J�z��������J�'o��Fy��U[_G�p����D�H��0|��AD0庾��5`�-Ȩ�ۦ� R%
B^)�$���������!l����{(SR�n'���Rw�ڑo� �W�?k(����`�e{���m�շ��h�]�"��J�ߑi���~�������'��N��ѓ�+x3�6�������9ك���6B?mQw]�dᩡ����4�m�! R� �i@��o"D`��-WAƒ? �V�п>8�B{�XųmU7�x��ش�?���)���B�F;=�#�9��_^nK(X
bٚ��˚�rf�3����>N��+��9��B�Ez�8��V+�i�ǸܔAޖ�Ck���� ®T�W�N�h���qk���`�U�\޶߽�?����
�N�]o���R���J�I;<���\"8�~qyB&�G�=n��[aN^��
��e��X/��Y�e/��AQ�m�"Wx6�s��r�����޵�w�m!��Н;(
��d�C/7@Y��6��zw�io77����~C�U����ZIosk'���O%��:~ �o��]�w�6�C� 
?��R@x/8ϓ~���l��;��>���A3.]Ϟ��ݬ��?_G�XG!@i���@�>wpr�v��u��/��׿qE�u����a��0����@��
��h�S:�*�|�%S�����q�!�xW!pB`Ekqq�-�_�F�2E���Q�P�^��Ψ��}���Q�5/����mU��YŒ����Eִ?2+�qyj�*j�a��O���5EZs����v��/CNv�H���C�x�:g����zWў%?t2r�ՙc�c)��行�^X����bBQ�w��k����9�d�cPpc\d��ͮz!�<8����l��~���,�$�㊳f"/c5}O�6�{�R����q���c����3Z1ny�q���c�mz�����T�J��tU.3�j��W��P�vr�	'7�Y�����΋�v�<��f��G��*���Ud�*F����%�Yۥ��m��ö��uJ�N�z����\������������?���x������0G/� A��J*�ke	-Y�K�j��d�y�����W���"dnVn	7Pqm@g���CgP���4}��J���r�oS<R�z%��͕Z�"F��i�de%�����.�ș,��q��W8�!ϯCДpX�qZ�j*]Ҕ�Ky,[w�3t�Mf�?M���B���g��v��L�ρ�O��R��LB�����)�d>��N�r��$ݓU0��%W�&��2�TԲbUg��f��aeP��թ@���+�������B���9W��;q���=an/�v����J�n���t���L��?���#m��v��l�p�e؋.JYE���*\�b���L�+���E��Cک�A����/Ɉ��`j����鏭;�U�b����~R^��yb��$�h\t��ӻ��X���A�#|�2|�;wِ:HZ�QN���Tn̙$��ζ9�ጬ
�u�l$�<�m5�{w���/�/�ʖ+/rV��������+x����)��G off��p?+X�o_�-������=9o�Rs����mN
�U�𵶄ұ᭮���
���st�,Dq�3ᢴ&�T��:���;��N=i�np�*e�ܔ1{��P��3������y�x���l��ҺC�P�94_@��A�C�~3��?�v��|�}��ޏ�C�u|�UA�:�'� �)2���=�x�����i�C�Q�2��-�bFZ�#��T��_)&�	��Y���Ezo�sw��r�0n�S���+�56�qF^V�iz��ƶd(���r�1#r����ܓ'"҄^���7B�!���_P���ٞ�w�m[[o�j$}ғ	���{�o7�sW�ی�� �+@���J����n�c��IaA�}x�J�[��8y{���n�K
6�;�vmn5���Dz�w~��lo^��lng%����Pp�����a�۸5�ի�:�3�_�h�m߽xپ����g��6Q�6�vI׳<��߈���Ώ����u�~�����6�����a�� _qKz��m�a����r��U�ö�����M)M�<�^�̩�m�Ҷ{@:����V{��|����o����w�\^o���c��l�
�3����T&ry��������ww����5��϶7���Z=WAbXȢ�[=3���;�7��4-�U�%<D�F*}
�N�R�	9dRwY��2#��k��A�N�z����������oue�)���"i���7߶_��7��5���\�o���9���I��<"#�G�Yʐ�	�euø���rs�uO ��Ord�z|��T��I2)�#�dɣ�Y�����q���i��_qd����A�g��)[i8���	��Pz�q�E���H8һ���a�_��[\
Y�W���|�-x�Ne\�`q�V[�y7���];��奕v��<{�ܻ��T�Ϲ���� J�,g�  ��D�YP0SW� 4��D�:>�J��[�h��fb�DR�05+2�,�6N�O!�ސ���0�G�w��C�֏����d���G�[7��dU����Ra�dh:�K�*Ynt��I�,W�./<�^a�H�:�.�s�*%��Y� �F��F"��O|�UC�Hv���/E*
Yl �SP��,�~v�^Q�F���g��l��R����i�e�?�C��\y�:7U
Hm�n���W�G�EI��'�=��;�i��/~�p��l�ZV�K����ԕ�(@*B���=���X�4�����(wV���uW���j�X1$l޻RX+�^��_\��v����h���"�	1Lѐ\�~5 o��I���N��/ ���?㛾��?-��]v��	Ի��I�o�p�V\=��_�FO;&�埾���}ݭr*P(Z�.j��1}��g�?n�(!�:R�:=>�����~n����_�Qˣ,��R>U���5�,߹�`y�A�w�r�Vpt���7�ڛ7/���Ag��7���Ҙ<�ۼbf������V�\�R��eI� q,�P�)9x�J�H�5m|����(��i8m*m�H�[�'
QYo��:[���SW��(���#J���{��k�K%+[~���0����>���n�0v[z�qCH�x�/E��e&t��x�t��M��/�|\�j��/c�T�U��U�=�������|qr��\Y�h�;8ǴCK��=,m'=��ۏvN��vM�:f�|b�<�3�9&֛��I'�����;mk�97B�;�Ga�\����m�#1�%c�;h��Q�v��7�Q��ѩ}J%�˷ȡ�*e���c��Q�rU�I���:�0ٖ��,�����&J�����북b��0�T�^~���|�E��B!��?������( *P�P�޼�@���(m�Q��rC�[�X'��Lc?����D�AY�@Yr[�
��'�&�o�SAR�z��w��|�Q�T�^�(�����uD>�k��~���
��\Y{��m{��u��Q��Fy� ����[��o֣�y�C��8�d�҆�쀂q[�8`��61\�x�"i!Ag\PQp%�����.<�-{�!e�흓��*����/]�Py+K�Dِq�HЀ O+j�����Q�pү�8�ǕSx��P9u!7^�o~gq��o>���]y�;<L}���߶��yNl��3�l�>7�w�(��92}mʀ�UרD��ȿ-�23c�<[>1��*��J���(X��K�����C����i�P��$�TX���i]3N���j�m�(���};�Ue����ȳ�?l}�-�Bg"aF����mk!Cr�ʃ��o��;��|&Bz^���A}O�����tc%��-,n+Y}8�,��gn�Q�R�'Y���(Y�=�iH!H�]U�e*�Պ-(�12L+��)<���*�����g��[~�����z��n���nD��⪳Z�,��=�%�����}W�P��_�Sn;�yG!�7��L/��	�U�@y�njM�0��]��U,/�H �q�x��8D���˕m;�֍
�.g��ȭ�]�ʌ��x��f�}�vc��>@�|-ϕ�յ�ٳRu!�6��'�[���LCO��Z�i��G���sY�|���R�r��P�PtbO�����զ�(FY�T��^Z1\C���+���2�R��O�܂������UF��2�!q�QI�Y��
�I?��a�7	4�M;��?�1��a��y�)ZN��O����IB�bDƨe&a�I4�)����]��Ņ/�]�IEʫ������8��6b'b�}�P�d��ȋ.�l���\d�2�*�m��<��*>ޮ��!|��c���v%�A}��1/�Cpx����wv�Y.g��;j�B�Sc�>./O�s�I9�si~�-/��N������͈&�;� #@ܿ���;vB�W�Sy2�ȃRA�U�A�p�(O*X��P#Hm"8�~�u���Avۣ�¹Ӏ:�M��O�2d=��V` ��[�y;�k�8�A��w����R��n�8�Sޏ-���>c�?,�.�qyR�r�N3�����r\��)���3-�`
�{���B�^o��V\��r�4���F�Su��J����ڲz��wCvվ�����T�?���'�a~#�Ɨ����� ���n=���ڠ���)8��:� �ͽc���c���]�r�ۯ��I�x�N]%��b�u�؝�T��/�q5��bs�[�6�(�x�\�ۻ���N�z���
��<��R���<�}R/P�@���J�Gv��H�J�[O����8:��vCߏ-o��%g��r�M~N@�t�m�*Yo޺�����������u��w�;ȅ����F{I�^��
J�g�<Kt�-����״�������u6�E59m,�6�ŝ�& |f��㧘?�#W+��e�!��IHu��n�ZB��{d���-һ��8�S�w��:��d��4�W�U��I�}�(��8���t��UW�Y~Wx�/�F����b{�L��S�So�Dց�z>xkg�}���o���Љ�UJ��ig����Bc�*K��9���yZ��Qa���!��);cjL*Z�Y,ϵ�l�*��t��8#A9�յ�_z�����c�i3�&��'�7�S/�U�z�!^�ֿ�}]��������2TOs������8]>��*~c�L?#^_Zk�+7���E��Ih�������v�6��c}�,�w_�dmnA&���Z%�
$�:�UJ��z��/�K�-��(X}��ڲàlP�B�U ;���܏����.�+�B��3
�n{���(Y��i7V����EX	˴�Y�T���f�]pk���0#W�<�a^KQ\:X`��NӠIc����È�?�(k��!U�å��ݯHu,;?q�����a��'��2ʖ��������t)ZC��������V!+Н0Q�<G�2&���*a�3G��͸���"�
Ӂw��Oe̸?�n
�&���70W�J�ܓ�s��w�[��
S�b�xU��U����gy����hf�?�?Ӝ�X��G�z�63gi^۾wf�EklɪN_�`
�Sy����r����o_�3�q�h�D\�Lּ2\��
3m��,L�q|��s����/�1��/,�T�T��Έ��>��'x)���۲j%��֕+V޺T��lͪ�Cj�qeK��J�&¢��A\���>kO�<��<]�r����7��ߴׯQ��w)���<�C<P<~T2R'��30�]��)2�J��`Eɲ��)|͉��:K\i�r���/��bol�k�sE�rY�*p���:�	^��s��c������m�Ջ�����E����Ca����֣v�E�j�<��*U�L=x�E=ﰼ���W@Tĉm����jpӟg�:��&�*��4������X��_�j�Q����܅du��?��J�-!��g��In�{��wߡp��3�xٌ��؞���e��LN�U��ItC��c��r���� M܉\��T�~x«�� U�@O/�&�����e���(Y�{[�Ó��&�s^A��
ɻ�c����w֎��apnw�r�]s���?�nm���{��JH)]�(nA��"���(6[[<{V
%DEf��A�?�
XV��J�J�+Y�0�L�u�9��X��KI�Y�����[�U���ϣ�l�����ʊ��z���^7䩄�������Э�v]�>P�p�x{*�������@�z�������|��k���3)��j���)�
i��Q�N��~��U�D�����e�����Ƭ��� ���Yzv��u{�}�����>mO�>n�+(���%�(Y(���1��_�!��簆�O�%��P��RE�W�]�����br��L��'O�g��=�[(�Z[C������ZP�cyMS�+On�v�
^z�zq�3�������]U�萑A�F8�*W�(���s۰�0ӷf�rUJ��1aB��},�x�;M�+<�^t'n���M���+�<�������iX'�K��"auG�����L��<�T����q�����-GB�/<����W�<��7�:��
��H{������V1�֥O�A�.Ĥ��3�7����1�짔$�N"o�F���s����D�
�N��<
�c�&���<O�Hð��\�� �9��U���G�Z^	���g!�B�ts->�E9"�R�Tt�R7 �������0@+��M�^�35i��;0!�X�����!`�Q�TZT8����jh�<����p������37�ek��܍�u�ׯ��î�7ꂌ�3��T�����%!
x�Ґ�5�w��݀yb�����I���g�ke��8�I��n���v;�qf����pK���v����!�������J��-d7LB'�Zv"�����7��0�������]�/1�����_�I�2�/A�YJ�xO���9��:�&�ԫ�`ݎ��d���,�Q�4���[ �����&�+2����9��MH�O�-������:uNq�g;���6w�뗯�w�~�^|�M{�������Az���x�}@n��#U�7�Qk7�K�ן2ܖ���0�����o�"����a;=@��|�6N_?��u{��;�ݤK攡[����-����_���7E��A�"[(i{����.J��������}{(x3��2��������4?06���
�c�)4)��C>G(�
����＝y���V�*��6<��4���~|{��;��^�fs{L	i3�\%�.�9�I�X2�)�讦�_�����ġ)�b��h���~���%}�p�m�{�B�m���J���כH���^]�����l'��q�B��B�gZ2a 1+\�����sX���|)�ʍ�j��tt�A�2�7�y�+��]���NO��?��8��-�~�ju�F[Y^k^�Q7#����佀P��D:I��nپia��-��˫IG��ǅ�M+ϖy���BQ#�#_9�}i[���wʺh��7Z�::�&�0���:������y��=؏�*pz�Ջ���������V�<���PTpҼT�>.<���}�=�mbXe\@q~ia�={����g?�G��(��[�i̸��(�x8Qg��G�4�S�H/�P����&@Xi�=t~��Թ�����x�G.*�\�#�&}�
|떿\��8�jm�#��퐝�;2����X��})@�x����H�%�#>vMlYNね兦�7�0���/��L��:�O7�}J����|�����&��N#L��p@��L�@����/c?�v&�s��e6}�����F~�L�C�F��+Jd�t�hٸ�[;<����8\��+�u��"�Z'��W֨0뢐��*�w1y_�e�����F���&+�yx��˽@C��\FE����Ue'7��<�cDJ�z��Os�%��'��%���Cf	�T�
1��?�*(�����B����̂@���P�sV�b$$`<[
E'W�b���m�ݗ�W�r�n7i�o+��Mo=DS��)P7^���;�t@+�z�{��dpȅ Q�p; 9�x��g*̏������qs���9�6=W��z�⨂؟UU��JU)��w�歍����V��}r��U�)�
݇)e�,�z��^���tژNC�������rt�ܿˌp��v���6�˕n3�����G�i�c��݄!S�0�g�J&�#N�3)�ߔ�I�!#�` )>P�[�
1a�0t�Y� ���yx�JR���	�`�1�����|�po�+q҃g���k~h�K��f�������֡��a?�v=��U�~�d������w�����io_�l��hG{���a�☄~b,��}�������6�Wތ�5�A�?�]#޼���KZ�G�mo��ͷ(v�&�_�W�~�6߽h��9���s
���!$[W�պ�g���+e��H��~ciP�9><h�{;��`)�����@QPn���(��O;�o��W��Oh����Z���K}��i+GA%�-�^o������pw��p���f;����R��� ��W�����kg���4�
�gK�wչ@z�n�55ʈ���T�X�mށ��WKǏ|f���ԭ�o���h������~�O:�9�������qث���LA���	��Cв�x���Z��b��,���G^����!o�S��;?��vp���=��`��������g�!��T�9�P�#��TL�����(;�ܪK$�/ޥ[%�|�ϬB��s��Ga9����{���\�藧����Y�����?�H�I��=���S�\���'�f��ϲ�R|M��A,C)P��	��P{��|�='�?xDIųPԋ�?9e���I7֖��?k����Ǐ��E�"mu������v�9?9LzN��J[�	y���:/V������<�_�k�	
�*~��{'��GwN��¶�#���P��1o/���-�ŭ,��[7��7��H�7��(��\�� M����J�J���4(�*��^���1Ѯ�¥q�r'��uH�c|+9U���(g�q#���!�+f��+c�,���O���c��1t謄��)��z��g��֌?��Z�G�M�b:vI3���S����B�4��5�^i]<�K��C΁�Ӟ�����uK��#�$���W v��������&��ƻJC������%��@A�.�N��Yb1��S�Fc����R(<`&~8�r���$����0�g/�UV�6G+�g:N���Hj*Ib���t�3��3t��Х]CS������O�	�[;`́�B�P�0�+�d��ɿߍ0 �R����
a���ݞ��L��p�o��=�Ę@�;ǔ§����]a��+�ʢ���{�j�b)qW��*i��_ޭ�iĿ���(��F�Ӗ��|�FښzU�Mƴ>J��gl mL�z푖�E�~z�I>WL��¬�e��&�j��1^�5f\���55h�����9�!��_x�C���M*\*X�g��_��(�A*p��j߅:OT�U��7�*^���f��K�;�(:�?W��f̠9u��0lo���o��/���iϿ����׿B�Bp�|�����m4$F)2����s(`s*U��(X���q������O�N����V;|���{�M{�ͯ��oۋ�~�^����{���n���C���]��()�՞~^�������I#�M]�:q���b[E�RX�½ݝ�����2�ǔ����mmEt�0�SF>�y��W����1Ew0t>�qe�ϖ�?+�z�.�M`+����'�#���+	��������_}��m��~��ݜ��M��6�Z��6���z)J�Zl�v���Y�J�4k
�nA�o;[o�:��������a'�\�fQ���5��Ь�Ź��sC^��N��Htr���*,=#0C�WJ���jL�o6��턯�����6A	��	g����c�G��9޺
�G��Z�.Eu�D+��Px��m�7�|W
#�+����Y�.P	�2���B����iWN
*������!ЫЧ��s��z �((��u1K��R?�������;�#�����v���F�J*�RR���PO
�Ե��(+�r[���ԯxͣ]��2O��\Yl�?h_|��ݽ�
��MC�������v ��"{	?��fm����8~*_*pk++��ڍ��"�%+��~����[_��������%M�5O�,P���eQ�#	��e�2�ۭ����;�7��,˸A�Е<���2y�����`22�d5�um��c��1,�FΖ7K�%�U��iw��w�l[?�9�'�w|�xL������?2>w�J���}�����6�
����B�L�
Saÿ�M��K?��M�I4��7��yZv�Pm=�5b���	m��6W�h3�G�:��-4�D��ax;I���ׄ�x�Q�� Ai�K���E�^c��E���tCZ�ZYG�p$qՒ�(��ҹqWX���ѻ�,I�#3B$�@R4c��i���qJ!�Q���k�g����ui;��0���_��j�	2�%��jl��P�yC�W3�5�Ս1�b�e���W��|Z�HM�T�욎A*��� ĉ��0eO���t��}0߄�g�m<�5�p�0�����c*�~(m�\�^qS-ڄu����<ήe;`V�%R�r��J_
V�QM�����Գn��t�6�G�Ƅ�S�`�{�9_&�	h�Ug�0	3Ic����t?�Grw��J��=ekE�˓���Ϙ!�"�� �<�x&;Pe�(m��)n�x�'c�ʳD�}�Mf
�I�Z�v&��Wb�4�`	Y�c��/g1�M��]�i���޼~ٞ�������������|�^�h�����;�Y<��Е�
t+�)4��3���k�(j�o_�7�}ݾ��_����_����P��"�nm�A��ng(X����2��,Av�@��,����M��UI���V/D�rˠ(��,J����7��cUpO' �Jw�:���ȫSL��w���q�t�� �2��W�㪿�s���U��w��!߷�d��vs�ö�;����n�0o�{���0x�vwݦ�K"�*��*P(�W��*hJe*J���#l�����v���!���+�7�_���/P�_gU����uoF�r��LV�,P)Y^��K���aU�ꛣ~2�a"O@�$BH��
��o8����VVpP�Ԓ�JEMa����#����۷o�v�W�}��*B�2�b[]vbe�K~,�}���2�V�/�A���h��)����q�*J�+���6?һ����޹�ܿ�n� ��s��Z�)����e�-��k<����n�m��e���;z�/W�Pȩ�Ў���X]m�o�@P/�`���lGQ�w��+wȥd�"�Y�t ���r�Je�|Qb!�K��3(4��o�ݹ���F
�V�l+��ɑ+p;9k�6D�����(s��e�YQ)AZ��~�CI2Jd��'g��h��[]Zh���8��67q��$�tݺ��<O{/��n�ĝ�eU".,7�'O�1��'(|c��	 DBp���䣦��_���������򈐱:�=�?����m��X��.���y���te�|~e*o��Mj:�a�>��������?	\%8�%Y��i}����+G��Ȓ���p=�����ք�Pzm;�x�n�Q����i|���\�4A�&�7��WHu?��V��%-���H�����r�M��?t ��ƣ�I�B��)[������(b�UA"֛����f��5@����:����m�����r���TN��0(\e��?<�-&D�m���'P
�pO��3�1$r���,��v�C��C�d���5�ix�Gs�{;H�U��γ�I�'~�\�>��4��$���ɐbS}Y�EM�_	��v�2��y.��%�����?>g Զ@�>+ӱ��mc�)L,�;��3mc)ˮ��I��w�+���������y,>�^[StW�W8]%_>���PO݌��3�&�b��T���cd�V�h[�T��_)��W:��C�"���<C%�6N򅎅b�����y��Rm�]=�l|��5<ٺ����o9R��7�K��*Yĳ��x��r������}���/�m�w�����տ��گ��/�7����Ei���p����a�nG��8����My�b���oڷ���������-i������޾���&�������Jԇ+
���3| l�m�.e(
-��_Uo��L֗t��B�\�pz��&W�W(��9
���yt:�~��Y�� ~I<Ϙ^���[��z�`&t�{�t�����}T��)���
Q�N�2�v�]���uF�V?m{<C�����F���wvN�ہ"lmD�Z�"g	w�GW��V��Α��GI��Ӿ(�N'�n3�q ��e�,P�?=+k������YI�E�::��j�[�eiּTTǸ�n�S����	�G}��If_���a����r>7ϡh�Ť���*ߐWX񾓷8!�r��̣Ǐ�'�}Ҟ}��=y��=y�=��i��S�>�����0׎�ȶ7��DyBA@��V4��[7WQ������[����*�*�>�˂��mP�uk�=}�����/��y?����^C���y������<��Z�ϭ"��X]nwn�l�n���q!�>ޫ���UVT&n�ӧO�W_~ޞQ�U������!M�!u�MJ�N�V�ma�p�cxF:�6��QHTXB��S?�k-�.�)t����-ӆ���'����*U�i�ڦ�d�+�\#�q1D>�CZ%� H��t����U-(/arK�+q���Ey�<�xH~n�t��l^\��t�KK~}�2_Cw��2����1�)o8ƨX�`Yw��(w�)G�U��Pò[�p�D3�}�gӊ�60���Ҷ_Qt�5	���3���iL���m�#�~5W,+��)���g<�#3�:�S �r\��jb��i#��'L�<�˫!���y�u�.W���R��r�c��l:>�������~��՛�|����P��B)@6F�8�C!҉��Ƹ��f<k@�_!d@v|����n�aW�Pk;<����ܨ�L�`� ��|T�<<��#"�X��l�>~��ˬ����#�[PF�� ��r�71��斷�1�l�og^(AH���s5�=��@��L@f`Yk��a*r�?����,�럖$ZO=zk�6ސ}>v�t��vf�{�@��9�ξ�C��3� b`ۉ�� ��P[EE����t\@��Y�f���$P�
���۟��в�����<�J^��oA`�@[�ި�ː'.B��ZyƳ>z�T]QOV�6�*�F׼��?8��*�4��a��=� yAiZ���K¼G(��?��%8D�5{� .�A}�@��tF��
Z�6����j����g}Y�(��;N���椓4��X�Β�W)9Ph���Y#����؞��A0F�h}SW�X����$����>�$eK5�ee��b���C|����2')�����=B��1wٮ1h�!�\3�;� N�� ��Q���� ��<��ϒO9��@�:���PJ�ipX[[mk7V��{�͛7ڲxy=��ֻ�n�-|�]���� p�~��� FڮZ�:5 ���50�K9@[a�q��Ү3 ���������`o!XnF�{Fޢ�r���p���N\U��h;��^�U��mw�-J�˶� ���_�_�����o�w���(V�$���n{qB��7e��g�o ]�hZ��q��~i;���+��}2M�K�FD��v��6/wG0K��9
����K��| ��M=ԡ�m�/d�a�'}*�?����cS��z�����1�64m;�3���7�%z��^G�0Ǹ1��:tbm֭{3'����V��|}��� �lѝS��%mǴ��������u��c�[�<�s��p~�M�n�\Y���4X/ƀ�}�5ݎ�m�8�2F�͒׌�y9K#44�2x�{m{ە��-4����[϶A�D�i+�3�
ڎY�;}R��Gg��w���ˍ�v|�F�e��vz���T}k�Z]N�*�j��#/�;Y*Q*�k7����n��O��$�����,r�\�{o�=@!z��a�L��g����(Z��d}���9���_>k�}��4����o�P|Tzn�X�^i���l��i�~N��?#������O+��k�oyu�ݻ���;wWx7����q�߃�Y��O>o?��<��="<q���i���g_�����O�~�?|��߾O9����]Ҫk�>�K��Y�qE������ڟ��'��~�����,�S��pw��%l�Fnmsץ2�I/YEY���?���������~���ϵ���J����N�)�+ˬ.Ϣ��k?����W_<"g�9h�1�|�~�������D�<�]~������VV��5����|J�\�v��(�@��"���� �������n��lwn�ὗ����L;<n��˝���<o���E{�z:���,���P2� ��:^�q��"/;h��:=>;	��9z�P�v>Q:�G���bo�m����9�6�~l�n'ڮɃT8�DJ��Z9E9��@9E���M>;=HH�
�(��� c2OdL?�	Cc��ñ�6�O��Y�/_2�a|O��6j�#&��ؕ� �f@�4c� �:�C�7�Q�(��%˄M�&�������ʝ��v�^n�);4y�f{��Q{����NM����(Y0�u��Cg���l���H�h��,���z�3dC#���2>Ҵ�s��3B�G�00��Nf,ng)*n�\^��/.p��fJ���	�y2�,���2J�3A����K��\�q���溵}���ǈ��)�����9�u`)�3�\�-�pm�`�_�[Ϥ�!{�Qķ�?�|;��o�E�Ō�:I�Ǽz?m:>v���;F	H���CA��$0�;�Eۆ��H	�7&��Ch)S�����R����]%v���$������%V�p=�$��D�<-C�l�B�cz�I��R�-�nv�j����� � D<��R���	�Nˆ#V�t�I���������{��;*x�m�(��S���_�K(Y�t�������U��S�`�3���z7ꤼz��z:�tz��P���B�-cҮ1�+�+w����whF�!d�?�R�>�ٙCB�̾������ʔ�V}5�\ɪ+����5�2[ppݙH�V�`$V��m���2h�q�=@	���j[�(@�����@�]��,�o(Ȃ*n�ǻ��؋��P<X��5�ʩ
��W��zz��>���]j��=��6Q�T��!֍7(�Uy�޼z�޼|�P����}�3	*��0���ÞM+>+�/x9�3�U�����ĆV3a�pU>J[Y=������2�7s0�z����*�9��Ϝ�H��Rvi��!Y�I�n���#f��|�I���d��~d�,�=)S��NdWCuG��+G�8�QW��4hLe�å�b�m�}�67޶���\p`��D���6���S+pd�������;�줤�5
�[��(�ߩl����5�-�s�T�#§�W=+s�U�;��~��e{�z�6T�A�oz�-��
?X�O��JA��}`��݃�����~��f�?��Ys���1߉����?�"(<_�
���L��S��B�Wt�m_�����W_}՞={��q�=���vV��I>A�2�g�|EJ%�U��?�4��?��}����<Ϗ=D0����b�i��?��O����)
����uk-[�n�v���y}��v�=zp[��	���x�D}A���)��ۧ^1����'�|ھ ��>�O)��Ǐ�ي���Jգ���'�P!<��� o!��E1|��I�ɗ_�_����?�)
�ì�ȃ�����N��2����T��8�e�B���}?�*JF]���0���3�����~��Oڗ_<�F�1=hso���x�ٿ������`�xN��l*Z3�P�>@������/�����GWV�aʱ(�)�����7]yBA�?;��잷7ow�7(W�=���6��;��Ud(ަ��al˝sX�e�A<�����my쬝'+�A��Y������l��/���>��Og���3��4Mـ�CC�[
M��I$�a��*�Q���`>�?��X#�ob/�?�w�u��G��w����!��I�pI���b��L*X���(o�e��%�+dM�����r�-�T9�rB��/x��c����{wn3�S���������%J��7�4~)Y�F<��2V*Q�I�*L.�f�\���gK�y�𷠵G_�X����"D|���ט��<��f�l�qe�ٶ��`���$��d2O����r���qQ�;͓�,�ە9�n=>�@���6����Y>V��d���WJ���['����L>YXb;���-<�{�,_�/�������F�R�� ,G�� �t��(4�nD�g�(M_���%ֵ�Q���6�m��e�`=�W���-S��8U����od��`�ָyk�Zi��S���u���Ĵ) �/|_�&��G��T���h#����_/Q 8v�ʾ�Y(l*�*;��~y6~�����a�����Qu��7I�h̭k�nb��֏)Y�x������)��:��R&�I���Ԉ����L��|�vϧ�J��qL��UYlH�>�L|��:�,��>@\7o�Ҡ����On�"��S�]�ʭ?��̴u�Kٰ�^�����7���WP��ge�L���P?,��,����d�U��4W���} g�� '��˳�J�Y6����YuE���;�:����ì"l����}�{;9��!�=��]����y�>�*�;3�}V�S��19�9�͂���l&/(�e�]�Y�ԳJU�p˖ ܡ?h~�1@���sճu�ӎB51��;y��̓��_������/�L���_�<�����ʌhS�suȉ��\�M�Ϊx�R��u���߹�tw�����.�[9��L�їz�V��c���PGڣp�Y~o����L!O��N�F0���v~z�.:���#����la<����(W�6� �`}%k��[�<��>�.Z��x���'(D�=��K�r���|��0οz�׶v���3���}:u��<ܱ�>B��P�n�WVQ �D����$�����|�m|����
҃��ڃ{w�I�]�?L�J�}�ݒ�K��C�G�p���F(�u�f�C8����h=y�$ʔ����mmu�ݼ���̟��}�9�����O�O��b��t\�������Vp�{��<h�<Ȋ�-��;�����h8��j��$̭[�6��%�3��j�'�=CI{���w�o���w(��!�<@k���V��ܒ��Y���	�zx�L�Cg�� ��⣒}�����OPt��&j�m����_����۫���}��:'#mCH�F<�C�[�.�O�����<�GHi]�TV�6�����~�n�<s�A�:y�ۈҼ�Jnm�@����o^��������붾����|������0'��6A&�XUu<P�sBDy<��.?��>��Rj��/Zo��c����\9�I��×E��;�:vy�	CV�du���o��|�3�)���3�pLE�r��.qM��#�c��3y_aR&뎺��`�]P&w'��h�I}��R�n�v�kT%�I	�����"s[j���P�^�dm2hA��Gik�gl��dA6�GJV�A*�8*3d�p�~���(��(F=!�nY��Cf�F+Ć5�D�[�,3��l��r�"�ER�RpQV����T���ʔ�@�(Yﶏ����{ҕ,��%+�F�fOf:B��}к}��H>6j	`�ﳅú�y��h]-�8WDĭ��$��}��WI�>ejí�#!�M�Tgx6��d8���fT �ZP�N�L�m��uR���V��.������o��>I1��`r(iA�$�y��I�"֖6d,���*���R�^J\՝��8(���;Ä��.m����=��>r$�*g«dQ���i�P%�=mm;�B"�0���;��Rg����d�ˉ�h>�ی[eű�N�I��Wă���W���e��w�&_
���Mn��%�,��x���CN��-�QJN����_�@З�]�d���H����9P�~�tueƹ�-�ޞg1M�w܇��`�щ>/��^�28R��0d�����Ҟ�XByJ��O��?!>�i�O4߁�}*+E��s���CQ����+�Ͻ�^�dP�/���U֟ʢuXJP�8���a�<L͜{U�O_�䇡Qz.�����0'(}Oc����j�����+�t�5	a�Vޡ[L�3|�qä����_��/�����I�t��u�g�����M  %K^l�Jsn�����ν�q��mof���(�����M��^�^�C�\e�vbT}�����&+ˊ%�\Mjx�J�
JJ�с�u��?���ͳW�oo�m[�������������*�����(]no��L++^|�� � ����Ѿ�OR�������7��K����SW�T��܅Cx���'���o�-,���u��};������|������O�/����'���ɧ��c��;��Eouy~19�K-��\���FM{��ʪM̵�e��ʵ��{y��=�-�x�?��qeg�s��a>��{Pwnߌ��%��#���(sQ|P�T�n� �F�_�����8�I�H9����[dZ��	��^�`�rs(n�Vٻ���������v%Э�˫R�������mnmJ��R!�o��`�mP�5��v['�l���ZIE�gu���u/���*���g�X�|ʝ痳�u��͛����z{�v���N�S��O�xVIZ7���\;A������%n�9��A	q�SK�@������2�0�dy�JjǏ7���P��}վ��e{����V�=]~I���
�*�]\��m��fy��s\��� �M>�y; װ,59W���G�ǭ��*Ya�v�p�}��/�1M�J�w��	��qbm(Y"����G�yc�X�a�4c"g�󴷦��;�ǎ���0�p�D1��/�e�J�;��j<S��0��wr�>�B�T�ZZ���&���Z����?W�h=����J�:���ma�WJ����:��3Xc��Y�:�e8�W%�!�O��iӃH�0O��x�ʀ�d���O!A�'�s�`�� ��+Yj�����-9WJy[}�K�I�zt�>�\�R��ݻR�ꃽ5�d99��*T�����Үx a:��?�#d�8����0�3�X���=�ԯ^�]��A���t��)g��'�^�.�UB�5f's����J�/
��{�Qq��PW���?p��%��u����j^�]���@%2��$p�
?�*xvH=��c��i��UQR������Nޏ��Tg@��+�n���vw�,���'����.���/^��Tl3�JCa:�O�# ������{i:�*/?6?�5�&��g�Q=���`�c�_����8cSV葇��fm���H)X���;��A/?�/uBU�Ϸi2��7iN2��6�S����D�PW{I�>�6��Un!�<P��we�F�LS����m{{�t�C���7ᗴa�f^���/�W�(Y�k�+��J�UB����0�r�־|�kj%�"�k�O�?��Y�u��ɸ�!S��1���VQ���3s�c�Mю�Q8�̤i��<X�
<�m5��ڶ&q�������Tcm����I7~��A	Vi M�Q�_���^��z3y�_��\�q��}`m]�r俯G;�����gQ�h�I2%�8�?�H�ms�UW@�;��h#g��d��lC�E_SХ�2�i�Uo��ue~Ӿҩ�G^�֣|��	T���<���w�d^���-���9\o[�޴�܄��m�`m���h���Ǹ}D���nŉT�_��Ms.D{�w���+�*��yr1�6w�������K���Ej����8���@3\,��A#�4,�,�x�Fr1t�9�N��J�u&�����3��tcf�`�?#?�����=$z�^{�C�����z�]^:ձ�i�iZ(�SS��PWqʨ8iO���k���^ad}�~������rI��(��Η�*�] ߃vL���l��w��iD��,�^���e�r��g�e�E�+����q�M.w2����Z֧)P���:�6q=XY�a�O����xj4E�B̓�j�a���є���g��8?���@JN
���Ӷ���޾{���Y��ݸo�W��������(�܀���`ǒ�1
xw���gSa�Ζ�tP���͓���F�����#�ӰI> "��p��0�Ω�lُ�$m�,�rԔ��������5�/�]�.5���.�������wԶ6������{�h?�0�FV�Q:�";�3�b�j��:Rv�v��eh���wA�����˽>�N�%���Ҙo�Y��ozҬu.�� B��a��6��QtJ|�p0��kJ���� @򿯜��^��0�ݹ�[�v�u��2[�����5|�+�A���|��*�����g������4٦����2�?�1���l�V_XZ�oc�T#� }�E����7r
�������UL��M�_�$5���ځ�^��`�ܘ�� APqZ�*��8�� �H��B�}G��{���� ��B��0C!�J߹��?���\��8Q�Ew��ɿz�'��;�f������\������	F�(FMH�Z��]��Rb�^������=�td�6��o=��aKc}u�n.��)S;4�V�v��t�:s�)���]��f���4�=��s�9�q>B�#��L Vu�� �q�0��q1��Qw1f46bw(�{������ѫ�w���5�KQz(1��z�UGJ�T�$��:��	ׇ'Lw��.��?����Bk����J��z��ݷ|���%t��^>�����	'���TK��L���ko��w�u||y�����s�UՈJx�Pk,�|��J�T��N�0��DER��668G�3������[�I#S����F�F�`ɢf���E�W7NaƓN�4�h���m�U����i��EK�|��H����O�5*u���JF�ʁ�� �+�l4_� �Jf�*c�R����~�E �
�
xf-�'wYs�O�5g6��B�z�}���h���mEٵh�u�{�\9��z��%�������:�G��k�\_���h����ٽ���QgZ��v��٭!N�e,IgЅ��Fu�(�F�z�V�� �x�Q����YɣtON�Bgx�n%w�V��U�_D���H�cDm�o{\��?�Ý�v������pgG�W�s�� �C��Smrj��?�A�t����W��
���{��_�'Wm��*��*�vͻ~z�^z��K[��1ޗ���3gg82��t��(R�<��-����E���l�)��V6��(��K���w}�1��Pyu�lP&ax � >=q��v�W��#�����D�CF�`X�Vg���F���9t�ī�#;"g�@�ӱl!%�·ֽk&=�B�����c�k���H�;�kڙ����^���"��ȩ������~�À>:rj*���'�I�M�3��}����
a��g�I9n�c7{�Έ���}^������7o����߷�O���#����t����|F�m��i�<�dM�Y�Ѡ�~<L6�2 L<��G�}aaw��Q�Ao乆���$ƘF���(i!�/Ѣ0�\'��t�����U{`�Xv7�� Ӷ��owGt��|�Y1ډe{�(�+�3�Lx���8�;h��{�V�ma���	����UG�N�\I��<iFw1�
J�A�ƺ�z�v�{��K�^W����*�r�2���� ��a*�z����e��'K�<�:vJI@�8�\r�F�)�[7�:�fΑ߉���N�Ј4q	�jg�p��N���>����c�H0�X��@E�%HL�)�UF@����VeŦ�����޹���U	B#�����|�g6�mŢ��Єu���fϬ����x�cU��*�Qg�zU��;��@<�i;�g���&�hG���v0�a9��;��NJE��;T�����w�����?[��������{���iZ*󊲈��S��>ކ�<�u���Vy{<s�B(�֍4H��H��O��9�����:<�iOx>힏�ug ]�u������sY�g:�ex�^K�Uù|�I�<*)�X�P���
OqRǙ�F9�g�{�����_���
���Y�̧� �����`?�"_|�$�X���o�5��ٰ<�e�|*�ذ��rCs�>�G�����/o�}�	�3��:0��ɻ�P�u_�E����J����|��{�G|�����9�l����1��}(#Xv
dd��{�G��l��Oc�����#�^_��29z*�:XŇ�V��"=v8y� �/<�8����=z��A��9<8h��h?��)�ÃCxh�ce~<��FP։sJ�[�]�c���g�hyNNF����'� �v�Tv�9��$����ä���*�P�Q&X΢O�V�3��5�j�;��s�<�|I�i���a�x����K��4��oG���I<�p
FѸ�QƷ��3���Oœ�)0s�ydD�g���Ǚ=����/������]��C-����/�[���P�u+o����F�F�
����~�v�ؑD�?uOD��T�_�
>�Ϣ��R\j��$�����#�!;�-S�]w���<ϕ�A� r�L$r��7��4Wd@��M�5֥��v�-y���>�/w�C���Fwo;���x���i;�(���1�z���K`��'?M74��t';�!�;�Ɲ�����x�dw7����G����s���n���]{�槶�Qk��mq6@ %7�Ѐ:�Pd�����Cɏۧ������������>��mm�=
��{��Da'�wxx�s��vض0�6>m���o?�בK#�671n�WvB)#����3�S�=>��?�:��t��H: ������͛�o�p2�yu�RM�{;�M����Pp����-F�.F3�jc�D�Ps�3q�d�"��Y�+�2b�{!��ec��rO���/�<�Y��/7$Y}�@]����v�Ά���&����Ae-%�yx#�to0��>�$|O�鼕ߠSeWߩV�P�2��'��W�Q�>��tK�WU
$���O�:�D� '�9��f����f$�-�:˨!��ĳm���)�k
�A�����g��-�p+���v���ueC����s���^2�E^���`�]/���;|=��3�\;�(���ߥS����{��R/{�J�����H��ŷ����I^Qa4�Q:���]\isK�1�΢g�67�s���1=
a¶�������nu����U{&�)�8��=$�r��;0��u
�Ø�T�*�a,�E����1�K(C�?�U�$Da��U��S�2�B�����O�eA��BX�	�@_Q�9U�^�C;��uE91��.���(�ɫ�bWl���d-\ޘV�#0���UV*M�7A.#K����t����OoP��=�H�0P�%(	|`\�m�m��5�����kz�m� �L�˔?��y� �'��^]��b�������'����^��p~��"^����t��*�4z�,�s���|-����m��ct)�$��J�72%�'�Y7�-�.�_��/L����J�C��� �)'H���-��͜�/n��Ƣ�5����BV�2�=�g߅1W#�<S<��V�Bx�P	�ũ���@D��m��w���~���u�輪�� ���w���r�ן�뢧����2ʪ���y/xșr ����t@�A�s�`��y��t�s'=UC��03��t�O�)�<�.m��uN7m|b"���>{�����2U��ӧM�7(Co�&�'�4��p;o���ӴL_�����R�N� �#5�)��d�rk��LK��e����\ْ�����ʗ�"�^�ԛ���?iM9�#��A{�U��4�#����|�̇���i��]3ܚv��]BUF��x�5c(������i��K&\�/q$�g����W�=���=ԃ��˷���7<|�y'�5ڲ������)k�<H�6˝z�1��q���=�8Ne�|Rf�3Eb�[�|�}�/���o95����]C>W'JW��?'�i���+r�5|�N ���#u�>2�p9OQp!�ލ�[��{7>Xߺho>�{���2N�s,���Ki�J0,��q#k�Q�3�l�m��͚��Zw�{��-fѐ�)020xv7wۛB.����ɬ;���qup�y_��Fב#E�m}}k����������0��n�����E���G�fv�q唷�O;��ϻ���{��i�`�aX�{�>S�޾��c&ܶ\Տ���C�4p���^o�yX3e&�B��`G��~��c��k����0�t���C҆��G�,V���E�Rob|�WF�BZ�-#Ԉ��� ��1hs�Ra5�#r��ͺ�&'xGg.�O�c�����Z���'�ᣥL]԰�\�n�:x�����T���C�ʢ�C�R䥥�^���,�p�K��[�K�Y�kYx�Σs�m��0��#'����_ka���|�^8�K��u&�>��Qw����9#�k�A��k<B�ѱy�����V��������1��eO���b(#|*�X�au%Gʥ��5��"Ϗ�U:ǧ`�o���4�����"��?��8w�����Dv��$�T>
�eK���x�#����mj~�M�η��Q�z.�r7��w��&Yʌ�,�/��S[�C��;G�r7>�7H� �5.2�/'�]�	� @�U��0��GrU�����X��P��x��h���T� �U+n�y5h�1�:��Y5��,��{FVA��,�F�N��Y����&��:uʋ`TV-+Cf|)���:GNTVKUb0�\�.L�@]�{���g�����	V��F�J^͍w
���T�x 	V5�NF����=���R�����&�s���cm��G�C���2�4�4�0�h�5��1�r�Bg<)��� C�f�z�Ψr�֛�n$�e�j��+��4�:V4��N�Z�^������;�G��*,�{k�P�-���U*�=c��{M�7���m�`$f�qyM��%,�
̝���`��t F �?=u«�C�$��;|x_���ʣ�.�]�Sa������H�O�3c�Y�)�W�g��G��9���^3�U�hV�,���ƙ�� 9�8���r�=
&��˭̹��B7y���@�:���s3������ׯ0��fa������c���(2��j�9z#�uU��Ai8��?�ql�Ijdʬl��YnQ��<�(�4�1$;8�OЪF����Jy����}T麫�w)'�M`��҆��хA�G���Gx���%y�L�˿�w������LZ�c_��T�(�}z��l����}8Ն�ń;�2}�h��;N�3_.��|����B�	��\��C���e�|���	�rJZ�����n��n�������I{wY��e�PP��+#�{�'}�m����uｗ��g�V��	X��\c*����Jg�Xʫ��6F�J�8m�8a�69#k�C�Р�.�+8�{c\�<3"�]�,���] �1F�����#ksC��i<�(�nѭ�Q8�.��a��idM�Qv�S����(�	�H[^Fyz�֞>]n���{k��?��mC�?x ������Ƅ#%�0�is��8�&�`��M7Ex����G�>b$m��6c`mo�~?kz���:�ȕF�O?��(�;�cl�庱�a�i��S�Ar�;��#�TN#������-g0�ݝݬ�������Ț鯓V�5��ã#��h�Ȧ���P���ɢ׬��OƑ;G�45�ΐ�J�Z�"�[��r��<�8�A��Qwփ�7S;S�I;==���oڷ�>o���8�B�Y��5Y��?x��vF�3�,��M�	�U����,G��Aԏ�%�J9H�~���`�Q��i\gm�����*q��SH|��j����fUg����ŕt]cgG@�U�y؞e=l�~�0r�	��	x*2�|�8鄄o�0N�<�1�^>��gv�(���3:IEZ&�N`6=`����1Ȓw����w%������$[i�� ���}���?��0ʩ��W�EZU��٫�j����2G�(gg<R픣�C㓄k�`�z�5Y�����m�q��ȿ��������(c�:���,#K��&?p��.�.hC�N[�(��W�Q�TdG9�H��qG�l�{!ja�,+U��s>�r���h��g�����F��]�v`(g幃K?��tAG����H���BH#KA�p |od�<��Pa
� g�+q��	@��}��s���C�u;�����۸�x���?`��bH��{����U5bUu���*nY�.�����n��P��eJ�#WeP��n�,G�4��j�^�e��ǰ�팥L	��r*�`TJ�@�5��=��]�|�,��� ��EGD\A`piK��сb�^�q�B���
�.����0uil�z�rUY�����
�q��5͔�Y��$�7/�gl�M�??�e��zj9C4u-��s
�g�)����ۺ�}�͗?��[p���+��b�}��w5�U��@ɢ��&��D�P�»�"����1���u}�!�8P#�z�xۆe1�Jz6P�Q���^/��%�n���I<;������?{��i?zܖ�g������7�Pb>E�s)���V;i�$�e6P*���W�dū��=\����M������)���L��)v�:{"�`�_4]�� XԦ<�(d��~:����ŵe��S�$C��H��)�ː+�,^����+)������
K6F ��W;���g�QT����l���^~I)���B�hK�xseW��Xχj�{��\b��\��_�^}G_���Z�7�۽x����5��YG�����⼎��U�]�+ҵ|�v�n��,u)���?�F�Ϋ�Z�����΋L[��"��ʥޓW�K������b��	�r G���Lo)#�LC�3��)��(������	�\���u�q��S݆�����ؿ�8ή���yy�:+��3t�R�h��x�xl|l�&\Y��:��ĸ���<����1G��O�1��*��~���o?|�=��^F��¬b�����xG��c��ۜ��5o�%o1�4���0�0����G�������������>ai\��r�F��E[Jw�Ȥ���~?�R��u���61��?��o����۷����g���{G�0�Lw�2����r��hx������`�AvB����%��]d����S�NN�-G�5�]��SN�g���3g��H��Wֽ�1��LeU�['g���%�.�_�����[��Gmqi&m�[�������S0�L]�C����)`�J��85�B�үtꨫJ����|�h2ȵ{�����P������W�|�\��Zɑ�t:ȏ�eҴ�UlQ!�vq:/����-�3R( W��2�J?�S P�<w�:��%��T�+�M�{,�/�������i���w���P��]A���rur<zU�랹M;����O.���i�A�������U/�̫��9+���{�5������0`�^�^�^����@�B�!n�u��l����rTԎϩ{���r���C��m�����Y0�s����D17��n��tPB@�4���t���==?CYw��n�?�!2͈B:���F\���ɂD�FB���/�7�I�!�#S��9�8�!x�+�)��HX�Km���� ��P�� ���P�ٿl{GWm#�茆�@C�r��j(�+�	���kXv��w�c�s�E�z��ĳʭLC�շ6#�D�l��h�u��`^�) �Ƿ�3�+(�� �9FIs{�!����!\�W��k}U���Hb����K.�4�0�4�N��Q���l�]���vu�M��|���m,�`�@@'m�FJ�����S��Q��~�S�����X�o��L�k�9M1an�TC��v�bxD�� ���ǘא����І��x�Yq(e�!��\���4Z ^�VW��oy��tL*�V#S���F����I����ОV��\ˠ�VaH��t�P6�ݹbt�Qq�>�JR�B
�Ѝ�a<h1dE����Ȗ���@�`p��Jۯ}�ɍp����w�~�]�-�]���������:� �5�M�⅔���9�6��
1���7=Q����@I�p@^DIt+�K��|lĸj`]�3J�ZS�̖G-�F�{�i���Lg���/��>i�8负s��-�O��Uyq㌡q��ʚ���o��.�.�`o]�Iكc�f�4e�;O�iG�4x(�Se�C;r�&Q6�ɰ���V����+dhC:�����1��ihTFo�Y��r���#�qw��ʽ�P�C�d�"v;�0t\�o��zCyI��L��IE_�M �G��]�t��0�k�%�o�Lդm�.����+|BJV�ԗ� �o���
���Q�4�Xr��"�M�w�������x'_)Á?��O�;׻������uW����핋�[w߻j����i$OeU�Ǥ_�Zg���!h���F�r��E~#�ON����Ƕ��E{�g�6r��0p YBW���+q)�O�Z����PY�m� [[~/c+g ��[���2��g��h�|z��ֈ��{�i�F�з�h��1���SxU/Oem�#����ݙ�ClG&y�L&/��G�A�k�#�����������]t��v|8�Ngh�&�ՙ*Ҥm&�C9<[��
���晩^xG�l3=`vaz�=\�oϟ��'W�5�����~�������z�en:p���wD������o���ƒ#S~��O�b�xr~_�7�=����4��S<�roDa8y��9xu�ᤦ�i��D%�^�!�{��EwvaD}X_'�Om}�)�o�G��m} �=Oԇ�40��9�����	�aFȤ!����kt�Wmqq�K�h`��~/�V͵kȤt?uEDm�v=rK#�m�o�74��#�٩ɶ07ۦ��8�G�DGy�|�����_����U{�2���Mڸ��m��7����}����޿���o���	h��4��?���I��Nq��Yn�,C�P�.��9k�D:=g�9f�\CЊ��0��ܫ׸��hy]�:M�fhc�W ۷�-wf�\yh��필M�'�gr0�,ظ��k� |�L�WV�v8&G0z��6���в��'�{�0�`���/�_���~���6�c�g+�y���p��#ˇ5���щ|"��T��v�Ns)Ŗ�:`ȓ_dZ(Q�T�)�}�կ9�M�#b��e���X��W����Y�^�'I�
�X����'�	 �D�q��"���X�˨���x/2<���(uw3:��4?����ǅ��:��ٓ�`y�_�'S��Jfb.��܌���	��"+��k���[QX{��x�~���$�X���� �y;5`zz6g�LC�1������:s�u/��_:7���Q�Q૨|�����h���.��}��}�׽�ԃ�A��?�cRR�$B�beS���U�v�NzELt���/>���WWV{����`�|�����6�����B�^��
/�ܨ�n4C� Ì�s�D>��0��a�^eC�b@ѐe4�2|�����v9��*^8�vv�y	ׄ��0���HL�S��2E<�� ����u}����_��9�p��V�`%R���E�P�{w���zJ ������	W�*è�����{�.y��?s�k~���s������Ƌ�<��{��Z��쮜��9s�U�C�ڧ�^3��@�XD���Pמ7t
~:]d�
AzU�'���3+�>pf����>E9��M��sF�OZi4�����yNX�����T9��Gw�H�������+/�3�'��x�2�^X3�!��q�U�иCp:��"��,���}���`�!��T�ܜ �I�A8��r�2e��,�|}r~�k��#{�m�������Ƿ�����a�Cz�%O�+9Ű()�Kg�t0@5��=��:����M������=站�{���S.���Xx"���
j��~b�`��}h��%r3�Fvh4�p��ý��pw�B}v���X/Zs]��������R9��R���=i���lO�ݞ���=�m{��[�m��}���h�����(|���3�9��6�������/۫/W�tT�^
�_�+����A�)%�/�^��+�?�1��\��q�Ai�U�2�������#��6����u�
'��Qc I�4�)̟D���:H�|(,u�xWsJl�Ά��ӹs�F�k6�?�g
���!�r��y+Ǝ#A��?%�leN�,�4|�L��D��mU�qų߲;�����A������U�r;4�ww
�cc������C�h�u�i�wp��������^��D�T�I~��1pS0�'e��z�����~Ѡ�T��~�,���Ô�	ߔ���53�.8�+P7�v��Ӱ�Ѧ�
�M;b�_�sw��S/��κ:s�$8w䦇I�M�|!1��o��ʮ}vT!�r^#��٫r�fU�w�?6q���6l
���
ݦ��_S�D�LG�x��ep�NYD��m�Oy-���h�y�B��	��,�]"S;,��X��c�7�&������)�HE����<�a�-�<h�����յ6���5��C�����Vo�	����D��|��@��$�]����;ǃ��e�>�x�*޻{7��q!mi�b������3��<���=��k\��v����.}�G]�g����$R�Y�$i���QWE����"*�QJ� ��PT1��/�#D�.����Ȳ�Uh�H�빔�Q?33�u:�Y���@=�tև��L�:�󾴄����K���J����>��oƹ�\n�9�q�+��&��D��� D����w�������рı���O�	'B��-쉻�?���O������t�[۩�l���O�M�k4�|�x(87�0�{އ���x[��,�0�`���p?�f�"��E���;f�V���D�UB��kt�s�A������1��8����|�]b ����J�\�|sn����'��4 ��Έ�`FE:�RV��7u�=O)K�l��/���\_�\��1�:W����1i�pPX��������.�]�Iu�s������D���o�����}��]�q��Pw��S�R^��ܫ9��>�N������PY�W����H�xjaG�-�:"_��*Ҽ�=ST`�!�m��dc��o���n�%�1
��#o��Ļ�"q,����`F�C[Ri"{�,#u�<R�<�V���ė��>-��F^M!w]��ۊ�����LCe�Gj�0�}5@K�+Һ����'�m�J�U����*wÀ���)��H�s���w�u���h?�%���)F����v���u����q{��S١B���
l�����|�������:�Y�|���p�H�>S�``��I�W�微_�JC�QqV��S?��	�3��%oL/�^���!�>>�k�;��>�pwy~֮ϑ�Wԣ����i�3Kmvq�-��D�=m�P��jO0���������_�՞<���w�g�l�|�V�^���g��M`p�a�����f$J�S�s�S�]($�>e:����>�����n�T܆Ε	�{��C��OǊ���^��[^�z�S������I?u���A[�O����Oi!F�4!� �N�+c�~���)őG��ȰW�3s��!kf(�
��C]��c]�O�w7�5�u=�12�.���V�4�5)��CȚ�<���gD٠�XvdO?�w��!G|�u�$��'���W�	{@�t���<�0���9��3G���fi�͟
�2��7���);��Y*�҉�(K�e�ޣ�a����gӀ�~e��d����N^j`�rTĊ��A�hȦk��Z���Q��)H�!�zՑ*�����Uޜ�;P��L�~���3!�'B�R#J#���l�l#4d�Y��5k��Z������N;���]K�vL����FYf(�s�a�a������A�Ț��;��FV��8�)3��Z
������<�:s�|Vm��<���
D���gG̖���ö��I[\}Ԧ斨i���z����m�|APa����ˇ�뒍]�Ȉ�{�
n� O-ܻ��!���G|_`���k^��q��O6Ɋ�-1���[�nhb���ϓ��B�]�g�X��P�մk��!���|�*�@�B:��/��� *�"��{N��-��ڽ5m�Yz�!�	{��]���IyWʹ��y�
2+��Z�ϝy
�Ť�u�o
܂1��?y������x��g�֊�\A��S~��u��
���0	�k�K^6���t�=0�K��'tnd��!����ʋV��`��iXiHma�|jW\/�1��X7W�ꐶ��~O���63y��gF���d桯=�kkk�.������å���� ��Y&n\=�@�dN�ϼd���Sz� U�igN�e��Q�E���]{�օ��^�4^�Q�sw��{��ݹ[n���
,����<���UF߬,kSaWBH'�{C:S;CQ��� ׄ�8���W]U6%����V��o:�wt6�O�|6x�S�t�����z?�.�𩒖�vAC�=�UB�p�]]"��#��t(�̠�c,�G8�UP�w��m�&h�7���k��M!��B�����;�����g�
J{�/��T)0����_|<H�rPG*
Z��W��ƛ���FQ<� ���G��ϯQn�PnP®�Q�U�J�iAz�?�s���!~6����rh�2���Ȗ�A�g$��L���;Ԕd�Ty%m�<��Ƹ"=�'�x����]�@�m�k}���w�f���|ҎPtN2�	�G\
1��[���t=�鑆§���]�����n�m�;����<�N'�o��/4檂lT�Ls���ȱ���m�M%!��^�_���?�y�]C�m�2���(O͖�M9lKx�W.B���{;�\��V����܎�#]k�Q�8�������m�ɫ���+�_�����Z�a|�\����_z�p�b���=���{��件��+�.�,=�x[DQ��Q���h;�R��;}UcĶ�*���RH�����{Gv��ԫ*���L����8غ�^/��S������9*ݝ�B���Q[�őeh�ؤ)d�!^��l�Q����׳�{)O���HGY0����Oe�&Ay`|!/#��P^eMvMT���3ƚ��ָ&���%q1���4��wڒ��ز3F��Ú���LC�g�ݺE�J)�U&�R	�N����q�Ɨ��������R��ز�W%�)������#=3�aC`��7���S�"׶�o[Yפucd��n1H��)�
C�qE=kl�T�2�)/�t��Jħ��S1�E�e6i˯�Qx��G�S���Þ͙��>�髱TS�<*�J�:s��2¬��^�Vdt�f\�8��IÑ�~We����F]f��e<�E�a����ǰy%���kћ%�nXi��efm���hp+�&g�,����#ףs��>��*�ړ�fn��.��/��گ���PE}O��Um}:^���'���˰�,�I�¤�n�t�{o����۽dgˇ��_������tk�05�t{;1���v^�w�G���L:I�������#�z�L���$ q���'���	�eDR�����#���"D��YV�i�*Z��e�뿄��"�C;ݳ^�E^C`_8���OAa��8��"�}o`��
���A��YWq�'�P _����$���<^<��W���$W0��cx�D��[y0��	�	����׍vv���S�����.r�(�'F��������x�+�����GK���E�n:�Ҟ<Ym��>X[j��smv~ztA(�z��E�MC��"��5�e�}��W��4����@Cp��blݜQ�2��<9F��WRF��ޑ��2�0̲	�lԹ��5�qd�%k�~Z���Bx��rU�X�6���+��[_
U�۸��F*]C/����n���g�_�6���f�G�����`
��1.�|�3,Jњ����6\�����r8a��ݟs�G���K9�ǔ%O���m�
.��P	����ϰW4�����M�g�(B|d�?X�\�V�Q<� �-��@�v�߼j6Z�VN��S
$S�e�"Z]濓^M��`J^𩽔���ҁ������]d����=�XC�4S�j*�F_�)�J9�O#�� �x2d�
��S���(6�R�͆Ru�^��8��'��P84�n
�G�,aV������J^��y>�Y;rގy>�l�NsRw�.k*$8�����M�u����v0�>���m��ah��}28Eީ�y@�FC,R	���GS)�V����[/P�;�'~qF�Q�o���n�������I�\TKu��I	Z�c�wڤJ�rH�L;;�o�����Ƈ���ᾛ���(â��L��������=\{���T=~�-F�Wm��3*�ٕ6>��B5߆���(�K��62��&�����S�W\�`d}���U{��oڳW�jIki�)ry?.�)
;0hdit8R\��jd��>_RF;4�U�U�ѓ�3���ăjh
(7�]������)�G�m���mû���$�ܨ�i��4�z"o��W*��@��

w�(�zp�����x�8�hdͻ�eq!�f�3e�^jS6�m6C������Lo��S��~MX���G}3���4����0��	_:T���)����]y�wzeOw�s?Z���\W鲎�����rz^F��'��c���L�T
t�y�=��M#�uoN9�-T1=�\sݞr��|8r�g��!�7#���
�e�<e�� p�Z�߄32�4,�xT?v�C-]7�:�����ҡem><�̘z��c�$v ���3�w��r'g�$�fC#HL����c�t,��z<��}F�xg�;z�٭YYH\0��Nkt���8k �����������������w;O�uS0��c�mfn~^����=3�d����dH�h���]tx
Zm_�L=�7�� �Fʗ�w��O�LIl?+�2��ߵg}�~0|����}&�;D���ǐt8/#�Q�ȱ�q�>9b���oF�1�&���d;G��ٮEΈ�Zo�	v�@��������m��~����;�D.A dm���,��S���ƞ�a*L$��k�?q����ʴH��O=(�BĊ@�4�T��[k��<e�=���n��������Z[Y�oS(�[@�	M���ɣ3��_���۶�{��r�y�x!�<�[�Pc�^�J��?I!.7�[}^�W�'���V���1�/4H�P�*�V~���M�|�4iDs5���2k5�N���:��Z�dë1┺2@2u�� [�j�L���ٚ
8?W��g��g(�{��^ů,-��%��.�E�>7�p�x�x����mȲ �:��!�A�k�TiJ_Lc��NS�`%dn��
S�Mz���f�.���et{������
.����{ϋ��>�Tр!t�Տ+nZz��8�05ƭ��#�����+(6䖳�ߏ~���-C��g<�M�W|yM�A�J�n�����Z�>��k��W�Q��1_�"y�����`��F�����W&���S��`�?�_����_#;�
�:
��@+:����  ��IDATS�Zm ̺���T��+�����r19vrz�vv<�b'۷EI�!M��-Z��Sn�P"���g�dh&���F<�����Ep��e��� &)���8�4W�+,���y>T\k�+��0���5�`�PJH?�0k=��|����mrf���/���D�\Zm���(�Km�)ES��aVyu�%
d�˘"-!���2Q��E���W�ݶ�59����\���n��'ɏ�I \)/Ň���^#�"<s�4��ӟu]~�&]�S��O��ϝy��^a�_���507��At���Q�6y�R�L?��¸z��?�k��������N���+N�Z�^V�\_�=x��/?��V�'���OY�N;�ڢL��S'�ц��sUq a���(���4�d�
���h� �@mu�G����%�������tY7?�S���4�GuƏ���һi�<�������Ë۶��>l�O;���d��E@����PE\*��~%jjf^�̴��$_ؙ�X;��Q$vH,,�e��W_=mk�C%��C��-�7?m� �cG�נ"|�H�e�9��������(�F#�nP��|����O�R0�Ћ8-�����RRV;M3.��i��/aL'���	�Ž�3���d��:�z���Q;Ez��3V�����,�@�Qd���8���?������C;:<#G�	rɱ9���Г.j�pˑNYG�albQ6
�(����N��Ϧ(����O�s�@���H4������X����v|r+�JG.]�"�Y�顼��K���qd=P�f #@ܿ�S9Ҥ���AךκQƌk���
��.1�OC͍i� �n��mN�SWٹ�r;{'��A�;�v�N���c(B�F>�p��]y���xq@]�.���$uW����f��;}������gm�vN��}���=ێ2���8����ЊtX�C�e�¶��Cۼ�^��M7���5��i��4|o��c���p|���|_i���B�$3��]���ׄܤd�£{*��i�c�V��"ؐ�7�Ge�l�����LY5��t�G�nx�ϟ=y�^<}�Vё���uNF�G���M�,��Y�Xu&��<-P��=V�
I ����P��mYK����* ?��h�"�,�zc+в��ϡ�^A+�y�c��[P��@O��5��Q�I
�.��`8�ՉF��U;<�n[�'m��)-���� {�,iH�p���"��@����ʪSJ�}�<���������E%���e8�k4�w �bc/̹����N�L#K��u��Vn�^gR�[�u��GW�Ç.�^�N3VW0���F�~q~�-���s��y~n6�����dj�1S?��C+C��7B��Ec\�{�sʃ�I�Sj��z��[��+y@��D�d�A^
,�G?w���kx��et���ԣ��������妯4���ŉ����_�U��>'2��w�y�%����Jv�']�,������y��ԓX�;_�qޗ:w���[�S��.4wy��{��/��u��x�2ܔ+ȏk��2L��LA<1�&2Æ���6P����
�������*<ߺ���6�҃ƃ;jdI'E셾0�W	�g������/fK��I�?�� у��,�0OG����#m��֯>�l�,q�a �Tt��C�c�[��6��7�7&Ai�_�������q�Qۀ�o�r�֍23�q����e�eh�1
ޢ�Z?�!/�A���b[XBƢ����=y��=ut�U{��%J糶��1����6���&��k�k�*��X�,���S���'�� ��~@�2ʦ�F]F1�o'��읬)�¬�h����)������q0��CQ�g�߅���>���~��7ė������r�V���7��1z�r?Bݏ�m��^���㇟�۷?���_g�����(GƟ�n>~Ҟ<{ɵ6���_n�s��9k�+T��W��ί��rr�P't!%�A�W֣��
#��@9�8=�r#�V{�-� �ã\)]6�_�_���/E�y�y x�2�:�M���f��_�������A�=T!�D1�pw<��Uu8d����Na��M'����c�zf&�SHҕ��(ԓ9����'��+��J)t讦��f���������u����4�\��J�,T���4n�.��� �#��Xw V��Qh�3E^Iv�EY�Ϳ
��C��z�<y S��4�s�a�3��]�x'�X_���,��8�R؁�=��驎�(~T���gr��ʊ����#ȱ��h�6����B����CW(���/� k,��Ny���8Eѩ��Q�g�x~Fxp,�*����E�euu]p	Y�h0S�+����m���rD�n0���Y�i�|:����)`?��6Vn���T���ѓ����i`z.�#���J]�*��e���i��#�J����*�8���ﺫ�6ɽ��S����պЦ�A͂�P�1t�ٶ�si���S�.H8g
I���%x���4&<v<A������˗9�@P���r��gn�p����jS�AXl��J��Jt?�J���R��/ᡩt,`��x�Gкv��y�%-�x-��D��y��g|��۴i+H�3K8�~�3���it:ޝv�d�B?w�k��3�x�+G�ҳ�:���b{��vɣ�<t90�����эdyN։�!���+l,�F�#K6�
!{��#��l���N�x{u3UL����XZ*榕8"��>N?tyi���S�#��=O=���H[ń� �acc���u��u�a���s����='��֖5�F���@�U8懰"��k*��dW��T���;�8uwgd�3�t` �`���ŰJ�
P��CطY���z�����Q��r�������ֵJ$X�2,�g����e>���� ��� Yj�0tXmqQ��E�U��+���i/�]h�!V`K�c�L:�njT��*c+[��@�x�����Ʒ�C��TT�3{i�:����4�NǠ>y_FY5�}�2��ʯ7�¨��/�.D���	�V���1�1�M9�C��g��K}�g�SOC������q��;��s]�����;��mbv�{����ƫ��?���uo{ �\��Q�i�La(�_�&�x��*6����)ȭr�uR�q�F�FV��>;e辌,m���H��u��~=�.�I$��4b}q;I�477��i�fh��3��[���zP�n���L�F��rˆ%�(��4gMy�X�GYBx�;eVx��a�Q��ec�[�����}�Wг�Tނ�R�Iy�����J�@�@ ��퀀g��wtDjfv�-,"[Wa\=�!���i[B>,�=�ѵ���������r����ն����Pd�PP�\'��_}��N	~��$
O꓊�O��l�`�=����2ڛ]�!_Y�.i�]>��:����7��;�H|���x��?�����%��p�J1%(�XP�C�rTم�>��l�6�b`�n��ߴ��u�C�c#�"8?�=�M��}��Y�Ob$��OCS%_�yfkh`I8ΤP��@�� ��T`�{ ;>w��U9�Ȥ���U����k�`�Q�}�0p
�2��o3�si���$0FA�.�3HZ��w��W�K}�6���90�ߴO{�b���#t���vq��U�:���(����'y����M��kG�4.�v�N e��W_=k/^=��Zojd��������[�dk�,2I|�dZ�BN��,Ӽ���T���n��s�i�RD��M4�j�Ӿ����1���vz�
��.Y\��dN<����Ǥ�)g�V��z���-�@�Z�a`����39�v��bp�D��=8<ho޼k����9�8��-��+������G\�lt��F�0��I z�F�#։����1�O +��F�O&1"���"�顗�@��=q{�ϟ��V�c��ѯ�.��i;|�	�I����@y��+�����J{��Q{��I{��Y{��i{�TGZY^F�-d�y�--�/�D�	�^��1y=\�?�HG>�Ki��:%l�8�g�4�#{�pS���V{H��ϟ;2XC�vʙD��t�ό7������U��9$W������֫�����]��x������vv7h���]U>[G�Ŕ�x�SS�K�S.��.[��Ç���U��>2F�}��v��Ix��k�Q���T3��o�=��*�=�:�\��\t�� k��T��7�V��x�wBǍ���*�իb�yu`����1�V4��F���Zw$k��mtA`�@����22eo�J0���rL��)a��2Z�p�C%X��VA�����=x.��KВ_�)�1���g,[����՜X-�����(:
�y�`+�y��uY���,�0�"c�_�O���D�����W�B�յ��,�KQ�&�z�P��`/o%����U0سR��zExR�k__��=�Y��q��~�*�Sn�T�6
Z��Pv�YYumՓ���s�S�£��-����sn��CÇ�y?����lzf�	�u]y�W��=�S�=�!p{,d��r_���k/C�ڀ�#[�;�0����� �k��!F��XO�(�Wa��f��/e`uP�.�F^�s1�\�KOzBt��W�T���p�c{gZ��k�F5y��p)Cn��Ty��:W�\�a��\�+�\���W����}ڽ�i���޿v��eޙZ)c�0�9�.��O��NJ��id���l�_��,���x �=i�1Gٹ�1�,�#��v
HFD��d#<�����4�/*�=<��y����Rz-��@���N$�?8LxaFӍō=zZ1v�H��cE�fn@�M2��(��Sq��Tɒ���0��P*�M�CӔӺ�=�9�D~�!��]Y�)����mN�6�.w�����PZlKN5[u��Ӛn��������,J��"�jfv�M��#0��S�v� 0�V�˫i+kx�
�u��=~@|;���3�G���̺�w�3�j�'�p:���RYe��WѴG?��.�.��������=�B�]�Z����p�c���`��t=_�^u����	�Q�mC��b�� �/���1��g�n����>b\mm~h�]N�k'�M����x��:s���6�q��PT,�!t@��: [�rq��� ��2��X%E���*~�M���a�)~�LCN[�ˈ+펝z��<�,��]���ʚ���n (�k�"5�2v*���uE��P�w�����Q{�qH�~��.��m�
�m���&iDq�1gG���؁#M�~H"^����O�D?�����#xcĈ��j���mow�����붻s���ARt�6~-�v�u�vʹ���P὆)e��]�]؎١
�O��!��&6�3��+}��=���9��:1�u��D�#�G��H��S���I���I�פahdC��ț�����C`��v�QqN���e���]y��m�h@�͈*E"����&:�G����knC�ݎ1N��]{��D�p�x�7h$��oc,�����hZðq$��Ed��y<��ɓ�	������W/ڷ�~ݾ������W*�ۓ��1Z�0�0�0^VW�����(Fܣ�5�<i�^��n��@�^}M�W�_C�N<�[B�2ߗ/��W�G?k|�?z�>�q��i{��%��+��؟�\�̹-��(�@z��I�õ��>J9)����V_�K��Wћgl׬o���|��� g�����vx��6Q�)k��a�Xq���Ȓ��ue7(C�yy�$��]�F��y���mK��7r���B�g+3���g�;�K�$e��&�f�|r��K���VeA�8=�k�`l!�3�:2:u�K��|����.���cL?�nV��-�ہ���?�&k#K���	A#��h�:�� ��HL����%�%��A,o>=�\S����4�D�ʊ�`fRH��4���#�i)KQ��cd9�bW{j-��o*B;I�ڰ���<��:<�j�����3������O�f)l���)��l���8��ji��<�s
º���:+Q��5�w��+��T\C�3��=�4b�)u�m����L�YXn~q�θB�*hI��b]�k/�=<�_�x0��-K�+�u���ϳ�L{�g���uSm id{��x*@c��:-�CO��k�+�S88�@��A����f�tyg#.���F�ђ�T@e(�Do�Ks�Q|��e��u2��[W��=�hJ����e��b��ç��Wh�(�(���I�K/�'x��"���᥷�Z���r��A_����ƒ�_r5�4i���Ժ�W�	��R�M�V�w�b,&�{��.~���4���S�Pq�y��3<JY���F�^��R����krV�V}��òw8F�tOeX�v�&�j��V�F_ڶS��S>�?{{{m��S�����~ʮ���eqz��l�"-CsW�4
��n��g/(-"����Q��Y�Ebwf$+�YDT�uj�����t���e�!P��؄L�G�Vv:�etO��%1��Vr>�C��G�Q�מa\�H���r��Š��Q�>�-�3��]�&�	ӄ�К�qZ�SW����ť�99�&�2}�J���˻~�^5�4���P~>��5����+)�e�fT`��i��Ev�S��-^5�Ow����/�g�⺋�[�n٥���[��͏8Gx�n��a�(ʡ���n��Y���mkk�}x�����{��-J����9O��@:}���ڣ'�2z��b��3%������FFޣ�(��\;��O~+%Eee��8��>=`��<]�Yk�U�0NwN�>��LS#L(_�v�rG�1��X=�&�<��ώ�9:���z,�`�W6w�ۇ̓Z{���(��(���϶G�[����ݚ\�Mgr�m��q�%-�G޼jK�Q��z��6�<a��ҋv�Զ>m����}�S;:pƈ�O���[�4�[q�4<��rQ����X�~�N�kme�������D�C4��P��O�i5]�g89ʓ�g��O<�{��}�wM:vlY��H�Jժ��;�����V�g��菛V�Fi~�@�����q{�a��~��}��&o׮����I���d,�Ҵ54��[�k<�BSD�$�m�(ޑ6wϼu���Q����1d�k���A�&�r�iu��+>j�}�uF���<Őr������"
���/^<��5J��k�|�����7_Q�/�G�5��DZ��z�����`e)ZfXa��O�|�K�����i:���o���0�|�|��q�^�����0�^��fzK.��,G�����<�dy��E{�������O(����Hۑؕ�8;�f���?�*yK�sŜfXg�}����μ�+ea�<!��"��+����H�bG7�u��f��LT��ٹ�s�+g�����\�����'��ߔQ�5H���d�ѳ'ӠG�y��L,�-gU]����h���8��5 P����=#�5��a�w����u������f[��������n6vVG���s s��h#�4V�d5���OzJi��a�~WP{If��sf�a���$IDD�;dOZiD�07��]_Ὅ��U�A���EX ]����)��E{��6D�D��C��m�xxr֎�C�r�� :2�$rG
�$Oo��rW`K�]#/R_���I�i���9e��Ynx�z�H�wo2I������	�8J��~�@4�Q��r�=�_�g�v7����,�F��i�k˙!t��ϟ?��h]^Z��մ[�"��s�K165���S���E�N�X�s{اP
�܉���e�M)@�Ӡ����v{���:E�%m�4�n�W
Q`�t�ZƤNm|�mv�ъ�p��*�D���"B?^���5t�B��b	.Ŀ����m���1��y�H����~�(��f���^F����d^�I
Q�z���I�"Q��H�7�����5ګdwμU� /M:Q�wR��b8���BP����Q�x&ρx	%�}��^���+���e5�_<���DP� �\��y��Ƃ�S)�H4�P7Llʪb�s{�t��p�$w�rn}��.�A��L84���ng�rJ�Ux+��Z��]XX�����gg�����?��?�!��%GRT�M?J4�[�4.��0Q�/{l�v��W�CO��951zӍZ��(M�i�I��	��Tk�N������zG���FA�q�8��TA���+i��f�l�ק��iG��B!_}�����>�?ǿD�xƷ�661O�x7�p͌�#�V��V�Ӑy�@���D��~�Ϸ(X�T55��Kȑɰ��F�#�O��"u	�R��:#�a��]#[N�[������Q>w=Cv��%r�QPZ��%�@5>��1�^����#�0������=ϻAаMg����_�o�I%�ɍ8��Гpr��������?4�GN]��˓�v���~z�>}|�6޿n�����BoЩS�GQ&/�N7Ȕ�/���/���jƀ����fN��x��$3=u�O��^��ܱ<|�W�y_x�0T�ҫK<x0�;�6�lF�M@A�������J����^)�HUFڜ@�%�%�m�.����3h������H��CfSmw���y���}8l;{���l��]@=c��P�CG}o�/�pV���t=�Ѱ;�i�9���a��̡�ԧ��v2#OQП,���)`�i�G�mgk��y�S������C�u��8m�S����F��P�m���&�En�1�����gm��"�)ΑQp(���a��0&n��mf�����n�S���ap<y��f&Q-P��q��3�.y�����e�r��Vat]����t8�ܙA�wJ�$8��F1�'�~b0����\������i[�����D�5t�R�̶��o2Z����s���c����.�	������J�㌂�����#���O�o6|�N�wzz�w�-�O�"O���N�b`�PN���H�Y�h�+������F���S���v�4��|�ǉ��f'�q�来�T�!���������Hsn��Y��MN��~`�1�u6׭�_���V0��3�lya�-�εga�-���3�h�f�c4���*�����Gȁ[ŀ[�?^s��j�Mk����',OA�f@D=^}��4g�}|��mm����-�3:楝��$Y��>�K�(	����Ta�U��6�AR�t�~���/��)f�g7"���w2�NF:w9�N%��"��]�W�╹��`WM�y�6#|tB5����V��M�uxh��<�6�T���mS��[<��������g��"|p�K��m�_��YA��n��;��@!P2rD4^
�ڕʑ,���qQ��=�QlKɳ���ȴ6@�2��n��P��vz����tROU�R@0��f���i��Z�>���H!^�"i�H$�.F�Y�X�י����u��'�1�bP֊�
�"$"�������+��\�۹�c�п���µ���VE�2J(��^�8�����&���CW*�n�.�PR��n��7{�:��Ӽ���:�w�^z{:4Z��š�Y!�H��La�#!�LT$V	���B$ڸ�-��0��|�Γ�8�[�@:[�°���L1z4Re"{3�k<�����S��)Ј�u#�c�iEC|���T>P�S֤-W�%Wua��W�x��/~�R_��6�y�犓�Й�UO���s�i�c�Sw1�����ݝ.��T"D�$~纴/ȨKB���/���C�җŻ�������>��R�[�5�E��NKٱ1��
�J"i'.b.�����w�i������Qe��[`�T�ǭ�2=e�S���\�і?�x0��ڏ?���;����)�6=����ujo~�,~��]�1�X ʟ
F�V��q�
O�Y5��3��I�{�Kp�@fT��<l0lJa��N��%-�������/�&O��^y�֞��?{�=��Z~@�Э���ZhY<���Z�YB��[�fݒ��>��}�W'8��k]�W�Hd�<oV�T��}}9%C#�u�d(�Νάs�YC��&�y��W�(�����j^>��kp��;���$�J���|��5yw��A��/��y�fƻ[�%F���n;��l���Ƈ7�YX[*�n�~�G��ԡ���~E֙����5���>�N�n�܆5t5\�^�:U�x_x�]���L��8}9�1��3�y�����K���.K����#Z*��%)����p�MsTٵN�z�����c6R���@)r'���ms����ҳ�0����E����fV�c����y�(�7:���bISn��&	kW��Ӈgc0cD��?�~��}�����4�#ϗ�CQ����;=/z��C�R9:4K{kG����/�!o汇N�c7Upk�i��,��/����cHծ��á�%�Y�I���Əmau49���b�2W��s�w>�:Sn���:���ˋ���l��wi�rzX�`8�R}bn~|�vt|��~ض��(�g2�c�4�OW�_hh��g�����'�t�L��1�T�C�[�����_վ��Q����ȑ9��.m��i��ck|B#9�,t��Y�U�PTF�{�G�`X�@�9�F�
��_}/9�!�t���Z)�f�ge��� )G�~��N�b��.�Sԗ�eYrr:�u]08��:M!y�m/�m*�ڗ�5�bY.���w�:Vup�5���~����Ց�QM������a$o�����#�9�L#Q����w�	�S�����z+�3�w`����%roX��_xɇ��~�	���t��ZR�8v�G�$t����a�4��C.���f�����LJy�7pj=;�)>�蟇W�Oژ�>F��V��i���wF���3�"�@��^
v����<����6D};wZ�r�;ˤaf���b�sj��l(�ȅ�X��
���Ʋ�V�]�[��GY+1���b+��Y!Q,.��qod_v#Y���*;� ��x�TU����I�R��W��Yy]%��J�O	��X�,^�V�
 ��|�l��4�4�(n������Wnr��8@�"�N�����P�WI"�k��H�þ
̥�Cvn��D�SC+�l@m��m�v&�,<�������(wה��mzf6����r��I�#j���G�3xd�
�R��>�Z�<�]�K���\eb�0�8�I���x��|�C���2�����������͵�Boh{>z�+�V��5��iIc/$c奔^@}id���+�.����.w\O��e�����^���^}��w�z����e��ĳ��gz���
S<ӥ��Kw����T�>6Vrǩ6Ҟ��z�ΤY�`xyyEíR�A�#n��3����;D9���/_р?A�YMϻwo��ׯ�ǏP��K�A?�(]�fᏌt���'�C��24
*o������:�f/?��u
ԙ��*!4�*��t���>(Zb�q`o"8��JC�D.x.��ʪ�W��kO���Z���?'U
g �ſ��T6�y�+�L�Ч�P�)
?��n@�/J,��'��P�&8�G� 4V�X 'UOv���e�MQ�u�m�eSau��
�=�"�����Od+�]N�$מ����C�T~��X���Y�;oǘ�e\�t2j%mc�!��N�r����[��n��`�����7�`��+�O ��k4�9�@�96�"]�=x��~ޖW�(.RT{]]ۄ��^��䝥��X��}�jO�_^�wyn��$�pՎI�*������8�0N���w�2f\w�z��Kg� i�LZ�*��n��gȹc����Y��1X�5�"�$�Fs净
�L`\M�cb��Q�T��K�2D�\�Is78we[{舁[��S�֎����n[���^��J�z;9�G�	��D{J})������v����Dq�	#�vv~���n�0��?{cj��C�eed�Ft:փK��溜�'܊ܩo�Un^����a;=9L������ �͚�]E]�>���X(�]�u�7��Qҝ6��/��w�C�rs�l� �*�����oﰝ�ӆ�o���t��b����8=���bp��G=cSY����A�t�������w/�_��o�W_���"�+=Y��<ʧ̋��茷Щm�,*\˙͖�s�"j�m��+(e�r@nΨ4��wX��H���Э�7Mۛ�Ζ �eKz��n��t��AΰI8�Uv49���t>�_ɤ~j�z�ma
�u0����$�=�����~�W���Ic�5�#�lcd�{�64���StM�ig�t��~]׃tR6@��v2�x�q4�u��7�+L	�3�W��g\a���O��[]��[uK�,�"�:�^�{�^u�� �����hҹ'�й����������K��=?3�5Y���ȿ�W�v0���3hDYAM6z1� ��@J��s8=���ɵF�D<�	�P�
G{?��j\ef+;1m���¡�j�Ő�(��5Ҵ�%���A�.X|�h�=\[I��Y�x ��i�1O��Bpw#YG'�i���Vo���
�'Sn�/�Si!��Jx�)鮙��_�J\�4�{�G�0��+>��0��2��v�o����S�1�<x�b�w��	@É|�*���X�`��$���-���y�+.��Ğ���fn8��cC:Հi�T~E>4������S��CX��[^Ea]\���p�Vi�5��W�^F��K���../� >����|	���O}運p�Rֳ2t�P�YW	�7[�Fn��K D_!%��1�KѪ�g�\-_�ýߓ JkW��PϦqgd�<r�_p�ֲ����ϯ{_��_�#��t�|W!�������"�t�?��}�yv0��ב�1뻧[e�Se���Թ�P�X�bL(�)C��SO�	��*m�did�ـ���j��s�$?I�� �ͷ���Z^^B�M�����>�޵ͭ�l�����o�.�>�������Wc$��Cx�'�2}�w�u�؝�\_��k#nh�a��j�frҌa�"��
���ʃ��y�_۞��
���>����Iv}�����3�RZlT�c\9��Q����%3	��n��Xd���P�#/�.�Qm�7i�������(��s�o�f=jȫx�� �]�+#!�|'?��ͥx�����������ő	�����+_�]���7�E�x�2[��¸�[��s��ϗ����v��ٶ=t��OU?���~��������s�@iK(���*���/,,�kXOx���K�oTb��	��$x�>����D/������u��*�����+>/ZO�%����W�V��xrt�qy�4�u���\.��,�O\�C~��Tjo1`�N�좵��ۇO'=�u
:�@QD1������)JEfN��t�&ƽkw�c���+?�%ok�m��=4"\��T��GKQ�O�O�F���f���O�ӧu��H�k���3�֮��%�<�o�M���SʵT+(h�^<mOP�@W�������R�N�w��u�����H�\[Y�/�T�)��(C�����;{����pC�i���>m{��"��'~7bp�r;�����e�@��'u��7a4 g1
5��u?; T\�ή2�������52�:�ɢ1�V��g�3�:���r�Ww�m�+yJ���>j�+��/������lO�8?Ey�>r ��� �=�I�]]#k��;���꒰�vRG<=�¸=��؇N=v ��OAe0�t���9��笺E���\�$!�Y��\�ExwR�PB������Gҙi�.p8�Z������ݝ�����3O��HW�t�JX�P�Iӎ���e��w���xG�m_�ǁ[��ֳ:�S�ō����s$kss]y�>���;�'��0�d���5������r]�yo�d^��}`�� ʘ��(g�}��Hޥ���nms�'<[=��3��D%����ȃ&�t�ק-�Q��|����Î��X��n#��	���ꍬ����n p4�ԜJ�HV�H��C��2���K����^b3^?%�M<�=����2k�T�كa#TJ��SK*F&�(��S��BM���~$�兄�W��3��@���7���:#YG0�FV?���r�d���-��q��UeM���CgSů���¡�N��rl�s�G��XW�rR�c{Acd�'d�n% ��	����2��ח���	0�� Y���8!�0WzFTjd ���e�Ը����	���z�g����2T9ep�G��8��Fم����W�#�:b���n�R頦����P8XCc"%8~��QP��(�V����G�¥Z�UwW(�=]%���Z��������Mp�'t����
����{�L_Wn}zU>�'F6[C㥷�+S��7D�|܇���s���3L�R�J�{�_��'ޛ\�4	vΗ���w��g)����"L�Wҋ���o1�{�+���㴎ɩ������U@1�
��wg�ꑭ:�s��V�؀׆��w��܄G#�ڃg}(k4����r�͢�IҸh��;4t�(.�4�(�(M��͋O��+ �W��x�/�$p&��ą�5�:���o�����t��բ���j��C����ndW��6����jW������o0"��,G�\#�A�M���7^��1����&c�/GFz��@M�"���~5h`�S�4_ʈ��x�p�rf���M�YY�zE�كyё�#�y��x������1��n;><���ǎ� �t��J��Z*J^��T��ɵ\K�z��+y'D������w�+���먕��/��9FU���R���m[�c{�������yw=#[�G�jXM;J0S[J{��TS33ظ��1� <��^ �W���T�8���"~�m�� .9(��'���
������³?�B�|�ܶ��o���WӢ���N�<C�?;u�9���S�D�W��6W}�N<��*IN���iGg��x�>m]Ү��cLg$��Bڰ*a2�	����$�M�_\G��Ȋ �^I����Z��P��a{����m'����洸}�e#KC�Y�v^�����
aq�.�]���F�0���ŹY�'�.舖�~��|��&�im����gk9��uYl�B�w�;�?�ǩI��%xF�9��:p�@p��45?K9f���3ۑ�9�$��{�=����s�+Fx4�:��f�#���.�C`L!�cP|���޾��.0&&�=WjڰJ��T3fT�]�#�{%��i�� ���[u0:��O���_��߶�����A7�@KƮ�9>>C�;��qO����=�-�$��S��sڎ]����j?����~?�c�S�Iif<mg0�V�$Z�������mll��>Ű��4dk3� ���i�������ީ�G�Q�t�{NdM+,�髻V?l`,}l�z���i��G*C�'|�������(�����;�}�./(;�D�x�]t(`r�9�$.�H�\�����0���q7��$�d)�Wc*�p$	�F!�ĬY^$G¶��!^�m������֯�^�;Y	W����uiv���W�o+��!
z�����b���ȳ���uS���L��q����6Lm��]�wn���1�T�6������fw���{1�N���2�a"P�\SS�u�RU��	��)L����:������t�;���^�ש(�zvԣ�r/S`�G���<uܡw{
Y�h[[���F��.h�J4 R�2������j0�F�{���n�^F�J�����L5�<�0t���H0�*Ч��{�TX�O�Օ0�@���n�>!�x�@�4�7�('Y���+���#���M�|`5�i��L���,�Ճ?0���0����<�;��.�{!�^�#�\y�����(�P��N"P���e8~��V��ܢgZ�V�<��_�VO��b�",d{M\��o[�:�~=XzG�*Lq�!M�r�4�xT���p2؀k|SJ�
�� �}j�W��>�������^�^/}�km�oʝ���g�E���lH��L)���ըG��x��b��ݵ{W�'���8��&�t�'�l�]���{a�7㚢��ǹ�+��J9S���x}��8�(����zW^���<w߲�-�F�FOv<wD�]�0��վ�jM����B'��� �K�9�Yf��twur+l�Aqz�=Ҧ���J%�o`U=�#y�A�{����w=��Y�'h)���x��A9�H|�N��5�ߎ�lS��lŀ-bq�w2��VM<�s8���7�h���_��_}�5X�"�_��)��̲�F�:#��)K��|� &�$�O^�V�C�F��X�4��E��;l�|���?�ZrQI��Dɣ�r�9��
ib	�w��	{�L?D��;j�{�������0��E�n��0J^�FƜj��8*x�1����Ȣr��<K;ښ�"oI�h�r��%4qN~VǇ(_�mg�#���:H�����Q|~l��߶��-�[��� wg�w˻9J��8��[��Ev�s�#��>D)_|B�<����h�����[�	<�%N�&����}}+��.���{�����؅�"I|W޺�<4�����\�U[�v����L)�^�/1�x�;����K�C���/�W�������M�`b`]�(^�u�F�q�,�kӻ��aT���|�F����y[h�`G]ݢ����Y�_^���@[0(��߷���Ȣ��Ù33��+��Ϡ�~��W�/���t����)�:��~�u�v���nA3�G��ݨMe��c�ܵ��::�wJ�S/���_��Ht����Ծ�ٶ��.x��/~�����+.+x���m�C�Z�RO�ĻB֖��,(%Ovݑ�W���Nĳ�d�Q�(�ˋ!o0\< إ�d95K��2]�*�!���1�f�݈����Od��o����M{�l���_�� $@ۿ��?�e�M;I"�m�-��-���'���PA�`��ܴ�����{ -��?|�����������ߵ���߷ݽCj�8\G�I��2���U��9l?�������}�}���@��hhbܩ֎:���	<�������}��O���6F�A�w�a���I�yxx��|���ᇟ������Ǐ����d�I�o�#������]���Ay��h����������4�}[,�4�M��F������l�?~������W��(���q�)���md��V�_�J�_�a�p|� �X7�|��t����r�=w�_y�R'hf_IȋK� ڹ�����D�Q����4h��<��U�~x�=���˘��$�:��r$�-ܷ1>N�d�70T��t�T�wz��BIE��3��l+Ӟ�)isw��S�x^�(�&v8�|��kU�>B���vʙ���W�\[�btNS�d�X��q{�x��{�CVY'W1�O1�N�_�Ԧ7�J1h��T��V�Y�?odE9'��V���y��"
.��}!�}��j��iI� a#��H6�(�K#��j`]_�g`� =�,
��'J	ēE�x���p��ރgg'�s��4��Rg���T�M&���ְ��Y�!!X�ޞ��m'�Sr������N!�� ]�0�:�	4 ���7p2>▴Z�x�ε9]�Q9qf}W���"e�޺��H^Ĉ'p�7BA�	G�{}yY�$O&I�sUm��)�\�)�Y��)��UiV�X�u��EX���C{>��4�����k��s*�}Y����������O>~/�d*\�-���k����սoBo�Q��L�֣��E��zݡ|i�K�Ҩ�:��Nѳ!���Q�1�|��ʢz�g�1��uݚ,�#�K7�� �����H��N��P9�����e�
�=VG4:�{�mwg'���|)�}���/ފ.�ú�1����ڇ4x"�+S�Pf;��gM$�FIɉ���;�Fer=Gs��k���o��XNEQW��Q��!��х۸�(��|�`�U��2�N�S%54e1��_D-�7�<�q���v 仝:c��d�غsN#Y#+S�Q�$�9]�d�x��#���]E��:x��xtЎ0���^ӫ����v2-�gG�PRUj/Ϝ��p�l�r7ޭ�=XŖ��Ӄ�;: �;��l{;RP�޴��(D�D��{��{���o�:����z�p]\Sϥ�LA�U.Vςu��i[9�v�^}�.WY�ƀ�D�.�B�+L�p�>���TQ����<E>H���Fյ���דּ�"]��p|�sh@ڃ��?��i�wg<��Uu����,�{�S�>N�TkJL��%y��5ZjG(�8m��J��y��s�6w����vv5��>
�`��h Kɛ�{|�4��j x�����⽚�*�[(���4.�w�[h��
����:��^���m㮑�������Z%��@e�k�<����i��ͯ�[~�S�v���ί1v~���붶�71֎��|�,d�m��ѶJ=c˩�Xg�";��1 ܖ�N�q�r=�{���+��Nϟ�_��71�4-�S'��3�S�����z�nα�|\�q��i�>�|��CG�����r&�u�(���Q#�̬K��������Q�����3��{�=d!�\�E6b8�-�ܶ٩a�ӵ�����_<͌�n��Y���F{�v���f��Y��������O��H���;`���C���`��!�����?h�:�����~��^���^���}��}����C�a������M�6u4��_c�B�{mg�mm�c�l�Y�������޴����2ڮO��O��ۏ�߶��Q���?������Ѭ�cd��32���C���'`\oo�Q�7�}���{��������sF�5X�^*��B��>�S7�����A�f�(��1�#P>�Uڏ��%�䷤ghY��O�'����3?�ӎ�^}����$�i}��]�_����w��%:�$��4�Z����k��k������z�J�7��,��%�<��:�Ӈګ�����Y�z��Z� ��,���;c�M(#Y
C���"A��mxS
Zk�nC�S46Z��G�IO#K#�w���c�(r4��W�'���n����n8�#~�x9���g*� X`D��1����6��u;:�5Y���`Y���pXa�GJ14������UI힑������ȯ�*�FZݧ
�ݗAe%��� W++��+�V�0]w;j`�/Q�0��nϫE7���)!�;+�L���v�����@),����<N�rZ:r�He?�SU^TxTdd�"��E�z�t��t>��:7����$�4
���eR�jz�M�0��W��YП��Q�
(�cX��U�V�Rk��W&tQ���Fɞ�̃�pQ@L�/F&�4����G�������^k��/���e>�#�hS_�����$��M�L��Fz���`Z��`��K��_�"��F���*�|�+ta�
��8�W�뗤��b��!Ҥ�G���څ�ѫ��u�ᤁ��WQ
T����z{��3�i%5��Yx�H#@d#�PUH��eQ�x�;ﹱ�����	�=�;�;u~�1�#D�c���̹�l5�T-��K��+>��+�����؄
)y��|���l���>���C�C�Y��`�Q{�����7��!�N��ĵyq��k$�3�Tj�
�!��H����ڬ'�[�m�@���2Y�.:0Y���+#K�Qٶ���5���e=��q֑�溚1|zJc`y���t�!;oK^9e�-����m�]�!G�v�?�]�Y7��r�Kc��0��w0�Pf������@���jg�c����i�m�X�)ރ�70���������ow�6o%����Zw�s�Ý�q���^�&���]�t�C�k���Qh��4~tl�R{�xT�!��Z���j�*��;�œ������Ϲ^nH�%yG�r�9�;Zl�iߠ4�Q���F�W$��m�:y@5�R��_�d��H;����-?�-�An�W(�W��>vGq4إ۽q�صRRN�:=à���)+�Trc�`Y
lu��2vᡕ�'�Y�i;o��e���$��x~�S�Iq-/��
���]���p5�u���9 ��W92�C~�;�8�Xq-�|�`�SY�m�(M��X�4�����n �XG�NY��ğ�kKȴ��6�������(R8�ȍ<\gv�|�v(Sܚ�]W��5�ٰaX"��[���nݥOw��
���]��n��nh��f�Z�/���3Q�;G[�'�C}�O�,u���K�О>Y����}��ﭹ�?G���C���+Uo���X���G��>�~\��:u���o8а�>�o�B���W�|:Ű�@z�1��q~�Lp�1��)���!���:<�}���M������������یJ�~�.FW����Х7���G�{G�7�����m�����6��A�^;��>@��Ȁmڤ���a�y�lC�l�N2rJYΐ� :�a(mW;\����-�u���� mC�x�[o�mA6b��y�������C�L\_��]�s���2�ڮ�W���Oy����[e��q������%��u�~򲽵��$� >��W�"=�a�I{f����/nP�/=����=^]j�������7uq����/�*dY {��@��;�P��{��#:�8��թ=+[�;d�D1�0�L�)>���ʀ���C#b�#�����Km~:GǞ<z؞yq6�p�h�,w�>�^��G���5wE95��cd������E�GyN��v$+�Iős)���TD�R�T`*<꣔�ǜ#%a�M!o�gKE�[sp}u�5XY�$xuѭ�r�q.�HFlҫ���6`��i*)�<#���9�����JԞS���ڛM�ը �xQ;Cc�z�OWQt�8����a�qJB�X��-i�u&w���N��l�E�'�ۛ�hVz��+�S$�Rg
֌l��;�+=�5ʢͼ1��` T�e�����m�w*,=C���u<P.S��#� ��kn�g��W�p�:���̓�"(~�=ጰ1w�x����_>Apҗ.07����a�G��%W0��}w�'FG�A8�w����׼�_��'n�Q!�;J4�C�X��[���dʞ���p��r�*��bm��%��,�v�����ʡ�+_�_���hZ��2���#���"�V^9�"��7?�AB��NbhI��#y���(�)ϊIB�H����z����N�gT�E�he4�R�����))��O�x>�ey��7���~ݞ=�
~_��5�I�u��BY�Y5�F�%^�f�x$���u����s���	��*dv��-�:��I�rc����v��hc�������N�6K���tn��hVXz坝:cî#u�r�>2�i�gԕ��G�\��<;m?���^�{����������ם͍2��eTa\}��;�����zW��z��`s���v�7�]�x(��;[�;���1�mg��4.l/�25F�ak`pM/�������]K'�#�F��R�]����*����MEy_o{g2]�?�B�W���e�1iŴ�}i�@�A��aG��]�r>59gL��"�� &-�UZոwd����m���n���#��h`�};J"�C0r���s�N!�"Ci8�7�B=`��~�,�����(3���Y���-�A6��u�ڏ����0_G�=���EKss�ŋ�9�V�Gcf���Y����_>�7�X\X�q����[�Ⱥ���&d��٨��g\g5;G[:��R���.�p��3K�w��v]�U���q�Y��~��V��e�&梤�+e�ۋ;
�r�I�� rM�G��7��ߑB���z9�ʺ��#�]��ܐ+���C�uݭz�����&F�������W/��2��R9G���:h?����v���z�~��n����O]!˷�b�^���㶟��Kt`ې�mn��(#D�߾Ɉ܇�b1���?�H�@�;�E�𷻋ᳵ#�i�����k=�/�����)zW�@��Q�{B���>�N�C�;uU`C���K[ogԹg�jdit}�=z��}�#nb���ճm]�c��	u�+Q��g�hI��H�&rNz�$�d�����������Q��+lo��<%��ī��x�z����a���O��D���D}I�r}�8BU�ܗ��M��-���m��0���j���h�v֙^�$�Y��m-N�)�C~T�L��P�M��+����K��GK�m�3Z���F+��H��;V#V�� �jML�x�)��rb�Q�c�C� �'N��a�5RT��G���
G(��i0�2��@����HT���Q��X��s�*���E>8��ɑ����
¼j������.x$��[h��(0]�v�[(/DK@U	��p~�u��0�cd(�@	򝢽<�<��]Cp��\/Ov�Ⱥ�I�7W?� �9{��"E��Bjdd�z�7�ΤC�*�=#�Ӝ:���mee1���N�
��+V	��el���/�Yh��\��T%���o�=��0�&��JrmL��+1;��Ц����aA�{~Ȣ�o̹#�dz�����C�u�oX����_h�2�5xv��81��k�ƿS��ȝ������r2���׼����{��W?�[ǆ�K pk�A�r��^x�q$��YI�9`��!!�\�V��d����.�<��Õ�|z&ӽ�i��4:����(�y���4���ϡ���DGm�xC����[�C�C)'(".2vj�FF��b��P�Hkgd�I����w2��j=S�#-H�l��:U{��(��R����1[_w����2�,�p�ue�����'E+�E�O��'`�%Y��=g��]B^��)e=.���O�-�uc��Jev�lS?SsS����oݾ�/�>FQG1'���M���_��k`9b�ˑ(��Q9I0r3�+��^�~	U����8��U���q����r8
�(�k��#G{�Q$Ļ��=��i�S(�v��^ĸU�)cP�=O��.r��ӎ �u.$5Bv�N�Υ# 0~��hd9ekE��.��[����v��H;�H�p;ܦ=�C���_YNT`\g&�ӑg821=�Q{��{P�Δ8��N�^}����J���L��Yh���yv�gMˣ�J	�ff=I�_Gy��-���������+\��y\=M�9��[1�����M����~#�h�#K��F��(�4��3.�ى@��8#MI^�����E����:Dѽ@�"�b�k�W��NE��8v��F��7*��S�#�(O{F���)���s=�y:�������������
u���__�˜���l�62e�4�Ww�#��}�(�oP���#����ڃ������ۇ��w�����o~�����_����e@^l�ӵ�D��]#�v3�d�ce�2�ܭ)�:��IH�rkX߾s�܏���>(�Ewpq��u�u���ӨW�{��x>�c�y9���~��q���ڻw��'�,GS�?"���qQ#��%/ֿ�$3&]b��B6�Z#�<�,IrE9G�E[Z��f!ϟ>�L��Vw�����^�������q�M�w�r}O#[�2j�"��~����K�о��1wN�;=sGj�O��7D�<��v��	�����Ԩ��1�=�(�[Ϯ�^qב[��-�a����b�A�Tmu�Mu���`��[�����ݽ=�tg�9�b�;�[� :��@#Q��uV�!Y�/���`cL�5��fm���
�I;����*��.��Q�:V��z��sYR�����k.ƭgݽ(���_{o��H\}<���gm�	neR��(���x��h/�7Ku�N�>Mi���峸P~9���.�>\k/?l�n|��bd�������}�b7w�&���Bq�]K<
 *�j{�Q�a$�,j�⊆ОB�Kj�2d�e8�� >����4����aK|v�b����{���0�潖%
�J�==���m����U{��r�Å�䑎�l|�� ���E�,h���3�,ޝ�@���Ɨĸ��Py__$C٭5.��;~��	HI*���G�J5<Be*ȃ�(V#�!�Q��C�!�ꫳ��<��Z �ߢ�8����im�����=�7�J���w�Þ_�U��=�w��Ch/a�,O��U����l��c�\R.��u
r������'/�nG�=Y;�p�ri�N��Y��gO�u%�F�*�]=}�-�(�Ј,��.M��ř�6�FԱF�uMn�E��ܥt�t�Q��h�yҖ����ѭ�����{`A�<�E�z��k L�k�B�s��L����!�:k��]O�I��D�Ȥ*�)�7��0��]�P��OZ����r�[]w�)�����˵�Jd���_����%��׆&~�5����fZU��(^&֥ۥ_ӕĉJ�x�*&5]Ե��`�}�V|ؠ���1988@	@�� ���	����V�����{A!�tS %�t��-(|U��kz�s_<D���S�	rÓ��QH>}��do����ܢ�У4��u�����7}���ʃh�xW��H�!�֐�)|�1�������4��4ys��Q5�'��5��d�_�W_���|�����9��kd��S��Ho��7N�u]��t��7G뼣��o}w�-�*x΂a��'×���U�hQ\J��
T�N\R>��Q4�%کK('�`�F��??f�|F��rnt���&iT�7ծ��[䒲<x��N7d��1�R~��seT����|zze��5z;���Ȟ~{�]L�w��-iޚ8ŉ1��K٩[(���	����#jL�H���U�h�H��rH���w�{��4(;�M��oנZ��9<�zj;I��B�R���\S�:$x��ۨ�
�����v�2������Д{t��F�{���i��ܐ%>�4.�bwFZ��}����S
vq3��h��m�-�7ۇ�H��X^Sw��#�����I���r���(J��ǌ�^ߺ�;����@�(�@xyW<)��Ip�ќ��.�;�����1F������;ƽs���(�gЫ�S3��E=���GG;m�`��̎��Hϝ�.���?���`�o�ɱ���ѓ��ɋ675�<��sM��hck��bdOalOMyp�<�e����e�u�D*7-������1:�o��w���Oms�S[��8
77؇�1��{�-�e��#�ӓs�{y����P�YO�I\�əm����h���}��B92~}�A���w�ƍ�3�-~�Q�1p6>�F'���I��_�IH��0���;���d��҂S)�7z�z�9��ÿo7�ڛ��m��S��(4 �\BWY�(��m�l�&'��2��h4�c\]�k*�%�|N�b,A�����D�%N̒�;�N��/^�7�R6߾� U�55�N���rJ�����3e7��f��r�[v�D6�A��0�	ϟ��#C�j^�t�_�p<�S�� ���#9rsx|�66>�ׯ��ڎƝ�4d��Cz���lc��Kv^�6%尚��~ur��=��o�*/Iĸ���>�	����
U�ſr��۞��"��)�\}�}�/�u�� ~7���v�a�0����ݶ��1�td-��-�k��@��A��XYZ�,�+`�Ȓ�����	�w���)E�Q�>+��P9ҥ1�rj}�
�&A���&M��W�HS%���F��	��������b.o��+�p�gQR]�*Q�o�.l�u��}�k|��������jb���Θw�����@��e�B���Oi���r���	e}
����<(Wm� �*)��PYJO����=񚆤v��i�NEXʢ��:5B���!���)���Q4
��/36�ЃĬ�0��A���n�ۮg��f/��v�FVv}�]� ,g��(��5��E�477���\|�_p��i�go������+�ơC��Qq�(�aQ������&=��>=G���e����e3���̧�P��sw_�B�L�(���A|n��W|O� U��a�Ĺ懶������(>����pa�1�յ���i�q��3(K��u���p'S�����'ߠ�2�I}Z�K��w�'��������*����}�J�2+��lq����Q	������O;�oLCy��{��E3\z���?�*h��F���2����ԉ� ���F�x�`AI�e��������gչ#���C�&Foc��+�&0��s>~Q�r_��Y��u�q��
��B�lN��tf��)r�Er$��5�(�ݎ��Ֆ�m�}J;�;j?��s~�w������Z�TSe�Q��Eba�SkJi�xN<#�{��D���5�ҫ�q�p� N�-�1�[�TW�)����:��W{�3+@:�#���E��IӲ��$�Z�Ѡ
m�]_wX�cg*�����L�օ?����+��%>��Ӌ�L�r
������^��Ő�����9�(pFxI�.�@8���Hn��n2�C�]#���9|�>���KiU���*�}��6�6�i����d��?uG2n[b\�X���IG�KO[{��?��}�������i�޽�TA�u�_uR���S�bPa�x���J����������^����q�6��2������������������5��Qbא�k�Q�e�d�y$N�x2�v�y�˹Z�������z��R&uDqU8�[�	�I/
�D��&B���B<�S���d~��������l���,;����|IL��.w���#b��L��F��5��K���3r��%G���W���@չT�6����qG�y��uz�S/��~YE��P�eipg��YFy3c#��)��z�K7�,.�Q�}������H��l���0��������{�����	�q�`M}U�!?�e�l����䙼i���=׻����i�����,���w�����+��k[�>M婞�C[�7O}_���	m#	Jl1���~��"�n�q��Sټ�p#M��'�v�g�`�;mT	�)E\:q�"+�J��ՐU#�B���4�F�	5�
��(�gC �T/�0Ј�MHT���:-H�X� �������I�������2�|�Wl�bP�~���{�T���;#?�'�J/�S�#�S^�Z��c`� �������	�8�ZX�N�4-���w�ȘN����k0�8 l�#(2��nێ�^Zi�˫mia�l����؋}{��o/M��"fr��п��k(���@��������{���l����mo�S���:��i'�K�6D�<Tx[}'~lLz*��M�)�Ň�̔�%�`xIo�@7^���|��!�$����s�͝�\�Q
�#{55�h��,�Oc�CN1��|$�4�G�Sh{�}��U�݋��]�I����u��B���}�@O��|��d���[R�k�ß�	Ӆ�cG���u�g_��M䁲C:��=����iiP���?�+z.W���4�I	�Sݦ��2}od颼�xtr���U:��*��՗#�/���F��e�h���9YX�gOe�V��x��=���;5�L+ûQ�J�#\��6���sm�������<P�����|��|�{�R�����|qU��J�\w�#g���Ty
��dZ�F����P ču|�5��~�pթ�g"C�cC��*WK�ꌬ1��q�5ӛJ�ovN` i0i詼T矊[M��s�>�xԣӘ�+N�2�>ky�#�
������sG����z�m���⛷ƨ=ҝA�ס��s�k���t��r}�gx�:��y� S��{�7�N9��Qd�����l�ik���ў_�6Z����GAӑ���t��A��"o?���jȻ�E��ȥĕ�Y��5sbǅJp.�TZ�ب���nt�M:\����꼉����o߶���w�>}�L���0ч:��T݂7��QLG�0����������,^�G�5x>|��y?���U>U���A�y��<��,�
��
�S���t�֣���O�YXO�vp*��_\�sy@�ǎ��q��͚�V:����i��@+��F��Ƕ�9mYY��j��'�^��7��h4+,���G�҄�+�t#�p�,s$X���oЫ��A�av�����PQ�r�q�8�NcV����dgIE�0�`�x��v»|�LӧS1�_O��UU���d�B��}O���S �yթ�?�ko~������u�gw_�Ŋ��]�l���S���
V雷��{g��o\�)W�(#�V�}��dnᥓk){PC&p�FT�c\QW�����G\V��z�$�!���Cp2�-4~>A\�6�q�:���I��TVӾ���E����8�-�P]@?�c&�v�s�Eڣg�g��BGp��4�X�
*�&.B�ѩ��bl({j��k�H�;�c����C���]���{�w
	b���A�ҹ���.a���kY�Ǯ����!0�J9){F��"�L�\/.�к��G�ψs���	�`]�䞡��pѩBb|b:S��ZYZm�+k��ʃ����9��	`�șub#&Cnx�Yf���k=BRC�!TG��'��`o;k�\Ӏ�u���ǻ����x'�E�P�\#��QN}����G��!`w��p��6=qK�7�Q5��'���t�;�}yi�-�η�Z;�s��U�P��Z�lީ�]cH�\��5�(����SZw�sa���8/���q,W�������ť���d���,�|�C�.��w����_��o|��
0p��[��w]�8�������=����<~�pVh�VK�V�]Yy(��W�r�/�sJ�;1�(�+[
D)Nw=�w��������Ѽ	Z ��	��R|���c���VK��&-��2yFC�:ҽ�S�.d&/+%	ͅ4�Y����OC��]Xh������J3�ahh)+���z�;��=n��w?������_�)G���Ɍ~�#���X�`|idU�����aqp��[<P*�ʇ������=���f���u3VA)Ym�l�T��2X��C%W��M,j��rY�*7�Vƕ�b�E�OҊ�g:���%�����0��Y�K���ˮW�A2U��V�(����3���^q	L�!����D�����&�q��B���L|޶���������D�� 5�)~��u'֧�U�X��%K��Ć���)���@F����еt�myy9�T��Mh�s��i��l��\(��:�<�G�A�a�k��~{wg7��u��?J�lԁ�u-J�k�OpH�.�,�����!��I��I�~�뉎b�8J&�h���g��Lg���@u.2���R����"�K/��Ұ)���[��ط�)o�~S�h�z�ii@��4�T>��;��wPh幢a(|8R��峺� �`x��Q�{Œ�0:��c0�u9u(��ݠc�xX��u�Zi��g:������t��BN�*����w�{d�,��SN��6�y�r���s�
���W����-Y]8��M�g��+}'�%Lћ��'�
9i�\�3Ӵ�Y�H}̓�7�ߵwo_���޴��p��j�=D����X�zw��y�7��������}�p%O�=��7�2���M�\�w1���Ai�G`�p!B���+��;"�N��Vu��K�G<�\q����0߆41��PE��8�1��;�d�i�>�g�)��Lrp���s�����Ql@�Wĳ ꙙ��XH	���J(acd�Ŏ�zN�Q�q+Қ����9G��$�kj)F�I!*M^Ǜ^����I��O�X
�r?eIz�W<������Y���K�g$�W�.Ěk�R�q*0�?0�\��{F˅Z�/�I?'|�s0� ^�<P��J�;��$D8���<��L���|[\~�VQ��y�3F��F�r�����5�!�j�b֦#Ë���>S;Ơ«�5:��gG�<�p�������^�a�nO�y4
L7��W�����7W���R���s��j�c�3�у����Z{��Q{��a{@ø03�f3u��M{FҦG�x�
�sw���G��J!���2w����A�ۥx誔9_��{P$���_�pw����%�g��(�\�np���=�.��G�/�Px��T�g/�;��p=hgZ��4�� TP���ZSYh<�i>�����c����%����fe�
����� y��p�=h�oUA6�%�L�*�*ؽ'}a��Ι}od�	�w��ip�JT9*�����̯?�j'(N��٠�wWז�i�Y����S�u
𜇃b`�|����q�~2�hco�J��; �����>�����8�.��Sc��"E��(\�F�`�8eЩ��+�����rS��}�X�P���v���&f'vF���uSƎZN�V6�)�1�@I���vSxީ�5�o�ԵKv�������q͑r;��){�!�z�+#q�_kR�y�qu���4��g�D{��F�֊�X��e�c�L+E�uU����9�X�H`��&L~5��0��5Ů]9��iGmg�4k��0�����m�G�M��K!��1���H�uP#�ƫ��|��k��2������� Y\Z�q����{�k���8=K��mW�x��Lz���.�o�9�^�SGUk�W_�ʆll�)���<W��7���hL(�ɛ��~�[�y$^4=�ڭ���'h���04?�'�Rʴ���úT�����Yy���4�K����ö���F5v�����Z���0r�����Ex�������
�� �.x��<�P���6;;�N��r�;:,�#�����x/Cγ�j��c�rɂ��4SF�4���؁C�s�"-e�f��D���S���� 9'�<����f�AY�����AN�t����v|�����l���6�Y�epgeQ;��2��P�Y���Zo�Ѹ���%�\����O�m���P���e]�I�׉kӐ>J����o'x��޸���샒ׄI�^�`��ύi!׍��9�wֱta��O/�G�Wf,^j�R?�Hw��S����芎A5��"�(�c���xB'��G��c��,��j��8t=P�b=��w�����/BTw~pAb�<�J�[G��룓�����`E��j��ғ�1F6�~�B�S�v�t��[��ޞ��(�Q���*5P��s�o8��2֕��[JU�V��7Za[đt�K|���߻���Qu�׻��!���F߲A�#���o�O���h`A���C �"{��t�1�1��f��T�RV&ڔSh(��匱�"��@�e���Top�bL�gf���֡
J�g8-J�ԫ
�umo�om@Tll�ςW�pt�p�>�0iT� T�g�k����v��؇�B{������:oc�mfj(#Yk�s�ų���7�ۯ�u��/�i�����W/��j��8�G�([*wk��N%��'�!�u�>�����[�
=���$P	���ep����Љ�E)�Q��O:i����'�S�^�wE��P\�\���ߠN��_r]N���:@�s��W��	�"O���{�Ëţ����t.��ӈHoq
e��~�'u�EJ^����HS����(h��T>=z�]����pM��F�)�N�Q���"_��/K�UF����w�劰P�ꍃV�V�Y]F���onF�l�����Y�'.��G	�|�q�t�l����,F�b�@O4�T&�7����Q�"���C ?犃;���Z����a���\� �o���!=6�F�Gv�N��Q=� ���p ��p\�B�Jܪ�h+���� S�+���]���X����������7���F_��z��{GJ f��4�2m�Q�Nѯ��.���ҘS��Q�N0�bdi/����r5^ᬓ5�*��/k�0�]DYu�/��~��I�Ǻ�N�(�I�Mq��%�TY��d��kǧݙXۧ�I���eT��	��
�r�����HGvrt4�]u������4���&Sc��z�Y�t$Z���RZ��רAhC0��'�>#*�c:k���(=iD�I�:�ݑrT7gGx2

��I���]�R�x3��&�ה�#�i�f2e8�Ë��:��)�G��UN
F��ʩ�F�,��-wV�+�����tϩ�s��Ϟ?kO�>�,5y�ٵv��%�w��vj�����tg�8��'Ntˎ
G{T����ų���~�� �a��K�����&{�K��)�ch���,�ӫc�V���@�k�e�C¦��qd)Fun�6k�ԭ�-�*2������eˮ��݂����B�V����^(�rBy��g�߰N{���a��W7���;�{κ:�V:u}����v
9`aY5\���|{L���ǜ��!�̌f�y�/p��:,���o�e[��S�8BK>�Q��$�{=�{ɲ�7P8y�C����yx\v��d�V��R�L��Y����_=gݜ�L'�"G��tO�y�Q*bܑ�q�u��(e�N���� �	 �n��%���N��/� ,�r~�/�;[F�=~ګ��b�f�V�**7L� E�7�#I�qc��[v;���=��'�	�Z�����n�.�[D�������`�k���&Lʅ�
}W%�p�',%ї �G��U���{��k~	#��$��+Tl�k��g�+����R���!p�-Ƴ�E�)����q��e,8���m�����\[^]l֖���Kx�0$aܮV��������L9p~u�C��+V=Y
��γx��%�KXe��}�;N�%�-S�\x��[+{����r�͞��m�l�ӣ�vyv�����lӓ�mia�=~��^>_k�~�#�E���~���/�i��A�jϞ>n+ˋm���U=�Na F�,=5�:q��
#�Ѵ2������)�m�T������-_�����9頯ҿ�=��ݤ�������}@��ʳ�σ�GN��YWٗ�>i��R\���'�����o8�ˍu�4ϙ6M���p���s	��ͼ�N�?a�<��j8ٛ��&бa�����'��j�i���^�������:�^��ٛ]�~'C�O�+���n%�k�Nث�t^G��:p"��G��:��nVg�x|~������%|y���h���H�R�P^G�������5Y� @��PI��ɳFD�^\
�������=^{�?���Ia�uo����s�x�m�ʣ��'cN����5��#�YeB����wݼ�s����c�d?�P[��R�
�un��=�@��B��*#V���{��%�$��������L�3�*]C K��d��
����>�X�*�n�`���"���|�"y�Ɍ��l����z�Q��� ɫ�{���2�r\�[�ӑ;c�k�H���*�'!�i�2�<d�����"�qq{�Q� �W�(��vD�R�.�)�������\�9�u0�&r��*��Q&���VڲC�F�9�@T�H��]�2�F��v?]�'TJ�S�%� �줱ӫm�G׸q������l�蔰�(yUo OԺ5�q˘���\���u�
���} ���</�ꤱ�a9�!��۰1�������2q7Κ�s�o���:Uy9ƈ���Go�ф�� o��S���$�Ө�)�v�O��Ƅ����|{��e���o�ɇp�4�M!"��8�uli3x+��4ǚ%��p��>k0�<|B�,����Y.v� ���`���׵��%4�;����0��]fT}�4�[��A">�B|��G� �������F>�H'z���|FQ^u��ѡxҸ���o��Y<V��hLÀ���x6���/1��E-��_8*Sx�u�b��r�$i�`��>Gg���#�0`�=u\ᄭ��]��6yG��˯��2T�:��]^���(?���y"sMG�q���݃kUiB���K[��]�2��75�4�lM{�ܺ�~8@
�W�(���"��j:�{�;#��m��;���  +���2|됻��~*�B��4��?־����_����_����_����׿j�|����ں}ѡ��)�S&*�*I'�=���o�T�*�e�oy'�J���|�=�����_���Ľ���:�I<�y	�LG��e��C�[5]M�.2��ׄF��,�,&�jhu�T�h��(XW��1��W�r�gb���n�:Q�4�!*&>�w�lK{X�[�:(�\Ԛ).�s�����вQf`vjH��es����C��{33�=#g���`?;�0�sjrF����V;�T�����7�g��0;�,ϵGk�����B{�b�}�����_>o�}�z��a[]q����g����4�J�^����>..��.��V���������������q����������O^:������ +��??մ��_Ζ��u��zuw�ݽ�垞'>ˏ��7��D���8�P�*߾��^�I�Ӎ����4����(S>x&Z�U�{eg�!o�Qf���ީ'�b={�,#��*$��l���14H71���4���w��>� i��o'������)��^vC���G�kڠk��Y;�7�j��~�'�Yc(kS4������@1��t�}��|T	䋾4w�w��~�?���m�>[R�ow���RN��Q�&�w�%�.+��U������pR�A%Љ���*�Ż|7[R+�
�H�F���6^���_�7�������XO�I_xx/���o�:�K=ߍbeJr����֒��^g�I��P�B��/0�ԃ�hI
��/<ë��__�����l�È�d�aFW��	�#]�0F04m�5���E��o7S�e�v^���Ҩ4�I�X^;�4��I���ws��P�HF�//MH����I[��-�('B��K�W�8�������oǐ-��V������w������a]u\<��
�H|��0�[����1nR�ipU���q�����Wq-٦K�I���=�~h�b����+����Y��E��Ōn�۟#h�˔/��h��6�F��wP`�S�����ٖ�{7�Y�w����NL���ԅKV�!�k��mƀ�ח%� T��k�QN:ʄ��%���!v���eCu�h���5b�S����/��0��1GڞuX�=M[܉�·Uǳ�)/4C����E��4g����2<�)4 ݬ%[�m��hɇ{
4�;5nŻs"<�=���3t�5��Jd�-i)�S������r�Va/��t�s���<�L姺�Y�.��Q?g�W�,`�Yo�ˈU�C��򼦈���~������5� ��h��4AG��%��˨"u^�#��Q�T?���
_w���$P�V�q���N� 0i�,��m�B�2��x<��믿n���o�?�������?�'�����O�?�'����_���_���z��$[���d\�E��pK�\*�������T��@����"��%��'�φ�#�dY���C�����a�Eʤ0R�(���H�۫_^�-���qՀ�[�m+V�V�+m��2�C=�E����3*�!j��<���tA�QPlpj
�=���BA���,}Ξ��9�c�)?�	�����!S��)wC��*�������ڡCko�[[�;U�wN/tN��D�,�#3��s�man��͌`@���8��̶�O�0���Oc�=lk�Zx\�o3������������g��8K���N��&M���3����ۿ�K�V��P�ū_\{�0�݅ϻ���r��]<Ӭ�?�VW�/�Y;��I��s��� ֍�}v�,׼8��h*#
v�d�y����c=��Ro$�X+���C$� 2�s���ݞ@dSzֳ���Z�,��&�{�.�/�걻���(E�����/�#����U�)s�(�n�|C���ӭ�~#L������9g�f�7�lDn���Y.�Q�����\�8�/����Ͻ��Q�a W��P�E�J"iȍ@0�	V#H<���
O�M��'���[%y(�IS�N�A	Air:��S�O�E��E����{��:�<��'#�\�˚6�G��|{ެrt�+me�ie��:ʏ<�9=�^�tK\�u(>҆A@��g�[> &�W9w<-J��ˑ�<Wg���������e�����Z�7n�=~GC���(�4�u>Գ�֧
��bhd�6F~+`$.�T�ߪ���tԄnH]��z���TL&� mعS�T�<�}^ߕW:
�w�~�9t@{�6^%~僧�ն+הe�qZ?Vg�O�l�,,y(��.��®�0I*x�]�:��e���i5��{i��j̖�(��������!2v���[r�W�4u�	FI��оf��|�Q"�O��ѨӞՈ�����暮���x�q9��΋���dwձ8�c�D�qf�#;zG�2M�H���b(��$G�2"Uy?�ic�?�{�R�dZuw�q?A��z��~�������+�*�
ѧ����O�s���ʪ�T�f4����j�R�6��z����x���u�ͷw�-؋'m+mck���8�g'V��=O��uC2�+�)v|���Ww~u֜yD���bd݇3 �׺���9}��_��}���?��2�>1��i��C��\���/��F%}z�2���#N��ާr�aez�L�2���
Rhz��*%�FF�Ua#� ���1������m�����k���韷��������}��ad��_�U��������ګ�/ۓǏQ�Qҩ @��Q*!V0�m�CѤ�����s�r�) �����|�\^����#�T��ҹ|3�i�w�
��"P�/�eOj�c$ �	aN��)JN%��
0�O@X��?�!��Ҹ��A{�h�=����L���%f�Go���}'qkh���u�:�޸�xvJ������e8�1�����dqr��C�L��Qb�:Ck�-g]7��9���'G����j�h�d�sm���O<U�BY���f���&'����(�2�Q����|,-���C=m��]u�GM����Y��w߫.̣�#�b��׍?]��m����y��>w��^��n��>�pϯ�?=/�p}q��{���Ջ���������g�.$!"{�R���s|�p��})�������a*#�
�O����ȫl�̆[���*N/(��b�PuՔ]�/r�gv}���r!k+8%wA��^h�0��2�5pI��&�.����ӫvtt��l�ܻ���pW��0<A���7�(|�h����u�E1:�}���؉�����������.��TT�#~��<��}��y�Ng:�-R��*(*'^UX&t��4m�k&�W�,:?A)sZ�%r������;�T�YE5�˩G���2W������wi�e�y�	�m��J[��L�@�k	��@�!$��|;paA�`�MUu����{����{߈�)L��$�7N\w�1��cŅ�I'2���i k8g����:�2x1��w�H��Dj�������ס3��ed�\֫㍄d��Z���������ƤT]��y�) 鱓�y��W��e����}��7�������l��n�����V��<ehiǷ�Hܲz���=���b(t.���}9�%od��g�Ւ�KrA%Q4�{9�3~*_yX���6T>�W�fTHt�iV8�w��#'�VD%�\!�ϼI�^��� ���yX�IdXmX\�JZ�',{-V&MX?x��Q���\�o��lUI�q	�3���\�;�@<Ͻuϸ���?�Y��"6Rj`���Y�b��0+~ڍ%���r:LC�{a~>��4��,p���	��nln��Wg���ѡ�~
4���֔W������EN�U:�DuQ?�d��H9I���u�;qu�H����V�9tB��*h0�8R��i<7M֡r�����34��e�%�"��$=�������UN�GO둗�X�P6(��t}	�	m��"����|�㣞�_�Ym���!�5�O�Au��q���LЖ7���Lժ���湄��p�c�j�z��Pxי5/��r�X���#/#s�gu+��:U�?�����!�i�ުi�g* ��v«�Yy�1|s�a@�P&a�t��L4�\�{!D�WoW��u��IV&���8׾!�"�A�*��s�t{��I���M���h����ߵ��������q��_>k?�����ŝv��b���Θ�X�@�b�d�G\��'��@J��ɭ=)����\Na>����0���9���
�BB:2¢~_�H�8@`�z�/�Vp�݇�p��'0�`~�odf�S�\���!o�y@�G���;2����%h�T{�l+�s0&ad���UV#�59�ffڃw���<h?~�߹���0��f�"MQ]���n�Jlvf���ۈ��G��}4��w�ړvp�q��>���(�C`|��(�����0N����RV��F��*L7��2�@9����|ň�e;%=ǟ;�;+q�TqNw��99����>�*���ri�*<.N��A��>k�����s����6�㥢p���i���C�]R��]�~���V�C���+���A{9Xx@E���a�E��eg;ა�� ء�.�Wǐ��@;�~��o;qխ�6x/%�GC�Ar���u(ĉg�K��BS�Þ�ZX����;^ q(@Iy0�yg��X���u5�Ռ��@�B1/��A��|Ю��&<���E��.��
X�'��5^u���
�E]�tfX�	���iIJ�UH5jO-���gYu�]0�
޷�h� �}g%)��B),�<���{���8�g��:P��!cs�����j��)�?��^���2M�`�����bcKm®aM�����vzL����j�\���ӡ�up�6����=��O���s�����C%P%����<��)tq�r ��PD)�
]��@����:��RBH�k�J�[B���:�Ӈ��(���9
�]g���
�yg�Q�!N�a���	���0�T��uwoil��U������3���q�x61Z{����G�O>o����=��7��g��=��o�G�������΃_���?k�����mx�ĵ ��O�	�$���u8�9�3!?�M���� V�Ԅa`�|�1b��s7o��i�{�������{A $h�y�w]���	�&^�A�_z���9|��BR� �T���$@#<A[��(��&K���"�{j����|�������v崽~�>쌴���v��=NW{�ZuN�)?[�!�$u��5��r\�Sy�B��#��=@�c�YҰ�ظ��3Ϩ�o�T�]8��t��5�	�b]A.{�}��%8�ƸB��gXD#]+����M��}2��ck�'vp&	{;mg�:�%�u�Y�"��R��\���I;>�O�����`$��� �&����b�[��)x؜����i�8I}�@{�t�O���)w�N �3h	��P�rT���<F�"�yMͣKgy��Y>>m;����}��6'��a`0�p�N'isNL��̷���!� �R�q� ���y�?>l�G8�Gf�+�H�)>�;��5ȩ��Ӷ����^#`ңN������6<���<p��8_md��\u��w���,�ƁǶJ#7��W�K @��
�3'@�c�e�q{�����\����?u��������0��i����M��E�E�ـ�����z���ԁ�ҙWǪ?k~N݈�SCn�O�c��I����(;��?��zNy
C�<?�j{��@z]�q�����KK�Y`�լ�߽��{�՟��@ݻ��#���wnݚáZj��n��k��x�~�����}�>}�=y�wwﴻ˷���tW��'���U�2=���!d-�4���� ��s(m�x�G�����4��[=�?����z~~D�؁�%$M��_a�hΔ;�Adr���+@���`.a�M�ˈ�(-
p3�I�e-�iD� 'qb8���"^�g�������g����ǀQ�8����S�mkh��mQ����W�2�+�8:�Ʋ����!����zW%��]���#�H���tG��������
z	 �Qݞ*"�G���24� �ʪ絰�AŁ����\[z�z��z���v��r[�>00�^b���fk�ҏݟ:��I��i�o��0?���Ӵ���I��d
��$�l�kb	�SB[�\aʮ����V`�f����Y��ҩQ�h����A�����x�|Ւ�.�z P���`��ā�u����o7�T�JKh9�
2+��_�2
,K��L�o
?��=�G�ZI��u�!����<*��TC 9!��g�#=;��?�/J�bt�շֱh*��u�]>]�s�Ի;��e���/ׇ���G�#��.!ϸRHڳ�0�=��E1h`Vk'8��Q*1 Ho	���&��T�|�aKp9���`K���;;�mss��b���[ yˣZ��.r/2��Oeg�eγ\׻���Ơ�~�7�A;>�p�1�I�8(���5�x�@�M�ǹ��tP�:e�*_���q���䟕Ԓ��DKv�q�i�"o���:���.z��i�w��=z��T��f~���Ok�_pT��
w�a}�1�[�M�Y��5�N�ŧ
����z�#�;Ġ��P���[�ޣ�8Q���~����_�U��/����/����7�������~�7���_��?��~��ɋ�ڝ��م[m|j.KW:���U!�Ч2�X�o�6V_\SI��D����VB������^���!���{��!��/�w��������G����rd �} ^9q�Z�h�t�a�H��8^�81�}h��D`�-�c���8Y<#��G�1QwH�BV�U^�;� `&�Ua�	MY��,#I��qJ����e5��ty���tjbl/g扒Oɡ�r$�9(����â���>��H��R�G�PA�j�EƂP�ؖC�R-�XDF����=B�k��V3y����"�"��fB�A꺞��R��w�w�o�t���&�N,��b���3�H�f*T"C�gKfd����I���ʓ8���ԟ����|�.���6H+�Q[8�BZ�J���T��%��t8���;Maҕ�q���s�S��<�Y:%A�v�rV�]�r���7�}�s��^�qn��
��=�@>VG�`�����4�O��av�^��e��_�(r���1j�8�F�B�$�q3߽:[���vf����,�-��Gz)������9�G�'z���] 'ԑg~ם#�	EOۃeϕ[8�� <x��>�t������h��i�=z�u����������/>ν�Qݻ{/s��w�>�>}��J19�cx��LC
��̠G�����g7C��8u�3��GG��<1��4"�����:�$f��J��W�}�`M8Հ����{*ˡ�$��C�>|��Q{��y�;5%��Q&�(ȋvx`�f�(FE�`,W˦0(	�.�X�}��c�U��zTu�yX���������$��ȗ�����2$K���dUa.�c��"l���od�0��>��k��C��������<����햋=�TLO���FY��L��-������jY-e
'kvJ]Ύ+ZIƠ��o�p�3���T��S
ɖ!r �\�'Zl:%`���JG*ΉI'�S�)�p)gp��U�f�����i�<<�"n�h���&���-����v�J����v��\-��ete��d��W�4x&�0E�ǉ�%��/b'x�x�F��t��u��iՐx~ӥRѺ�@i�n�m�tpI ���e�S&�ٳ%4ND4�V(Bz��`Yg���J;�仟8x�g��ι'r��)����]�yh�R�F��4�Nw�;�K��AW9"j,�����ՊX�L5D�Bpqch�������ssj����9��1��H۝��7�c�����e��$�b4x=h��4��Å����&�T�h��( �E!���z^bĜ�5����D��CG���UƀW1��?9V���H(��pb�YGҔ>���V:������0�?)e��.�=C��e�I��ǣ��+ZjU5UdØ ��)gЄ�Сv��3�쉲�kʕl����h�?�Y����>��oڧ��M��g�^|�������g~֞����\?���ON�_�O������I�y{���v���v��Ӷt�Q�[��Q�؆'f��-ۓi���5��e�ȴ)�$�s����c�`��	{7����{��>��ts�ÁI8���ڣ`,������[G��4�����*�7�7p����ņ��+�����=hۄ��ch���9���d�6(׀��/i�/�Lx�nY9{A>o&��2z�Qm���Q�Y���.j���e��tu�Í�{�3:���6��1=i��&5$�����.$_��/�2�� ��*nI^�φg�l˷Vu=;�N؋+�Cɏ�t�*����
���Ȝ�w���(��O�joR�}+]k{g�}X��V>�o��>��e�Kw8�!�O'!���y�:?�8
{І#���/��S
�ڦs������מ��C��9��v[�I��i� ��ɂ]]�'��.u		�Y6�1p�l��qTŁ���	��^�;�p��0���8��ſ4~��z�cV�(��� ����*-C+�В�ΥV�v6�W��&�6���^%�t���������G�EhB|���=�-GB�F�B'�x}�|%��s�3/O'�H���*g���4�s?yv�=��z��I�_x��yή"�3�p� ����Ę�L�gOǩY�)����K����3�"��{n��L%�8�:h���P���p	����BQ�3�
�Ͽ����{�^H�Q�-��db�N<K+�#��3���XR�萹͒{4A�*L�����v���u�K9J��k̲�`�G �I�!
˫b������t����Dr��^vG߸�kc%��3�z�G]�:��2b��b\��� ��H9�h�H*ܩSW?�܏%6 TΦ_�M����,�p)�;w�ڭ���I���@��.��N���q���m���ެ)Ҙ��ɘk[�`|��*�
�έ����VZ?�w�3-�뜹"�Cƽ�d�ƴQ:q���4�u#�e����u�t�Tn-vikX���^F;��u��:�{��CY6h�V{�L�l��M# �]���s���v���z�8��:Y�T8TIo���(��s�m��E��מyם����k�*��F��L�tQjQR7���+b kbzͳP��'�#7����6�d��3��4+]���Q5�_��eטWY�YO�yV7����))ulS�w���=�O���K�f�K��NO��U��o��A�|�n�v�C���7�%l�����:W�k�%W��<,��0Ӷ�oc�u�Uo�)/�q�*���ƺ��L�2�Lkl�w�
q���c�yC��g*��`��87���Ň4J�w���*e%��t�)ܟuX��a��o�y��?}��zX6i��J�ցw�o�����"�]=NGKY4��\���߶:ga5�:i�x�N{�E�����?�e{���'���O��G���_'���6s�~�\��&�&x=�|���z�y�|�q�s�Y���E{���g��'�����O����mv�r�V���@��A�A�Q����ȴ+����gA"'��hi��{(�a���:\�^-�mP>h (�:���)��O7Qe�?�_���!R(��:�$�̴�{|zĽ�v�\mn�h��xJ{�%e����غoc_�*���6��)�O��x���x"�r�h�7)��J+��W�&N�Ʊ�vQ��K��W}��N�٥�ӱq�w�L'�?����˰$`�7�X�u��YW6y4q��2�V��4Tߺ��?~�1���vk��q2�AH�K�e����W�ѡl����<���Z6ʙ�P�ؒV���N���k����7o۫�or��X�҅��¡Va3��p���\���'d���D�;��xʴ�㣶���^�y�޼{��W:D�l�@�5�XJ�� �H��r�����CrʵMLe�d�(�����陛ã��;/�9��B�P���0N�Ζ�ؾӑ�n�H2�G�A��J١s`��)p=ҩ�q��+W]Qn�=@�@�|����'8[�k7�/֧>!�wҭ����g��A�� ����;i2#Ψ�
YM;�QUK݂RΫ��׳;��sa2�-*Ãq�$���[�Hs>~G��u�Ql����Gٜq��@���t�gW:V���}�`�`|�uA�ʡ�W�ǎ�0v�鵰\�'�.�QX8��� ;���z���U}�M'�H� ��_���T=S2���D���srl�Dux�1�'+�����Q�O�B�"���	R1�����CLf� ��AA�a}o��_��m�8R��O���#�r�
�*�z�y�%�BgJ�WKG�s�|��$
��<�86	
h�Q`t��"�/+�@x�ߠce�Ռs=0�2wy���_��:�Ѫ]ϯp`]�/�Iښ:�J9N���r�BC�Cp�m\?}4�{� ��
����B��8����!�wV�`%�{�ep%�n8��4�N�%L�̶��9��������V�������B!� ��O�Ϥ���+�7w�n�KsmG���q� ��E�J�H��=W�?,���DC!;O�\Il�T�u�wϺ8�~�\��ad�k[֊j��@Y�i��o�܏�u�9R΢L�]��z��Q����ו� $��n��bW���/G:�^�t���Q�n[Q��>&x>Gii���IG�\�"�E㜺%�Z�L8&(�����M��m�����k�SJ)�J�����O�4��'���,yTw�.��m��2/��VYE��!�r%H��B'���u���3�Qt*�h{�'mk{�mn�=�W�B�!b]�?u>\��J������Q ��vǀ.�����A��R}��P��6x�w��1�<����0t-�l������qc�:�3�,���Q{��q�>��_���"�N���64����<��Y:k��Xa�$h��l�Ghc�mtr�M�߉å����_����=��������ď�5�q��&)�鬻ܲ�'��.�QC���%
���w��Nw#��3K
��"� P�X)(L�ɣ�"�^#����_���<y������-4�F��&�+��8<:ù�o�[:X�m��^
O�<�O�Up=2de���֢��ơ�̃�����B��������z�4�6��gM'G���]|���r��I\dH�����Q\���F��z��K����(Z&)� ����P�d��!/eT9�B����#0�x��y�����'�|�>��q[X\D�a����G_�����������?<��|n���!W����E'F�t,W���ŹZo+V�C�`�V�uR��o�g��w�ő-i@���ex����m�2���X�����S��o�i_�m� u��N��l�g�N���{M�/�!�9�����L{ OC�lٓ�&e���<K�ױ=���{�
Mz����E���Ay�L{�\ �_y��Ƴ��N�:���~��q�i:�0����g������ !=�]}U!9����?���ix� r�Y�D�F]��]�4�!Yy� ��XV�~t:�+9ϸ��t�i��ż#��NȠ3ƙ�.;_��As�����������h�S鰰��MB�]�>x�3E@N�X%p�9����;0��:Z��q� ����e�O<��.��͒˶�:���k
/ c@�о���Rڶ��d�����T��#�[q��Yd�xU6*�{7 ��rh�F�٩�*{��{}JU�5�Ա�
@�NRr���]��Uޣ�J�Q�*����ϩ� ���wwx���C�0�_���3�����1��2�@��1��� \�t)�)�Om�X�+����ˑ#=�o�Nnt�+���fv��dG�Q�cO�p�}��t���אE�$�+���&��IUB⡟�M%8MY4�j&m�N�B����BD!c�	!e�
�ᠥ5F�5i��R���oedh0y�r�m-�i��C�ҋ�0[�Da������͝q����^R�C���g��E���
7����T�\Ĭt4��c�u�0�}�b����G������}h��8���c�q�j+�҅�z)d!ΰA#B���.���#���L���ypXN���e�.t�R쮼���'��	�ً�Ekj�+N^v�H�>�=������*'�Tj�2�.�W�<]iW9������B&����h�|�
�cH9��[ʛ���O�=W��y/�Ţ[�¿�u*���@ܾ�Xl'���\��V�?#q���u�8Z��J�P�BG�_8e�ڲ���!�n[��j[;;Q�
9�*��O�
���!����P P�yZ`|ůz��tNW`%�g��)Ƨ�H]j;+�O�j�����v��������ӏ�a��S4�t���,b����8?8�Y$i�����H��3�[�8���!����B��Yn��ڭ��������O?m����ݾ���q焐vM�/����`����{yvr܎���#\�G���ꃕ5�²B�����O>�S���o4��J@.zo9��'��߇5�] �57���9i;���.�ao�sR��UO�� �+��0nK6�rd�.�r��#U��yh%rP'+��D&��Ω^����Z+�e�����Iw�ۆ�r��r�>��ֲ2��j��2�C���O����S����4�x����-��Ȇa�춶7v�����F��۷ۃ���'Or��t[`�zu=�	�YeH�@x�N�`VHM���=�_c>�<�9����.�a�0��s����C�R�j���������m�0�m����)���j��i�N9q�����ۻ�wݨG8U���_>\�4z9���e��Ck�
�^��}�2�CХ��v:�pX��v��U�^�pϷڜ5�B]���rG���yaio�z�U�-����Ց|"ۺF�.h[��Fm�J�M�$M�_�<-p�J	�7�{����<���#�ꏀKXp��j�z�G�c�� �N��I�8�s��Y��ZMp6W/��s����{:��C���������7[pH�[�j]��׃"SV��F]�W�/��J��X�X�8\ [�3�#3��>=�!�i�����'Kh�׽��L)���>���ƯF�]������Ug�tf0�I�|aM��vw�۫W�ۗ_~���������mscE�.D���+�e>�b��Ԓ���O(T��u�'O��R�����P�^ؤ���y�s_���{���b��G�H7��;���r�H{?b� �Lh���t�Т4��I���+UB(P�� �ע�8����r�;�xL�U}0 ����$]D��ޓ��xԖ�ZhDf��5a+Q�jL�(F��� '˱��83؛eW�x�[���n�e��FY�J�u	|�%n��q�&�;�&-"0�93�"��b��
���L-\��0uE!M��\�����Ңc�q�L�=�lM�,�M%�3�e��.(��r�d)�s[z�B�J�'A�{�=��B����:���$R���}�U�c������+B�y�qVaG����a�`O��^��a�h� �,�#��RoWt,xO(g�b��
�Q<t}�������/�:�V]��Q�H�-ˠ����v�a
������u����q��1�(�Ű��"�f�i�b�����,�����t�R�3}W��@���$�b�U撓eXH�'cW�K�y�º���t�[�1�v��ِQƥ0�B�,<`W����0�p���N���^{��gK�F��{�A$�e���w�J���J�����G��
7��τ�:�F1/ʉ��q��o�
[���d��|���AsO1�+,�D=x�G���g���y�}�	r�t>C��ۈsE���+ͪ,�	�q�fV�3������0������CW}���k���]��p�|�"��ࣶx�N��vEUWaux\Ѷ�T90��M��P0w����6睬2��������	EcX��}��:*�� ~�������ݶ���6qvv]>�zuc�̫�;��9�i�M+�� �8�����P�~!�{�M�N�RG�D�!�>-Ya92�4�Oy�M�<�\��,=V����V{�f��}��޼]�~Yi/_�i++�����U���h���v2=�L�1}�I}�7}#�Ζz+e� ���ol��P�mo޼&�7����#c�ki����r���g���/ړ�O۽{S�C�)W�	t��q�L�˘2$׿��wAü����ƌ�D/#QН�"9�PHxd�5���F��d�(���-4��w��JGY�$6��V*���4�{�5��N��v=7����D��v�����u���3"����hts]�ƅh��:h8w6v�VH�rea�����h樗L3 ^�8��-�OIu"ӤK�SW���y괎�\�]��U�^��vU�K�v%��q5+\N^����FJ����-�U&ȯ��U5��%C|x�b �s�gҐ�MoV�k�W/g��ݧP;�:L6�i��o\���%_����9ҹ��a��6R��lO`�g;�#���Y�W������݇���w�I׆ϲU��m��NCav��������mmc�m��
�w��˰3�U =eq2��C���O �Z^n�d����޽~�v��B`2��#�8(���6"A?Ɛ���m���\����cz��x���G�a4�"�8s���I�V��r
d�/|���/�
t%F��4+�)�C�(��^�P6?:�b���.C���A_`�_�
�Q�b�_�
��lF���R���D;�� "���@��GGeXC@��A��T[�ٸ}k�=|p�}��^�sk�MO
s�g�Um�+��L�L�@ĜMGak>:¶L_8i����􊋬��)Q��a�S#�v�y�1Ht�)��p]�BZI��]�:M2�p�Z
*�%�ƨ��Pt'�C9\Pe�k��u*��t��⤟督B"$ͷ�C�K��,�P��:e+���
t	�j"BH�P{*̀�_{�B`"����q��Wu�C�����������s�3^'ʢ"0����>3I�`�tq���z�
��wHqB�.r[o�ֈuIfES`�ϣ?����h)D���um�3\�xydy��L�Ƈ�M��2��:=�꺧Q��W��%�,��A�	Փ�"��V>���CL-e @Ὲ��W�:���O�w:�1X�o-�%��j�Z������McRn�$iz)�ƹ�sa���k�+-g0�g):��pD���rx�����e���j��'�ɞ3Ȃ奥��?H�+#�H$F��x����H�}��˹
+)Y���@!w��yFG�ʧ�����ݶ6��z��`�]��#��@�� �%'��d�m�(6�-"��{�������v���md�<<E�p��6�_��xY�͇osV��kݧ:U��	}�g��Ael8|IC�	��֠�R���ʁJ[�m�x��oHe+�S.�C���p����ДU<�pP�/u�E�{�PA�P�?��'�>=����̄;��y��fNO����
��8o����8,;ms�mn�탋v�����p1��xS>���סVN �3�\g�O/������	w*dn��Y���;���h���V�Id��|N�$�� Ak�PC�	���Z���������|���t�����7uT?�@��2zOaO~e_��:G�_<��������")p������]����O���t���-�S	�����m� ���gmo�(�#�}i��9^��Ws����R��c��cy�>eo�B50��u~�]�1�4�s�L���66ۇkؔ{ѧ��j�	�\�p���|����-�l��8#g��CL��6;5֞=��~��O�l���PzvUʽ�ö����Wׁ�N�e`./��#���{J��Y�*�5��B����aʱ���1Y*��qÔyH'���:+��}Fz�O�9�W�;G�t:+�L�y�8q�͎.�^��Bd������$������F�+[0̆���Jx����(�eΑg)����%��l9�佰�7Mފ���/m��{�j(�t���w!�o���0=�>��kzH�Piw��q��������zz0�KU�my�m�*ZhKh����?J���<H{~�-�bDn��ˁN\��v�	t���mt�Bd�����6Ý��������8�|�+�I�)��ѿ/�\���db+�8ƻw�/'����|�-3��[-3�b
���ޮ������?���������믿jk�?#�������~f�
	��w!��Nm�,�F��)[�cy({�"�8�" ���ǵ���ϯ��DX�N���*�Z$�,@W�������Re#.0�8��"K��ppU�M%`�h���ݻ�p~1�t�`%ME~��i����J;�3�q�^�J�k��+�L:�z�0ѦfP�M��EBF�X1Rp�@=���5�|�{{�2ˠ�O�YY0-�t��<K�?���f���N�W'-"�����S:Z5�������!|���$���Sm~a�-.����1��(��6��/hT'M�ǨE����V6�����[p0�W�=�uU�#���Rp�w0��8�-JY�+gp��tz����v���r_,Q��n���>I7�A��>A^�Cn�b�'+��B٢ZV/,���C��S���[B)�|W���������^��}v�T�1 �p	�JO��k`gP_�=NֹN���*����ը`�e��������� 8d�o�y6�٧t�\�AS�EEF����� =i�#J&��C~�/9)��h��{K��CCi!���Fe|~�·�=!��N>r���
�⠽[y߾������/���:|�p٢�x��к���%M�0�A��0��]�]��Vz�Ne��YQ��aE���fl ���� +��K��r��x9V��
�Җ�޾s�=��Y{��s�c,:To�of�օs&�v��S8�p)��Uɹ�{���?hJ���wqx��1~��9�e�s��#��6��2F�8�q�إ��u�*v��'y�sEа���k[�8�[8��3�v�Jw�L*�Z~B�ऻ�s��:�yQ��D�nK6|���sW��+y������������������n#x/�Ygg�|tC4��sv��B,���fdC�����y-)NV�O�_\yg���Q�B��H�>{^������>y�,.Ա��C���h����_��������/_���|����<���(�O�-���k���ޣWgl�wq�r��eQ�Ir�����S�����`����ҽv|`�i�v����ԅ]^|�yZ�n�!?�s*k�S�ʹ{8y�p�.䩢?IFʁ3����YI�چe���9�1�f]|e�7���=�}�9�d��#l��l~�qj��HV:V��#eS�=�:3S������уmia}I�2K��9���y��N	���Ć:�8v.�i�I�[�8TW�o���:?=���S����'ޔ��|7���"~c�Xz��r�9�� �Iۅo�K�jN%�9���6�[N�5u���`��@]g�bz���2.���Qtx��n��.P8pW�xUW�vfF؄n;���Ց�R
�3��^B7�㙴�����Uc�k����6vh�O}g��M����2�iي��txۉ�N}�G�B����P�'�A��9!
Q��ƪa����~Ǖ3Ȋ����m��{���@:�y+���<��=�����)gr%���a�yd�7p�84J"
��s�������?��o���׿k_}�e���^6����m��
�My����,QYDV��ܸ6$�༯�E�R?��W��E�.���?���2�\�}�zF)��C�+�	�����r-A06���Tn��B�}z9D��. X��8Y8�� �t��VP(�L3�
N�D$
��.�~/+[��t�KWg��	{�df��Z?�!C
p�l%��ȗ( �"�+�:���~���Z#י�xPB��3�-�Y��P�&<����.]�vff��ty��P{��D˥�Ŷ��'kv�&Tf�`O[�)�uPq(<	��h�U��l��P�!X	/��EV���� ����w�:�N�.hb���&�'i�a�7�*��c:��u�3�/�.2�g>����[D�W�V'��z���� t?o�#U|T��K=��+���pp)q�N���?5L@������D�dx���$�����Z�.S�>jY���"؏q��3��e>@�����N>�/;���d!=����J�A�mi���f@I��&��	ig"t��m��qX���o��W:Yk�d9���P�!m�����/I�apP7|��[xb��f�#p�+uC�[OKf�΅9t��bYF��7���7䫼�Q��%t����-./�{���[�q��4yNP�1����a�n0��eÈu��u.�vu��;�����I�F!W��׽P�Tbtz��,�*G���w���|��f� ��7D�(C/��Y;Ĉ޳'uk+=|.U��ʣ�f�̻sw8�׏�����"�}��~�`Q�ԗ�Ds�����{��������a��B�m}��3:���W�(pȹ��)L�O�r�Vx�����,{J��O������d�e�m�����#���!�D�I�3\r5[)G���&�Ƿ�|�~��?�`}Ѿ��;�֎�\�Q9Z4`::]����D,��ԁ�s�k(���'�|o�N�/�/������n����z��M{��{����7o����J�H#�l٫���FC��շ�Wẻ"�T�H����78�,O�p���f{��u���o��������������#=>���N���K��p�����6����pG,��8biB;G�{��f��=���"v�+�)�T�G���#�焙�ϕ�:>:Z�A��G�����$n@�V��&x�9L�h�m�)�	2�q��!���|�C�пΓN����'Ƥ�x�q3""6 |��D��w
�+�N�-�Rxx�h���ز�\g&S:H�G��l�j����3֛���+�����{^���3]Z�@���Ȝ�W=V��W��(��K}����)c��ql`��Ķ�\�X97.Go�I׳2 u����U���[L�h���:\*�}f�E9b9�5Om�Qር���t��������kmu]����K�0n��z�p���vk$�\��i�q�{�W c;Nמ, Q̕anP�ڟ���&�wu,�޻� '�r�{"hS��ߏ`����2�0�9_�aE�T
fV�B��&P4<�c��h�쏴��!���o�^p�M4�8{�2��R@|^�!f	E%��B�(0#vqA`ȽP�����t4r5x�1�ҡ�0`;��
�#4�;o�J÷�7m�&��R�p�J6�3��A�
����4�߿۞|� ;f�^v	tҐ]�{�h߮�Cul����L[ZXD͑��uU/i9
��ؚjk�-)s<\%��O�O`��-S
K��y����L&x�M��+g)��VŠp�EH!�P�G�eR�-���U��`������g�+[V\8L�q�**{�fR7{G�3���.�8�SѮ�w�%rA��QO̒�g3T]R%Tʕ:QZw����4��)h�������t�4�A	L\�dTÂ0:�\.m;�'�cl�Ä�Ki	%`�axؖ0�8h��\���:c�p�����p���l+Ċ�U��%��de���"	`or�Yașt�d������Cf�6�)l3IY��u���OZ� J9���-�1���<�Z��)�����qJ�D��U��~�R��T=�|s*]]�������������=y�4�źI�s�֑Ao߾n�h���Lٍ�:�T�2P_�ZubC��<z�#�?8�(T8+s}Eyb��G08�������_#�6��. ��L/��YA�+5-,���E5�a<�K^��ᮡwG�
%K-�_�����N0��k��pC<4BΤSJ�zW�r�(�f;�ͭ%�Νۻ׶�޵��MʥA�l��ǟ|���}tr����>�|	��~�Q6~��E���H�C�ܖ�Ω����<�`���k�K�o�!��� �a@B���*��oҔ燑�"�3�.u70PfXu��4�g��:���ră�M|~i�Ol�u��Ĩ� ���3`l�,ҙ��RD�8d=�]`n<eg +�Y+�(�+p/�����@_.���P�n?��,evn�msc����՗_�����u�t蜫�8ӎ�����(��������!	�%�����U������9?1�x�>��"��f<����b�`�63��á!��Jo���n2;�&ы2�{0I�6~da��SWH<�K�H����)u��6(�O���Vu����Ω�|O�o�߳n�U��ߦ����9����6�޶�g����6N�����]y���vw]��lg'�2��w��c^=��5r���64>6�>���*6ر�����JZCo��Fp���k����8t�=�qg�e�߼}�66�IGZ�>� E_:7R�jJ#�[�}��T)s�|��F'��e�Z͵�唝���E�޿���7�h���q��G�����j��Y�����v���	��J&�O�j���<N���j�# ��%�ۀ�,s���o��gcsĄ���Z�=J���l�H�:�Y�ڤ��V'�Y�B�[}���3�]73�
��g�tx����G(/$Y{�6�@hbl�-�.�\�Pf�[Fm%�)[u��v-��\�b�M*�B}<�R\t�\䨆���Q��C�S�f�����RsQ�`Ք#����6�"��1iM>��K���X�S����Cg�Al�NtR,J�E�	�^����md����f��S{]��N[������t���<;�̃�H���Ν����G�ދ�
�jM� �Z1�甸{RJ�����*l����X�\�5lE�D=�º4���C��"Ȭ}υ�!�2���o�i����K�?�������O���]���W/q�j����X��V�)��]�������\�Rߺ�m�s���Q�����e�Q� i&��~=�d�Ʋ���}!!����}�����d	{iI��U�f��3��d�C�Ã�i~Q�J�DT%5�P`�oY��`DiW�zO�ޠ���$]�0n��@�����G\�3�lH
JCG>#A˙z[6`%�Kg:�*��ZD����Jie���"}�hOc�ɕ�$�hJW�̳�ґ��	��O\�]��m>�'K��;��b��ugqH����*�K�q��*i���ѯp�������������O�]��`��q Ntv��8��s,�%��{��&B�"��8����Lz��W
�si����Q�=��[j(P:xt���?y_)���B�Z��U�P��8~_�u�@�y����ɑa~/~<� H[{�(�j��p�JyD~p����[�Rɞ�Kk]���ay�H�n�}H� �x��Z�נ-�x9T�RΛ�(\4�|�V��p�3[�5,/1��0jߵ�߿�����D���HDyp>�S��F�j=�]�.T�;�C���)?hVe�|�h��$'��N��_,��u�e���M�ڝv�w�F��{c��DS�+�=�T�\��Sm��Ν�my�6�p.|��A5s�`����Qu���T����o>�9x��¼�ːOO;\�v[�}�-.��cT�Hg�)n�p�qB`*��p���`<:��u���M�°>=؉l�5k�-8�v����CWrٹ>����\2�`�=�G�&�w�S�>h�2�+���P��%6 �cؿ{׾�����7߷��޶6p�����	�謹_���E�X�@����X:�a��ʆ��i�5�9's��Ƹ��'giT��O�x��bi�c ������Or��"���3�ߚ��|�`�,�#5vˈ3M����P����K��R��=�^k#E&��e�Z��(7~�����,�L͠ӏ2l�[{���E��?�����}����N�&<��ʛ���Y�(;cT��o�d����`T
U�6P�����f{��m���W�͛x����	�r��lׅ'Rw�н<^y]/�v����ޒ��ʾs��\U�^YN<<Yt�Ӵ�n^�z�g~�U'۴�#l�vh$�<����f\�aMs��Ｏ�
��4:x�@)]�LI�<������/S��2p�68��!������}�:�`1�F��+l㭣�l0���h�C!#~�Wʑc�p�x�Uq#��Y�V��o�'��M��ˎ�~�C���9X�Oq��T���/���C�)st7�z��l'�N��O�Q��(��u�Z��w��ܩ?u��}Bt�<Y�8���p�މ�k�x���B������#���6� q:��J�N�?m�*����{���"�'�!]����	��^~���}��o۾AX�y�&=Y[����B�V�@
�Y��Ah�#uI�SU�������ֻ�:��������#ڰɄ<�c�d��Q��)g���C�R�\d�&jd���0̚[�\${ŕJ���p��h�8i�Rx$��_e��HE�$�9�w��Q�Ǡ�������q�#�k�ih��Yc��E���("H�/^�h(bHG��e����[&$�P��̐��"-��Q1�yuפ[�B��g��cۼ�P��&�<�'�!����s����]G�)��h�&S��a��ҷx���	�
[,a���:J�s�#��N�����V;9�h'G�ͺ>X����s�]�p�.g��4����K���3�q�@a�edh�<�@��Rr*���a�ԣr��on���:�;Z�3i�4g�U���j�8�lQ]`����zP���ꮥe��Wү�(ly�u�v��p����)<ڷ�E���I��O�\nK�K{Ewuo9��˥��1ם�O���92Sy	]�&�?�F�L5�$�(���>N��7���߿F~��B�5���fCD��{+�C��N�+����!MPw|���`!���^�E�s�f%`�N��[*<m���U��Wѳ�p{ӡq{1$]|��N��M�J���ёsN)���r{p�Q���!rp~v?��U��A���}]��C�ϊ����o�4����
�pO�����/��%���;��</G2��}����Y��{'�E_vq�Vޯ�7��}{��5��0���?� #%O�R�)u��H�F*�l�rk�����3�Ɋ��_4���d�u�����_;&'�;�qwo��nDw��o���h|����`�`���Gp��/�54u�4�MXZw��-�.4�09i��.4��u�KR����*�W�����yP�K�^FZ���Fz.�P����~�G�R
ኝ£�K[�,��l�6̨�]DA��3g����wp��7���#p�CV^��t�\�Z����{���u�mLq[�1��?��<���S���_��/g�FE9����l��_�Wg^������	�羦n�~x�3i��:����� ��
?�w�	˰����A&�c1��QIt��Q�zR+L�-�e���{^9
J��p9Oɧs���^OG���y��ڃ
�;�G�<!S�hbi�dEd�������ɱi�W��pm~ԕo���z�|f�Eͪi�ƅ�q���2�%�F�fuBj��m*�h�gY�ة#�kX�o� hI.�,Z�3��7=�y���G}ȳ.n�>���+q�����vYI[�RK������!����x
�vp4�a:q��p����8��%A��y|pT�){X�ԗ��A`�\����g;/ʂ��=��yb�X��9���
�'��
���2	���P�|h���Ծ�1Z���J���Ҵ66�+�"(v�q�p����aeź"Δ��%B#�%�T��!7q�p����	�t�	\r���o!�ϯ;,GW� ӖCB��ԕ�T���a�)QI���:F! W[-�������G�W%s�#{��LN�2�8R�#��%_�N�
�����|#uմ)�*X{92fZ�{f
%0�yz�M�٢���5t혚�4$Tz�ڔ��,muC�t�B
�fb��%��u��q��:7O�M�2��z��z�v��JO�A�|�l�[�[e�K[�	��B�B�<��<0�[����:��:�},�{u~�����Nvp�p���q�����*�C;:�Ǉp�V���Z;��<����V�	J8�oC���q ^O��'oPG��Ԟ
�` K���Ԑ��y���[���\4�����a�]�>+!,�����/+�zV�=�"W�wy�ùBX��uG������"xN%GO_��滔��+_��^wi[�Ez�'�ԟ��w���4��+�Q�,JX�h5@ŚCҎ�����n{�v5=Z++���I�ߌ;�z�r��x$mp���^f9����(��"X
�9Y�N�^��gZ�:�1���rw�tr����޷+o#�m��p2X~7)��GV�nqb^�F/`�>h>n��<@G!���h���#%�)[��]�(�W�:%��G�,o�b�o� �y�t��Xı�����};e���$�a������gը�p������������m������~����l�__�jk����#�������5�� >�����k!)�5��2������}���W_}�^�rV-r���s�i��,8��1�1"u��,O٠���2�(�mX��Kc_J�JO��#Я�J��PotB�_<���y��qG�k<r#�F'@G��U�"` �׭�d���E��'˅tġ�*g\�����Y��!hV���;4�"u訬|���~��[�n�{w�;�]�}>�G��}K��^I�HS�"��L��4-�שg��_*����6���Ѣn�#�g�k��l;12E��8��Vvi����n�����_{zuL��A���R>"ʿ�:9q�D=iȷDI��+����B':[�]9���cd��2_�(��*=�7�H['�z����6?2����!���tǰ�*m��Zcl|ǋ{/���:����V�-���1�L�S�9@�0�<�yՁ�\���w:�_��}$�o�� oz��@�0.��. l�X�;z����>��P�\�!ny�=S&�����QR�;Φ��^g8_7�J��t��b�������9x��GWF���}��_N]�^�kQPN�#[�-�$���<*g>*G+�ԙ�s�d(*:�+4��T�̌'
3�}/�zc�����{�auβ�M���=2�3�Y��yC"�ɽ� M:WTxQ �P�4�He�����'R�!��~U�A��ﻪ�������d?�������`��we ���Qy�4��03ugOߋ�����/jrBT�0f:V��ս�"	��gl�á\E��F���ĥ�)�����Y�*�f$nz<?;�q�.#?7�Q�-���:��0��uQ���D�'��[T
nHWg?�,:''��#4k��$5y��g�(�_�y�������I�N�`o�$�蕺�`���rT�-z"��B�r��M��R��y��8����-�)"��c�+��8�ʹ)'�8L��:�_8W�{�9W8>x�q���Ώ��f�]��L�mq&�n��g���7qරޭ�6�F�����ɜsۗ��}O�U3���E����η]Nƿ��@��C�I��}=��^��X�P^6bR��7�']�P�W�F/�P��?�ڲ*#���6T�l:����x��hr���c�7(��G�0�z^y��i�
��#q�˩��5��m����ﰓ�h��E��J�8�D9122	G��+����
F�붶���?a�+y���(`��������zGK^��k
eM�8�$���uD)^��KO��+�y:����9(��A�����𪭯�����$ƨ{ߌ -�ɑxrSR�'���65�Ԗ�w�;w���%���e.�Ԟ樳�
�|�Q���G��-ӯ<���{�a^��͞�9�0{M���4v9�_���ҍŒ�T?��<'�mo�e�]�ﻶ��m��m�����sW�E�_�B� 2$��B86|���1��I����Sޝ;�� ]��)����y�W����[���h��ǯ�h��w��K�k߇�r�Nw��Ip3����;"X���w�� �q�ڃ���R+�]���8eVQQ<�!o�B�D�W+à�m�~S���ߒ�^�L�鹜��A�;��o�%�y(��߫'��Zg�T�.iB�νqnϽ{wۣGڭ�˙���a�6�*��q���*�6����r���{ۋ���>�Y��ŧ���ѳ�����I��^�j/�r����l�#��7�����ޜp�ԭ��pݿ���|gp�|�cy�m]E3��x*C�.ۍBBs���3�a8G���c`�0Z�)����9q+d�d�`����>������vpd+�H汏�� �u��/s�)_�y�o�T��P�;�о�i���v�9G�e+�M5V[�䷰��q'؅M��l���� 9�9�#ҧ��n �Y�@zRo��`��8Y��[<&�ؘL���eϿ{�j��,��(]�橍���D�c�b�p� �6З�E��8��Y:�n}T�.�2i���;:�s$���{�c����_}�V���%c��>-��k�e�Y�];i7��?�GW����kw#&���2p�e/��'txWZٌ���(~�a6L� ��R�0�e���2:��/x�M�w��~�+-�Ad����U��xR�+���c�u\T����5�Ɋ\��F@��B�"����C�����aV UΆ��yoR!��>>\'sሴ��4t}��*O��*���HE�3U�GbtN���-., XGLN$H���O��Vg��p
���m��?tB�=^G�Pg����0%��A�Y�8	~�ɲK'kQ'ka�-p�f�*�͕�1��iv��S�:Qxx���x�X��ɵa�=簌}��5tۃT܈�~�]�4�:��9�|H�<�g�V�2�{fgZ�"Ԩ��Li`Z>��Q�^~��$��|���)����(r�X�+�o���-��v���c���֎9�����v��t~R�Vg8L�8L���=�F�܅޶�m�n�uE,��V�?��JO���Q��o��ǘ.���q���CZ����#�'�#ɳte��xTZқ�~(�ڛ�r��Pq��,ՈRJ"2�P9��ru��r�&�Kw����Y:V[ۮdZ{p�^�L%iϖ�Wr���{���G�5�}O�QX�G'��VY��Y�zOz�� M�b��u.��8V�p�ɴ���,�9j��;ʍ�����J���o9�k�;��9�B���|�r����*�4%Ot���U��?��=�C(x�C,iI�V�^2����C��𲭼���U;:�n�����r�%�
�lp��u���P���e���֭mn�v�@������<Ja˙2�L	ҡ��5���q���O�;� �>T�R&dK�0����ΕM����aWh��­�QRtl1�k���j���w�1(�}�޾�&�[v�[���r��y�N���;2'C����:�� �-�7*G!��}�^0�N�?>:�g֠�W��n_~霠������������I8s��qd�χ0T�E�$�XW�o��+Cyg�#-�s�y¼(�d7�\�u�[��������
����c�!�Ž|8�竡�w��}�	�+:5l0��Q^�v9uĈ3��}�s��]#>��|>��8��ɓ'��GeO;�^	�2z�9����ޞ�3�q����=�Ct�����ً�駟��?�Y{������ö�T���>XZ����K}���	����6��m]JO|K_G���!�gQ��d�W��(�t��_���ƨ��ߓZ���v����)��'�g:V�Q�N9�q���sD'q���4$�샻��-�M�;m}!���$m9�P�2/��Ɩ�lK�$9����ؤ�h'�N�6@"�v��Dx�]r
G>�V̨�4�Is��z�����᪈60�{!���<K���X�	oy@�Я:�&�G�|�uJO�~�Nᡲ:B�����O#��(��g��4|�c�уeOE�tw�Ly����U�9�ynv�_�!_�n��ًm��n���9�Ps0��� �ܤW4�T.;P��.��>��*[W��H�9�J�^��X���!,�F�Oxh�ʣi��Z�!�t��LX����A$��U�2�L��A��>�;�����J��$�J��|�Xr�#'`J�
�!0kr2D �m=R8I�{5\�bk��J�^�PG��Y���q������ �y��Գ�<�e����g���7�t� '�� H���#Fu���s����p��(�ސVv��̶��		�C�qt��W�sN�D/q
7�̸����\�e~s*�)O�,�pV�s��!j����^��řvky����8Z3c*l{�Pz8Xq�\a'�?ʘ92�N���*�!���;_
�2�8�k*�t�Qz�`�\��0!4�OFpPx1���<5��m9W�'��L	+H[qxC!Y�RJ��Y�/��F�Үg�Q��H7TP'K�ͪ�]��,�v2��,=YN1>}v~�,q��;tq�϶S��1�9<�������^8�k�k�y[8i:j	����"(p��p�	�z�!4�;+Qx(�����t�:>!��rid_ʧūy�蕐�4��2wp�vw�14t�Tf:�%g��:�
>��-�̙��IxO�<S/ޛ��2�>�!G�$���4��+��$$������C#�]��e�4݂�u]����)��ߞKׄ>�@f���N��a�#U���NCn��+���o3?�����
��^�z�)��o��(u�q�ïy���� ����S�։���aBUy�!��ڄ�Ӹ�I>׉�7���l�w�j�}���������Qe�@n�sn]!̤������R[Z��u'�;ohXY����̐AR�H�4�W�t��	�]w�3�Ы|Ч���}�_s��<��,�H̵��}�8��iH��*�Ց{T���r��p�-���U�x�V	k���ƻr��g���="s�@M�4�)Y.���(����M��ޕM�p�]('s8y��fW`;<�M���Wo��_}۾������oڻ�k�C��!��h��z�r�v�
���=��/��c�s�KG=�ˏ�E�V�f�Z��P��_l]F�ِ� ���o6M��r�^����y�\�Up�RVp���5ܾx�z�;|��8I�}O�?���Ϟ?k�|�1��g��>�9z��ݻ��=�%MxT}JF8��>.KG���:����X�]De�N�s�nV(\^^�q�zQ�}�G9U2GY�<)������q�"���8a9~���)/��K�
�[�T|d����{��P�j�;M��#���R�g�<��g��ئQ�|u�������+��HP�@��g6�J��+[�4/� �F9l0���v�}B��l��a�8���[�HA8?�y�ɂ����=;�y�V=��m��OP��s���99�l<��׆�g�F7�w���~;8tz���#���1Z��,���� �ЙM/�M�.���j�l�6�ý�i��='��,����;J��N��j��6�qZ��ҩZ�ϋ�i H�~y���k:��8Y�O)�|Q�4(����k�,W�We#�q ��y^g���:����p��ѽ��L�Q�R:}̏�#���w���F[ݰ��X �r�e@�ۍ0E�=%zڢ�Ve'%+��H2��-V��X�0�D��ي*���`�\lm����1�H��y[{�|���Ǚd��y@�5ԡ���z	�5xG�!�.���ݵ�m�О�7΋{sT/��lzւd�崬Fp9��-V�|)GbhD��~�%�� ���me;?ߥnss�C9S*
&o��5D�r�w:��n�裇���%�Dn�m=:h{����=c�U�8�2�x�����C�J�����h�:�cu�!�|�a7w�dck���据rh+�Kr^1�FCm�2�J^*xp��ȼ��@	I�K�2�x�Ϗ
����QIN�h`.��?���A�aL�3ʮ�eV�3w��-?���m�M��M���+-iz�}���4�w��C0�bR�(�dUdt�O|N�I�V�!79�%Y#��άxlp�@���8Z��.G{�c��D�!����=.������#��Ә2�*���7�!Z:���(��k��%��^,
m*T��}����g¦��-�Uk��C�q��D�"@�kҌ��h9ֆm%����0202�9:#1�ɵ����oJ  ��IDAT�x��x��s�|��㚼ő2�C��e�5�5tf����{����>k�+�V���j���F����.{�c�<U�H}�i��.9|%�H�W]4 '^��~��G�L��F9j�#G�5�>*I`���=~�j������o�����O�4	�zG��G���!��Pq�[����|k��ux«}������/��7_���U�?��8P.�c����*�-�iń�����?��-,���4�D��tޅN�4]zAZ$��i�o=��u��������'G#X�f��+t�'����6:u�ԙq�����:�fx�����y^�S�M��lAGz�'r�+G���F�F�G:C1��S�Г�g�|�\x���pv��vrb��a�qks#<�������/����+�N��q�Y�¡_���ad��{���d��Kי|!b�ԯ��L)c����>=MA�T��L�g��8�Ր&?�8=���}����s���^NIW�O^�����S�Ka�����ؕ��H���yZ7���F�}k�=F?������������t���f)kt��ѫ:�ƛ������j0��|��NV�otQ��A/��j���T�"N2�(0�QSʫ����"9jϔ�䰾�n��;���N�{0�
g�G���(���5��et��w��<Kdx���w��:�(�W�����*M_:dT�=k3Sc�u�=zx�kz���:iۇ������z��ܡ��1�rJ��)sޗ���]�|!�I�668Gԩ�}�7/��T�A�������#n�VK/�������v�9���Vm�#>+��ҙ<���q�)ɀ P8�Z�Y �V��i�+4*��]|{��'O��/u$�>mP��_�s���mܨ<�a2�p�?p�������ݺ��Wuzj:=�.�'Mڨ�=L�O��:WY  @߿��N��r��н�6������L��\��S�����w�]�?uXG���	�cx�tB{F��761Ӧf�+S��kS��a������9�������_���}������rLaA��ak]�5����x���H����vۤ���(l��0�K�T��-lω�~��!�8`�/�8#1ޗ�z�`}��GN:
0�� F�A'�"�����UC�D���޶w���8J'Ow8U@)6��Խ��ꄎ��0L(ZBC�/D�
2�N��!"C�y�PꝬ=� f��TV*��KVǲ�BÈ8��9�aiq�ݿw�=����C�*J�߹V��m�8P*)�aK
X��bg�d�`u�L(S�:�G�"!��R1>٦�I����o+�8v�r�4��ӄ�ʹ:%�aX�9Y�)��O�C8�]2w��&��2Re	T�Q��\���=?M��DK
�ͷ���v�E�t����P+|� VY
FF{'�#.{� ��[�d���&Ť
'a
d�Q�N<�I���R�c'K��I/��RO}4��%,��Z��ڐ��ȸ	�'��}u�c
4P�Z� E�	��DfL؄��*mf���:�M�������������9`(�Սw ��d	lt��R%�tk(�b�P�=�� ��iԆ������x
Ho�����o� n<�\���*�\vxiy9y:�G����z��}[_[Ok���!X<O��9��vC/�M^�������gF�s�v4g�Ut�l1����:��P+;���BW~��qzeg���|�P+� ��JQr�pN0B�z���_Ή� 4�8�`��6��s9���`'�=0��}���`mn�������J��A��|MK�g�J�3�S�np��i.{��s���$|�d�д �����:̹��q���:����9��yZ/8�d�U~6�Uy��%`�
m�T�������.&p8&���c�k Kw'-NVV�����U9{sܠ١J�s���}�(�E��x*|�� d�>����p�V��~��o�7ν��M{��C[��j��F+�`�L9���Z�,,���IqA��h u��Ј�?�{���4��=׼ŧ�.b�I�K�&�|S��w��o�i�v�_5�Om���\�&N�J��ؚ�8z��ni�%���	�������>����W?o�xў|��=��޹��ՙ�aZ4'�e����V������h�r<\��F����{=��y���{4�.C&�[�@�V�lσ�4I�5,/+'��xBҐ�z~�0ۆ���K�.��R��������=�g:YPq�o��r?��(rz8�^�w���K���)��$v�{ �_���d�\�.��eOq������j�G���CU���+xxޡ��i�O�Xy�
���Q�w�gj!P�#�Qv�z�x���c���=�}}=Θ��z����KHCG(���OX��A�ǻީ2]���g��rD#�rF#�W5>P��m�䟆Hu9���*]�KWMvOčߧq�wi�vUGq��d��ͦ����[�����e��Fԁ��m�����p]kcE�QW�/��i����c��x�,'��_G��b�����t*~�[�M��N�YA���>��5]N�����?p����봜��ǿ��w6���^��uVV
@��;���p<�C���ڱ��8Y�TT��_J`-�c ��b�a�_D�.�!� :UD+�éᾀ�so�1����'�r�{�6��ç1()Ii�	[
7W���+�K,��p�d�p��s�i�B9YԊ�������G�!p�9e�JE��x��F8���>�|q��eKBY�1F 9Kh:ZD�`��;ZA��	�
�E�ͻw@��-�m����i�,��!0�������pu�8�&Ƣ�8����°�FeIM
����([�&Ł�7N���p�ys ��F�i Z�Q���:'KF�o?V���C��r��~S=^*;��7�-N�J�g>���p
S8�K��/W��ɗ�U��V��gm����3�,�U/=b�'aP q2�9YY��Շ���4�w��0�sq�gֻ��Y���"X�8Y�Öc�\�9��s�N�Sq�xqj`
Eh��;8�vH:��u��_`'�34�Q!�l�wZH�҃e=0J�
�3T)����]�������H���T&����I+��J�Q8�=Y:����9^+{̀�"{Sc�?i�ѸDad�Q���UHʉɻ�?� #�����(�۷o#4oG�oY����P�ݹ�~~'�uK����}�K��x�s�>��W׾�?��+N��-��s�#�'K>���)H>B�+'�!�!��Qz=T��n&����K��0�-�sB-��|��*�1&�r����������=��'�\��:�M[y�2�ߣS�S�C��6�L�A��C՛��3ʾ�e�,��Y\Xj��ϐ;�F�f�Lz�Έk�1<4����@w�a����ß>:H�����*�I��JNX'J'��Υ�������j;�߅�1y7�L���FIi�5>3��t*t�ML�����$��!��3�k�w��1��iM���!h$�-��Ycc��.��\ta�m���_i�߼n�~�m�h��˯q�ނ�u�B�#*kNI�xj��"�R'�,����f�u0��z߫l���D���8<+����$���CgBY�ɢ�����!��\=�4��>���;Ӄޫ����t�4�6�e��J��`�<�7�Y�������_����?o=z8h�� ����k���9�����a��{�.K��p��G��t����@�6�P5��wLbK-,d薺��d���[o�9p���&�8Y<Ϫ���9L.�!�i [��i����-�S�
g���:M��g�Ţ�՘��c�k��4(Djp�%p�N[�a|W��h��q`��ٚɪ��E[�{g�N֛w�mm}+���м�R>���h8d�F!yPRɦ���a�'ǐ��w�k����W?]��@:WSĝ��x�V�?9�?k�!yDOQw��a~s���2����gp��}śN���x��u���Z�!��B��4��dQ$��<��-_?L[~�:�xS�*�\��s�R٤\>:X=_ȋ�L=�^�栵yh�!���o�g���\�B�����Ӽ/�$�ki܎���Z�Ş,������6��)8�&�Y�I�ҩ�H�'�A�^C�u��G��8Y�}O�Ll�8Y8�:Y�-'����������+8Y�ܵ7��Fh�C}�z�n�.ځs#� w!P�ƀ42Go�	|Y���{���  y<=�ё�6��w�~��Y{��E{��i{����죏�f��ťe�	�]ʘ�Fh}��Z��l�N�>U����޽h[��mg�����W�N��p*e<��J�Zs��8w]�~!�C�3��� ���pu�b@۲�0�3�F��/1�5����+y�8D(���1YK6;�%Fƃ��.r����R�$,,�'���h�q�vQ��da��TT,�2BZe��f� q��?TZ5R�ԯz:�n�x[��� gfl-��� ���n�ZRNd�6#��aq��h&�Faߛb��{�B�D�!���ٲ�=����zT뭂�R���s?�鉙6;�H�б	�O�4s�p�q����w�z����B,F��Ȗ*�{���-.:[�_R>R��X�����)=�^#��T��q��u���rueO�.4��N�\��[ma��X��]]A�W�ouL�p�I��<@�<.�
����J�h�y
�iDq�Y#?�V�����rh�'�r���18�!�ĳ�9��JK�L��u/��B*-��xVA�1�R#qlL%b��s�e��Fa�pD� ��^�K_t4蝓��?�	W�!�s��e�!+��<�h���0�8LM�"���ގ��U��g�8�z�?1.Hϐ\��4����ɹ��^�� 8���A�8�|}N�2TH<ȩ�h��C~��H�m��%�mlĉד�3��l�u�X[w����˫&��)���.���/g�+�cRI��`�p��adBV�A{�Zm[������mm延��m�Z_�q�C����%_�Dc�2:�a�C�Sm�v�����C<�s<�2�f�i��&]
�>�_f���t��&�|Y/��x3t���w�����i�Ġ���Q�!ƹr��w�����x�����QA��d9�r��cp��ΰ+��@�.p�jc~#Ϻ��ҍK�A��<W���:�$�#cW�=��=�o����w��������m��B��v��ޔ�������޼{�޾[i/_}�޼y�c���c?ll���vr>�N�����pC��m���	�%�qd9�=P�vA��t��a��܆��Jn�Cq�~?�Ɓ����{�"����%�E��k����1�N�N�[�wi�h��k��9�#��IK	}�	�<��C��c{:��j"���ϕE��y����'����/ۯ	��x��<Iz��!N�B��Ҏ�#Oy���!����X�~6({J���4�S���;gԢ[��S��:��]W���v��6���vq�׷��p�& �	d{�b�# ���^.[�9�#U��A766���`c��|����>RV�+�T��9�Q=؀#�ހ�L�;�jq����!��(�Q����H{|�����ὥ��8�&�ؼm}� �����+msm��R�	����ʹG~��a�"Oű�t
-] ����'�ۯ~�i���g�S£��1���V������jS��<�i�?y�~���ǟ>nϞ>hO�?lϞ?j=v�H�r�R/l����g�?��>��t�}����1������8_3��������	|z�}�p?ʛ�[М�]���+�3���'����6��:X6ꄮ�O�A�Z���S6���l��gB���P�0����V�C\�biѽ�n�9�2��(y���c)��C檟P��p��r*�ΕN��Ѩ�2dpg[m�g.�Q�U��6�E�^<��3���qTV�K�����~Iv�&�	f��,�
liQǙ�H;>�#ש�����C��5���]�r����	��FeJ0L�w�T��`9�
� Q��~�4�?p�x�R�����wB�C��0ć���"]�����g��>����ٳ�[���8z� �`8�b��1H�iĖ��p�*G����U�۷�'�쫬��ep�^`G�h���'����Np�� ���Ǌj��ƴ��΂
5���c���2u��7u���.���w�0����!�r�8Y������&F`�r�-Ň�mwBu5"�*��-��_��z(�e$���9/UW[�h��#�e�'0�2|���A����E�b�R?�
��F�� FY�٠Ů=EO|E���DeL[t\�ұ�NL�gU���tg�Ҥ�Tu�%��O�J<�3��#�0���u��mcHom���q;t�-H��j�K(
�`H��a��p�T`X�)���,�)��N�UZI�⑜BL��3��B��w��loVmD�y�;����[A�\�q��Q`���>8 q&H*�*l�G5B�p�F\yɠ�^(yY6�G�g��.���5�,P�T�J��{))���w Ö�����퉎F��P�'��%�Z�L��[��e�����l���Rϡ��$�2Kެހ�����������{j~jk�Ʃ�}gg���k=���z[��Z�Ar�p]���8}�k��-G��s�u��e臗�,���<����*�����Q�	���S��N0mp�WӲ�!�������a�7�+e��~��c����<�s�����C��mm�b a�c<�"��n���
MH���뤤����[w۝�8�n�x�ո	JTe�<����R��N����O�����s.|�.=�U���`h}��:B�>�����l���x?�l��K��T+�ymZ�4y��[܉{����3GÞ�cx'��\�˹Շ�X�N��tx��쿵���C�1��67���ʇ,p���a�j�!<n�1=��S�������N�)����� ʫ~�e�����t��,�`��o���� fIO�5��}�|3N�8�McP��p࣢^k䥬���T��o�����,+?��?q������ �Vz�����ϟ���9��sx�|o�]���߳U^��͛7qd߾y�a�>�f)�3��t��p8�����:�p.5��E��'kjz�m�l`�}hG'89�0�'�^,i,0�`"5����.��e�3ؓ��%n�l�G\�	�ޱ�.I*�����T&	[m��#���Au�=7x�i�©X��l�����W���w�2�X�Hb˾���>6�姽�Br�ܹN��u�����ڰ\�q����\����/�_�~����Ƀ���=l�[8u��������ѣ�8HOc��c���O�p���&��<DF�nK8g�:��ړǏ��Ϟ���q��/��O�\=~�Q{̻k��9Wtn*�{K�(�kH���.h�C٬3��2l� 0|dP?Js�:�:X��9���>����xօ܈7��+�$���:|�ӳe���a���@���h�g{��@��?�kuS|�qޮ���p��&�@�EW��xD����o~�w��\�|��S��S [���q�$��rE���36�a��d�n�\���kO̶���ayr���@ø�1.U� U�t�F�����R8_�=F]Q(+!�c��P���/�е�B�n���`	O�<n�F��_�`��s�Y���1֎��Ę��T��`�dMb(���f)�ʆZG����:Y8X�����B�d���;Y������NV��#�QuX��(!����:8�N�=
5\Pӧ/DUF*b�ƯP�Q^ꩣj��F����8[��ԛt]�����-��L�sC���	����$)��_�YR��~�Q�X*�!�ُ�v���w�~q�:G.C�٪/��d�~o,	!��̕"Lʘ:Y�O��kYe���`9���s4���⪘�V˞�i���T��FX�;MO�(�-�
潽������ǰ�E`T>:Y�jÁ���v� sr�2��]S�X^�IW����ɂ��Ѯph���%�2��x��yW���.N�6�}�I�{�OC�QH	��>b�R���DA�VϮ%VERC�zB7�e����霬�y� ��9�RV g�'פ�� 6Sw.�]�����75��~//I���u��+��]lh���CWf[��o�(
Ex��E|�uN�QW�Y���PI�K��q"��;�������G����J�ʾ�}'޺����bե�T��O>�K:>��r`�¥B��<K:���R�ʪ�ǹ��1m_�qol�@��+�'q/����qz<PL��搡3�!�!nF����(Vs&��[�'��=�ФO��[�	��P~���{��������m������h�X�ޘ����4Y�Ӭ���s�����|[�}��",��aA�H�,-m#��3:��+"l:��?�����ßq$�DB�R��{��R�.L;�<�ɒ��p��ww�۫����a����rɞ(l}��w<�U9��3�+�38r@T�Y8:�!�6����wb/r62�������N[]]��:&�t���.�	G'+C�ϥOe�21`'t��GV���ٍ�����y�����X'�d�����C���8�:�!bWO��F�rJ+�C��*f�Zh:����7#qdH��a���8����)G�T��ԁ��^��s>����7�Wi4vH��t��[y����"F"���C�8��ݻ�8	8�����񩎖Ԅ��M����	�d�Wy��oe��[����n�7C�����d�^l���_���0���hz����]	ZY����/읊ܰq�F��O�����<υw�� �k���9��	ŔyL����J�8:e���{�گ~�i����y�sk.��\�.�^�2�lXb�RG*A^��pޖqvn.�R&M�S�#��;�׿����/����v떍ٳml	GɅ�t�޿�S��=�az�S������2�^�����p@â�/��|�o��L=��}��q��/�n����s�@�A��/9��֭%좑��c�~ãvVs��ʌc8��9cna�T���;G���=��M��Ɓ�7���AX��ޥ����^�^�2=.����R[��֡�N�й:����
��ۙ�X[ذ���W����|�Z��=>S.�EN�om6��<��/	�P���	-�����\��>Lalr���/g	�~�/��[]O���X=�����o?p�N�HBe�ɩ$�:�oo��?Ĺ��ىBHK���01P�^F��4�5z��XS������1����/�����_گ��D�f�K��J#�$�e�G�V"�im�vn��A�È��";�l�ty|:L>�(�s�g8��dEl���G����c'��Ǡ@ݙ�����d��ʐ���ɪ��h�E�\����kY����OA�1�<#�,87m~��k�A	��´���W�d�̩���'�T�d�[�Xjt¼�$�e�.�c����PX
#�(#�\�:
c�@U��%��uR�q9R�e�*�{�Gb�+��.��?y4�{'˕�4~ŋ����8D¥��Q�ek��S�6�(�)����+����#��Pt�1�
D�I��d�)pq�f�,��J�"�O,
qY��!@EO�1��f�1>�����L�#�h��9Yv��Hd1
!M⼓fᱜ�~8�G	Y�قCc�*�� A؅������>U/�A���F5<�O�Ϻ4�5V�9s����SO�#�A��ٴu��������¿����u+~�F�w�h�#�:�8H��Y�� |�3C&x�|���=l�I��q?�I#M�1�?9\P��19,cU4�ʣ��iǀ0���郇,�{��!x�/��Flpn����^p�}'��)�����;&Br���R��y/�ИF����c�JPe×`�����'�Zyf/��w�O����s��G{;� ���s���m|x��?�m�8Z�x�[�CPT(�ʻ�V��t������E�,�e���"N�ݶd�/V3���̳���6�^C7�N#��y���zH�ٟ<�pW�Õ�b��/�)�AI��T�����z�E&�_��0���/?�m��`��7=�; x��wDB��<l�p��sh��������У%��#���5x���9Bm�uc���#3��B^�@�bC��Ut�*;B�\���^� ��lҬ����m�\�s���ܧ�2�u�_���K��#�.�	t��a���&`�#a������"2Fi�T�,ō:�<ß1P����vy�����%��g)����T7���o���1�gf�M��y%-T��	�3WO�J��8��bhj`jlʋ��C���u���ij��^(p��^�#L㪼Zu���Ł�����_�,o�[h �hs8z�_�I��N���T��������I� ��G�:��N�<��_�:�� 0̼`�	#0�����57�FuS�v����{�#�W��8Ys6�kH��U�0��������	��N�L8�"/�7�vN�zGmfj4C��!��ϟ�p�w�#���IW��6�L/��[˱_u���u��e�������ӡ��Q�ns��䨣;w�q����ot����2���42����&q�n������|�.]���D�X�0.ٯ�V�QM�(b{��6�	wG�8]G���V�rԌ��������+/���%_|�m'&��^�ǥ��A�A�J��X92����j��ͭ�̷��\�R�^��t3@��W�$�SuV�Q��bٺvGx�'�ѻ7ޫ�st'�>15��u+.��=�;sڝ۷���N�x��_���}������X=Y*#7	tn����/8�B�[�����p�L*�` nf�y�� [Aj���t��(�V��������7��w�}�z�I=��e��� 1��r�����S #cz�,iw�W�謜,{�vq�����s�d�����A������ԇ��a���GQ�䦐����O2+'Kq�de��9L�RQ ���\h(�� �m*bE�35O�,8A|�О����;G�*#��:�]�b�L'K��AꜪ�:�m��@���v2h��D��`Ӏ��S�g�ShH;e�*VLP��4����8Fi�|'�&N��|.�d��a���|/q�����A[-�vU�,����1���(rT����밭�m�-��C�GF��:Y�7����3���S '��:��\ F��!	B�n� ���,~��ؼ������n�	:=�ɢ�Y���j4[�({B��R�l&�� =4���Ç���Fm	
�2�W`#��`�0J�S�5���K�ץqH�uo]}ZGw�Wtp@o��!]�EE����qa�s�^�s����^�(���ԫ��4�����e�Iޢ�9�7��IߖA��4Y�R?{�����r�CLG�A�0���v�X_[E��du���4m}R7{��I��J;�?�p��WY�@�p�]��AX� s�(ɳ��B�.)F�d5�pMԴ:��°�n�����̫�q�w�������ƘF`N�!���H�S����61ڶ8UV��Ԧ���[�˹��x�v6��}���z�� /�����(>^�UU-e��tLP���N�Ƈ��5l�z/�0�-;�W�9�0-������+!w#�?u�P8����G�����K#�?�G�S�s{��3WX�	ՙ>M���U%lZ6
�Ou�8N#F����|����{52/�o���%�EB*D���_�G��e����>��6a�m�_�����I����#*x�������'�NL�,G?�HU:���=�{y"�(G�1T����3G�h�8��}�u7l(�6�h�e�7L����ڙ��ǮB����Z^q)��ۢ)�_ə�˫ccC�x5^�T=���O>~�>��Ei�+C��D��⧽�6��v��kXk7�C$��]�yX�*l$�8�s���̾�U��y�9o�"_�~_c#�de�=�q�v9!��8�nW���'���'/iCX�8X����ƅg���j�J��u�"�/�V��E�m��������X��]���h/�>l����_~N�?x���t�v�ή{���a��o&yR~\�ܹ� '�Shj�=�����ϰM�%���!x�\����|s<_�w���\���C�dQ�t��Ϭ�uu������Q|.���:�:b#�l+��8]����<u�Ơ�҇�ll���L�,��s������M��vX���p|m�a��}��Vf��ꈑ,�ei���;����]:$��s�ͅۥ"���6:��ār�
sq�^u��>����:Y�Ngl����S�C��	Ҵnq�ltn u)[��Y�3(�>7����[������:���8޳�m�����m����u:ߎJ*M)b72� ����UNl���2��Ŝoɱ��$��2�b(:��F�	�/]�!{<--�{��A�w ���qpp�p8C���j@���T���uy-�e*f�gY*�7:B�P�z�{x����SG����a����rܼ���=�^)F�e���,0���l�'�pP�r����Tݨ��U�et^*K��^$$A��8$D��LG$A'�yK䍀�LT�*B[Ӣ�BN/���
TQR����3�6TK��A�#E���!�Z��m�!j�J+�K'��	r#��2;��Q��?q@�W�ɒ�(s#
;a��mqU�:���{B_*(l��ڧ�P��:ӺkD�C�Z�G��9I�d|��|�Q=Y�� ��ܥ�(@�\���ßYj�i,�k����>�|���Ҟ��4購�Ը�o�&*�*��o�ۦ��wiy��x�\��Q���`7�R-m�I��!x�� �賞v�C/��	��<�Uh�뛇�A���U�ҕ�����d{�m�ո3���^�덊5��;H��W�k���6�G��}N@)eJ�u�g���)��� ~�K�´��5�U~r�7���|�A���ui�(�����K�������I[]�n߿z׾���������o�h��߷����������_�/�����_�����}��W�/~������~���������]���׾��ߵ������7_������:��đ8�dme�s,_K�1�{��PG���E�ꀷ�r���\:�X�� ����O�;K#��f�G%O*����*K|"�����S�����V�;��^1M�+�k� �J/��-�6xe�W�`d�=�=|�������  ���8a�n��j��+�|ptM�ׯ1�_��w���Ɩ+�6�����vx���
�Ǘ�o���υ9�K�4��m�Ơ���� T���p9qu �eh�Et�>K�S.����mT��1���s�]焣S\�ť�ӳOB7����Pނ����o��
?8|�/xQ>u���\y���7�w�Woll�����C����̹z��7�{��F{��EZ�j��-��)�B�x�˹r$�.y��W�_�/�������O/q���|9��d z�C`:M��o>U�AO)ϤTm	��gW�sD������SI/ 6�D�AUc@��eC�i*-S�~m��)=��y����K�maq�MLI7�x�2Rzѭ=�Bn�P.�,�� HD|[�*�>C��hٲ3�V;A^��v��mg�����Ņ΍�`ʮ:LK'6������!��;�ɉ˖��SéCIO�㳻c����WTT� �&4����%�������g���=>="'��}�2?#������J<�yh�� �����ÇqW�o�߯�ϵ{�}'�i�^��߾�����&�|�����xG�Kg���n�@x92�f�/�̆��Fo5k��*\�!�����G��7�͹�xX?G�i�H��r	��(c�ɒ���2&�}�r��޾���Ն#-� �x�P*�u�N��H5�G�VKU�*̥��FeEL=.Q*��V=���c��v�?�iG�8���7�\��������3~AX�v�H�<�ß:�4}�s��>*n.xȀ�btBU���
�*נ�Z�)(�Fz�� ���V��Dpi/�p�寜(�Te��O΄~Br�P��X�и�wJ�ri`Ce�f	U��|,�Q�r��_�o d\�W�Q�Щ�7NGO��'؛)��2:G$��MgL�̝��f��B���;k+�J�m`���K��;�;t�F�>�z�>�Au�� &��&�ly*E�qzCN��ӏ�G����b�N���8�6 �oe�2�i15"�HB�#!����T��8� P~L/�Y�OL��4�vu̇)OW�+�;y>^&P�r2O�|��ƵG��G�Y����y9�ų����2�iM� ��'Tu	���]Z��<KO�|=���n:GһB�a{h����+}̳ϧꞢt唗��N(W$j���7n������pت��H��ŅÞ�k{�	6`�R1f�Kt�t�t�j�+F��r}vn��E��>��� Ĩ~�G�e��_�������������ߴ?~�-�����n>���{�}@qn8#����t0
֛𸝄-Ŷ��6����54^�r�C*G�B�a��a�T=�e�G�qj+��������/�u����/��qmY+\�Ax0��Ňy����=D�������'�Q���h�ޛ^Z�u���^��ӧ��Q�Ѳ1�غ����a{�a�{�}��j�������N��v���S���c��bg]�݀l���)�8񬑜��6�a����A�Ҧ#l����QdyB�#�/JV!j���;����K��^��*T��1�.�E'���0�S�|����	�X��y����}�N�A�FXQno�+���w��3��0(G�8��՝0�j(.1�gfgg���۝;CZ�܏�o5O��AR,�`a��	�9{w{+N���z�����{׾ǡ�c�Ç5�ҡ��Oy���F- ���`��M�r�a������U�a��O'��U;%]��.���Ξ�����@C�4l����O輣�iꏮ������w�s2��[秗'ι׈��Ơ�q�I�Ot�mx��I���c�������v���3�u	\i���q6ۛ��mee�mn��ce����$e���s���+��!|���7�2j��P�����G8
avr|�V?l o�k_"����e;��Sp���"���	��N�\�^��4��O7���Z��e����w���>��{t&��=�62����[�e!�~�7GLػ��q"wkxl90���NW5�,t�ٖ��ٚi�%偅���U��u��B=�^\?���'m���ҙ�t�Gو�@������5\p�%���2:꼕�6;_���n��p�%:��R6[%�k$X��Ka"	Ma��+����~ O�>n�x�>p�Y>��� ��w���F[��4�
�㙧.D1@S����r#Z�i`�O�@R��9k�ݜ�C�i��;��\1f�G
�������=J�8��&�)�li�b%�0.���,�X�i�~_��U��pV���o�z�Q�hSً�s���)�
֜�	�.��OVĘ�t�>���D��"�t]Т�E�P,��/�T�)E"ê���,kװ��q�a�������tЙz��a)�B��O\�U�T�Ywأ�!�xO:rr��W�A�%m���n��⑎dd���v��<��nރ�3�i�X׸�G��d�A����8'g*HǴ[;�]T`�2!=���	�n���~!��t��Q��=8�W��U6�p�pXOJu��-��ӣ����)|Lb*�]��Iz��H7*���8|�+�^�i2!
e�B�0Q6!���{4:��i ]!��I���ԇ�"������Uߦ0�z/�x��B�6�(\�N6�X/i�^t�e��=m�$�[�u[�v��z�3���T
�1�I�r�+?�R�C5bT\�b}xok�۶�>FE�^NU7q��� �Ň2P�����Ƿ��_\'P�]+�.��~ŗ�g�>��W�g�1I��G��Pe���,��a62�ak���F�o�GG�0�6�(ăݽv�<�?ωo������01���=��R������a�4�����vA�����/��o�V�i�(�f�]Uu��Q���a�w�g��&U�©;|]Qn��OF�>��z�k�9��'��^\�����*.��Y�u��#F=JG	/+�Wn�1	���\$�a�z��+lz�#�zd���0i�ԯo��������~��mc(/q0Du�ћ.�9	����A�B�8sֻ䒍y6�ڠ�ӯ|2��U��rJ7�'���TT$�$�Jf��J�%^��s��qˊ4>�j��E��)�Y����sE?i�tMK
͉���Ū �6tMYl��Po�n�3��ߐcY�By��T�S�e����\����D:6j@:GN�^]�Z'��yԏ7��ki,�MC\��������LH/��7O�a94޽�v�i}�u����E.p0����x^�[���ġ�eu��	�Z�����,��c��(N��0r�tlD����aЉ�ђ�O��i�[��i��Ma3�iϟ}�~�$IC@�n�Ỵ����z��3x��F��!{����Η�tn�6��҆pȝv�Ę󠔏C8�C�@��Xm��/�㰾ko�}���)�Ii�j5��w�q���A����v���v�9�y�y��ZG���O������՗ߴ�������E�8x��(Xؠ�ba�4��id��]�ys:ͺ�Il��7�E/�i(3����pdtN1B��:/�9x�m�C�����OK����Y�0F��sf�5����<��4SqL>�+�7���Z�]�F7�bi�c�T���%�S/p���P�8����r�&Dp����<6��P��H�]Y��}W�\�GT��������/V7v�U�lz��f\���mm�:�W�:�!��c�����J�, B�n_����(]�a��g�~Ҟ?����ٕ��iƵ�a�}����w�7������X�EX���F�x5�Bj	j @�	�:'k{W'��`0��N��e$���M���)�܏��BdnS��@|��9Y�)��d9��=��!�`!' �"��e3A[HPq��d��L�/Չ��,X�Dr �.�"«�]���|^��iL'�4TD:;q�"0:�N�wN^��N�%.�	+-k���L*�	C�c>=(�1�[���V9����W��-��5�k"�+a�)Hlvj��)`ht���V pٕ�ɶ.R1�3� ��F�P��8��:�6v�1�-9DA'K��w�,�F�-m[�2'k"Ck4�zC7 ��]����}��DX���¹�j���Bg:Y8^*nC$>���)�p|b�DX$��\�W�Bu�bY^P�γ�z����|3���˺�ꉤ=p��ڢw!�v��n$e����CDˮ|qN]�����8���S�9��k�u-� �����\��`)�T������5�䇲W��`/Y�У~s�yh)=�qЊ�im��I�'���F�L��E��C��A$�J��O��0G�+|��/w����1�#M�8�����9�4�j��J�4r xa��xMa��ė]��2�5�:���t%��={�p�ڡ�F�����\	�cx�)S��K�ko�έe��P�I��rd�5�\�R��s�UvA
�D�P:?��̜���t��ߣk�1�e'!�:����#|XG@�H��'c���J�}���cI���]�Ϭ��#�ܿ����w�Mx����(�!*��4�=��u�.��P${O��Gqr��� 	q���8k�d8o{�mlb �k��su�=��.���c��=��v߱~T�F�K(\z��'e�Q�N��A�-�F��`F<���])1x�h-�y�����Ёu�i����rP�Lx�)�h?
+�D嶺�{�t2WG4AkɷGd�B&���P���O�B~�4C���*��<�;n�#,.�E�(�l,:8��
]�&qġ��[饝��*Ŵ=|^�\|~�gUV��ſ[��t���1/{	6���p�]I��H�B�\�p"K���W�V7LL���r�W�������0�u��*����#]��{��Ֆ������:�BJ��)�����Q����"���p*>=9��8�>��Q{����
�����U[��o߽^i�� �������ꢼ$i �0��SæmT���8/�wʬ=�z�s����^� }�����ߵ/�z���W���3��X;��؋�Șml�u�y�n��|�Ҿ��U����S�7�,y���;�ǽwp�����6���M��߿�aڿ��{��$MV����R�֨$w"]�	NV�0��C�	��~Bg����ʂr_D)IcRS霒[އ��Ǐ�P\�H0~���)���?�4n(�A1��yR�L<L+m�1F�8�N�Ձ��~���e�����1(R�d����)U�f��[~y��aO��4������5��8S���qv!��+l|Wp�W�����i[;N.+"�_����ZVvyk�QӴ:��h���_ �Uܥ�I�I�*�)X��D8�9a�铏��~�y{����hG}rv��	������K���_�x��o-�Nː�R�h�@�H$?e��O��>̱cOV��Ӷ�Ԏ$i���CF��^{V�fX�)Z/�D����B$ԅAb�څ��'KcP�.�2�R'F3�C�w
���U0ֲΘ�8C%���pC`{��@�k���1��. з��Äd�2��L@q���:��$.�.
�2(@���Tx+�u�B��AZ�-����:� X%!!��(A�����c'���A���"���`�2O{�g�"���;TС�1&�S���0�8Y#(y�f�<����@�ͭc���C�Ƕ"iD�x؊f���dzN��(��_PH��N�%B<C��d���i�7�GИ�1p6���p�g�?N��d�Åf�4BL��x�{�$�`it$�Ƙ�N'��:"���PH��u�~��:Xn 8�L�6��v�LyC�)n8�P��
%�X����jy����)s�Ҙq�1�eC���Ө�Y�{�PWJ�:Y���3��d��+眤~�iy���Ic��r)���*��<]�VZ��"pL�]���w���J���J�>�5���H�O؈*߉�ß��.��t���U�����`��5���AZ�1���,��9�fE}��VpP�2y�B�rx�6iȗ�]���l�1�N0F�+�$r]�RW�م8���r5pʒ�aM�g���`��	�4��am�~_�SjșC�g�D���6�򋓕�����x^�Mi�kj������G������wU�Ks,�(�RSǟ�0�ٳO֦����@s8YнE!2��C�^"[��8��j(:|� �Yl��s�0,d�pS7���6&.;wpԶ5���3�cӍ�wt����}�����3�
{���A]��+�rYtq���Q�����ټ+���1r��cѪ�)�w�9���芒EE��eg��+p��#�}��rf�+�����D����;�y˹J�)��c�S��r9���_�5(E�� �rߎ44��q��@��KP���p��t�4B��<��R�jE���W�u�~U��9:�Vu�G7���:X��vHֶ��8H�\ҹ���v�??��݀��)q��q7`��ψ��əȅ�=�t�LBY<���k�QV9-ꑠD�4~����2��������{��9K5r��3���]�<Nt��h��meu�}�ݛ��oۛ��`�2E,�h��AK�@˱a	%�K�A�5l������u���n����ͷ����o�ە�mum=��8\�q���՛���˷���^����)��e�����ն��a�� Y��먽��޾}߾���o�_���~����ng'岧J����Βy!2���;�\]�Dm��j �է�ՋEd�ڠm�;�׃�8�ޤË�E\�������VB��N��K���>�A5�9'W�@ʭ~o� �4������p[;L�]�6�y���]�ިBֻ����Hʅب�ԉj�y5�d9�T�h���K�|nח�]��J�#����R�A�6�1����8Y�BƝ�5,�b�aK�v�ݫNHe��'��Z����+ �`+�I���� ���$
 �����M{��k���o_��w�ݛ��f�Dh߿��w`�I��6�ҝ��A2�&���!�b{�mn��D�LP"�0��V���$�p�L;�z����3)�h��+��!B�õ�\*�;�8\O`g�.��#dw�Q��#�$�_Th����(T�(N��\- �14����Sq���Jx�J>j(��U���U2���d��"�vfI�KTRj�bA��(�c��G~�P�'��!&�w���ft��i���q)b0�ÏNtz�"���.�F���;F�jy~���"[��,�8���U�2���:��/�v������˶�u��6Q>nR}�n�;�mo'J�Z�Jg�S�E�\�Ѣ.�Ӥ=��KϨ4gv	�FqX�p* ��P׋�穑u�4����^8GI^Q��g{�3Q<�r�%�!��Y��Z!Mj�A�C�!�EtN��8e!�es�F�F:�b�^N^^��[l�s�
aC1�@<���G�\g��zC�B=7��}�B���f�_�Gu���Eq��h��2nP�儭�e��^�M]�QMz&�{�S��R�@J��C�UD~/t�d��5�!���������
q�*�e<L��%`�:���J(Z�˽�=�M}�x�CU�$��PT�G�䛢��%N��$u����,��gWL��1����L��������&�9��#��y7���_�u�a�Q��p�
��r��,i�ߍ����4u4-L$3�u9#�k�SW,Sz����U��p����a��|i���~�ga㊽�6h�i���Gg�B2UW�7��4��"y��-��"��%xm�����(�ټ�}�����X�8_�w5�h+h&m{��oW0�^#w��*�N!:���?�;W���vN@�N��C��돡,L�un�n��x8�j��`\o���a���y[]?���[8X�m�x��M8�d�=6l;J��C<��3>2�̀w�4��nv��I�&22�ڢ}a/�88���������F��2�κF1ur�`�����!�c����%:@���MΎб!�4��p\y-+2�>)�5x�\\g���1��,ϥ#�����S=�}�㪤o���k�W�8+�x:�C�7���:F�F�������N�8b.g�MpN�[���\ϳ�zg{��&���ǚ���^���A���Cw����ct���H;BqA�ĉ6<}��_���u5�NN�z�U\����=%5|��y�U|���#�����6��w����A{�c<��C�0p��:�����)�A �&{�u����:J��S�mjf�4\�e��_�i_�kDx��=v�a��[�H��.��E�3mxP>X�����ܧ����n5N���Ǫ���o��������ŃN�׺y��՛�[!����W+|�}��N�����\m�`����������M9X�
�N���xՑU���@9��\�gn%���Q9�\��ϱ���ay��0I�G��H��wل�N��-=�a��$}�'�6З���9����ӛ���JOWæ��ӤSU��6�6SBl���VG�;m��{��> �ٔXz?�6�;�J�)�T��|/���+g�W=G�D`k�u�O�GF,9��>q��+8N�-g	���4l�s�G�����vqz B��'�?�m!}g��J+���m��d*�J7� �KZ�� �t�^
�E��]eBĵX��0��>��Q{��>2���x��~����ΫW߷��u �\�{ia�=�������L�ތ� p��4g낍L�k>�C�\��@'��@w�'W(���!�����z��PPtX�	����-"Z�X��=00d��E�Wc(�j>���ڴU4A8��=B(���ٚ�r���9�uxL�O����N�ecP�_�+ϬBw�	,s�b� ��x��i!#��9����x/cس�5��Ғ8�t��	m��YL��R���P��B�V<�5��A{�\ahan1CG�O+eg\U����Τl=xG�$xw��E6��>�6 vx�ʺZ�N�[�u*Ӻ#Qt�̈́C�0\b����J��=P���U��x )x>:|;FZ�+$�S��a�'�A�Xv�~8J/H�Q�&
�>N�|���P�8��^����U�p|gg�0�M�KpO"2h)i�gjn�,O�f��6B�|V!-H���8C8�6d^�JX���U�g�
=r�Ғ7"\6`�Р�e`8/��ҁt����|ÿ*���*Y���T����9�N��(r�z9Y]!�_���Ǧ]�o+w���p�{x�yҴ�>螥l����45
m��� r�+h�,�^u/�0�.'����@����DP�r�tRJ�_�� ��`���[�M��q��N���U�����*&�&��#�K�(#,3�HM��%�#�\@AE�(Gp�'��id�v�����ٕ��)��6��\����H �<��B����?�Ịoj�^�H�7�\T�j��¸�C Ma�ool���o0�>@37� g�����B����Tl�w�����a�������b�cw���G�mxܵ��ph����~��`c|^ \G�)������ƫ��@B�&�^|&�h��PT˭!WF����h��v
f%S�<�Ƀ�s:X�c�u��<Ce�o���ҝrм�9�u���fķ�d���~���r�6�1hp�'#�A�q����3�A��u췯���;p�*kkY��=�ֺ� \�}�mm�*��Ȝ5d��z�Yښ����kH��\�<�t��l���ԧq*����L��z�yX>O���8=Y���.���K8;�_����G�~��-�q�&�'��W]!�9�h�_���";|T��[������A� G�,�N��n�4��vEM��lpX���U{��^,�o?��wޓ����j	 ��Ϥ/K:�Fҫ���<��_��78H>��#�Y�e���ݥ�]�Q<8�m\8o�^?�C�b#��(�4��[c� =U[�-xoO���BK~�N9Yf��8�\��Ϣר���	m(�ɲ7+K�=7���9굸�ׁa������sūp�>�
�c˨�ã�,�S�2{a�ٳ�Η>�x�{K�؆�ӯP�V]���@]�=nT�+7%�h͐�S�~�H��g�u�v��f]��v��4���"~̃�&�{�]f띋6��7��o߬��x�{��Do��w��nq=�X`$�~�n�ѡ�:Yz�U1��X�,A���io��
>p���ۙ0fK�im�����^� ߴ������}"dt�ݺu�=|�s��F�tz���Eb��c������d���*�2A��d1D�Z�P����!Ir������?��1@Zk�Wy�$}!��,Av�-�qԼ����?�둟�� v���"���1�d9,!K��L�0J�a���1xiT+S�Ͽ�>/��3��r�nr�@i�R`C�2��V�?�:8�A����4�%��y*e`�`U��=~zz��C���lnKy�ޡ(���*KK8YWY�U�G�e('��ɢlap[�x��\[�����p��v\�R�g++���v\�!�'�u�Xؤ'$�PRW1
7[��x �`��h�P�/=tN�����?�PZ���Z����Ca˝B��.��yΐiq�J��)pKY�sqB l��� �WO����k'k��M�g�"� �8Y]H�4��q^�,���<]��I�y&p��T�oN�C=�R����� p��>�4�H;�M��ټ9�0�5y$���b��ܫ�t>�1��r��@�v����і�R�.��˧I�Ô*���ԛ��{�"0'�>x��{�|0�?���h���iFv�`�W��0V����Y��~p���&�I?T�#n�(�KWɫ:t�,ύM�M?��aސ(��3�U����Qɻ��MH	^
ݒG���!S�C�"����	�cLZ�d�/�����O�-!�=�H�}d��:��7� 
�}�|T�wy҅�����Ht���C^�8��< ��M\iN����O������rm���(P�9��=��^�"e�&lpsI���0zܠc�
����I>N��N���E��}f���kh੭��#��v����Trs�U_O񑡢�s�"1Ղ-̕�|�Jڰ��$u���ENT�G����"y�N��'A4C�����P�ǜ��0�1��N\�0@�7] �����Bk�XU(��a6wg�W���d��:ћi�fp����|΍͵�T�#��e��0e��:v��)�NM�?,#{��F��H?F���j�n���S��1
��f�3���CM1�A���(_R'�"����.NU���=��"���<�u�z����o�ᗆ�J���	-��Gm��!pw���3������ɳ{�����L��mG���7m�v�K����vM��|�2�+�l��@+6�;j��M�U\��%�4�Fq/mJ�?\��߈����`:W�N�F��o�����C.h�^G��i/[>u��ߖ�;UV�����\=4��Z�Qk��*L�(@	od5���3�'/�A��i�vw.~����\�I�>���HA���y���MR[/�a��4���C\mԗV��^Y���C��dy�\��y-��>��)��w���q�^3:YKw��$��f�w�9����.^y �z��D\�[H�����,�`_�����z^��x�xV��V��M��~H�S.��ot����Z��K�λw+mmu= Q�05Ysnz���� ��y�7���E��<3����Gwm<#u�<���s[Ő�}<�����d�>{%܄]���x~��KW�V)���7B�3��D��Qa�/� �
d���)&L5����rw8ˆ��
��u]���Pc��	rr�Al����
�|�5}!�M4o[�Lە#T]�[�Tl�ȷ�S��ʒ�����P�Y-2��A�)T��LE98&\�������\'�Q��|���_KP��:���2�
����L�Y��?"���_��Bz&bh:�9_S	�^8䜨L�E�åT�W?�-�ܼ)hH~�_��u�^7�t#�iҞm��s(^�4��Yߠ�Ҭu�v]����:NSpไ������2��:�����]p���u|�B�<?��_^�7����tp����3�{9��c��q��W�-����߽s�p����g�^�y�=��.�ů������K���yZ�4������K�T	���#�����,RB<���6�����sR�jF��	����ûp�Μ�a�����hw�CV&x6c��mힶ����N{�f��z��ެl������yԶ����1Ɯ��t�g�k�x>��l���G{NZ;�a�:�Qj��A�ʷ�1� O������	v�I�hZO����
#u��Ѳ�*�{~yT(�<��G����_�	U�F�/E��0^W��ߧ�{���K���iϻ�Vz	��Y�<�`w�L���fH�Mf��t;���NG���E�±Z�>l���+nn9W�
'�!���j���'����Z�q���KGF��1�l,C��s����Y����#�רM�uB�bx8��L)�4r�����/� M
�r����^\���u��85]�N3�]�5���e|��"���ʍ�1f��C�5����{���)u�1A���#=MЩKU����q�C���а�q��j�v�H��52��b/�7��ҷUOc�bȚN����`��n ��sY �!1��a~FK�Ҩ4 �*^f���U���klq���§�	g�'��~%�a��G����#�v�2�jo���min��Z�isScmrt�9:�����Gq�ƈ3�&��(t�t/�)��⊨��x�tR�K�mDun��d���/=܈�9��
˽�-�euX�aP����|��W�{wx�<��K��:��:�!t!=F���lx�FH��E��[	=ژ\�Z�K�=��R)k�A,���<��Wֹ�!tgi�B�����t��M3?	_w�4���N{��ɟ8qzS��ڑ�)��LOg[4�kѹ|Y���U�\���ewT�s���{�����u�����A�9h�K�&F��W|�#�9���[F����5a3�}B73�\�ɵQ!�K
`�E^\Zn�o���������,I�41�Zk:2"Rg���A,��3�]`93;�;�}�z���U�]�]"Edhu�������7kz�{y���9Ǐss3s3���R��L�ίW��"(H�
�r4�4$R�ɯ����_��8`�������W�O���Ǘ�����'��U�����%�g\Ю�6��������U�dj]=+��\?���˞`{]� W�c�H4.��Iߜz7�����5zr"��'o;mtA�!�v��̧��{�JOqm04�lL<�>=��,V+�d�#�c\�H3���d��P��r��S��<� �N�9O��v\�1�u&C5}�A����(�Dfd\��_ʷ�k��x�w��T�k�w�I�Tm��5Q��g��4�=�(�*Nn���~��/J�T���GΪ�Z낺E��,�9bL�x}�Å8�h�d�e��0��1�����R�
�bh��+��B�x��z��r���%g���tR���6Q�(�0b�K�o�|F;w]�6�n��,�V���S�vVL��pW1�hQ�ʔ �]�� ��iee������F�^�Ay:xKt��z|\7q����{��^�y����4(-q`�g$��uX*�5U9�W�0�"���g������<N����b7���[cGyco*��V�Cn>m��~����=-��篷�ӗ������������n�m`,�aDa�s}�����c�:�8=�s�4���������ȆCY��8gg��Y9F�d�\�>ęm���G�����W��TVa�z���w^�+���>x'ms���ѥ����7��L���F޹�j�4 �1�C�!;�w��ݭtY����5�����q��1�c��a�b`�gS�-���9Ɩ�m�\���>�����q1�H��4�5��R/��t#��u�j8ݳߞ=�Rg��с���IY'YBO����|�r�و�ߥoT/��9G:�y=�g0i���J��7Q0���~�����H�5�*Hɇ�����w^���{�����%�K޲U�8�y�o�Yk[������o�&��Z�23]���Q����S�mEG�+�t���=9'rf6Jl�}�"_�c8��|K�9c{%p[)镧́.O�\����O�4i$��WI6l�:��@u�x�rX/�<e}��#��뮹kd���4�[C֛zy�S�K�N\m�"�1��e�ҍ�331�f��,x1�4}�@6��)�����6
@.(����!]U��;�D���]�U	��(#�|���Fm�pҚ�î��1:���鵎�h�D3}i��H�pq�����N��Q��1;л��m���p�*����Mu�W�u�V)��M��P>�z�:o�4[<Y���q;�V�ϧo����j5�]�1�����H3��O���/6y%�>��_����r]�6��.�[�]�����'�L�)�r�x�o��R�<�2�l��U�qg���p!�HR	0�(���3�R��;��6?����n�;������Z�n�e�:J̃q�|;��DA��2�^X�)K!H�sP���v�w�(�Kxdh����+��K.�s�h�'�X�u+D�f:K�o8 $\�U�ma�@)��]�����r�N��/�3 +e��eo�F9�Q���i�h��N���n[ۛ���*u��5�R��g�^��r���l�ah۩uМ�D)��<��[z*���?���(�=y*I�H�MZ�VeP�Upn<"k"tćF��ZM�#�q�.(��H�Ο�^��_�T�1�G�W��.#�(��bQ�������wD!��p�\��?�Ϻ�uD�:ze��
�=�Cc�2MS�c1�.�#���UJu�Y㽦���Ak7��I��40�..1�4�F4���F��J�\�]�Fe0m��_Rpp���Hw7����%,�ϑ�׏
�^x��S��#U�*���j�֞@q�P�)�#�q�a�@V���]�o���2�r�89re>��4~�5�M���z֕��sd�r������W�%��E�i(��4�'�����|M]ؔC���K[�i���jl��!�UX���|LKG����7C0b#�P�I��dX!�]z#^�I���N��0r��=�_��������a{�n�={�۞��k/���w���NƠ��v9<Ӯ��17��௎Gi4�4����0x��>�3�E�Ș�r�����F��thk�:R�����Ҡu<Z��{�������Jeq����? �5�*4=`{w�����]%�	mS֍2ɩ��#F�$������Lf��!8�?��U�Qg���I{������o����C��Ѷ�7�vv����q�&8�Q��R�k�q7iڈ	��L	�E�f@��)��1N��
�V��5{�k�[�
�<��n��]T/N�w�G�;�bt���;i5�
���O�<n�t32�b������bG�}�>�&�<�͜�%R�(E)���SֲM��a]�~͜2ǚ�^�-�9=�0���wy;�:��5uk�p�/�ݺ��ܹ�hg��&xw��s�د��C��.���?Κ�[������=�"�I��l����u�A����S�ڹY���?�M��k�q�|SF�r���?��%|01i�k�3�Y9�kB��4��c�q�S�e��#�i�L�/��~�G�&_�735��V��Mr�Ҙ�4q��҃;szΜ�t����#F�5���	�8�e9I/�!vg;�N:Vu]�z�{H�Ԗ:�ʷ�|%�2���ӓ�a����YG��;�B��60k���/|�Ͱ��G�s@�V��z��g>��dCش���0ҏy�Jdz/�{��jC-G�	�^��ԻΟ�q���m�y�˥_�{b$�\�RI�{-G���o>򗎇�շ�����q�s^I��������	���g��Fǈ�~h��3�u�I��(l� ���nu��=�%�dPJ2A.H%a��D�V�'�MaP��|j�ޖ��*������۷ncd=��p��D��̆	R�\��~��nfOy;x��\�`|�F!�2�?���]��9��*��ӪP�j
�~�>SBR�)�d`Un��l���KE#p2�/�NX�2��bn�B�8��$#sen6�g�%9u�~���-�u�ٚ�P��F����?���.�a�2i�2\Mՠҹ�&i�9����������a�*Gnn�+�C��BB�7a�^~ݢŞA�h�Z�]#m���`�H/*����:]��c���M;�n���8/�a�/t�q�i+*}8RvsC�E���!� ,SZ�4�0`��_k��1��Ѭ�hB7���9�"��3:Q����2���U�,^�ޫ��2J�)��v
�i�9k(ܙͩZs0�Bw�ĥ6��5���Cc|��p�۳N��߸$帮n�_�&�D���m�4R��]+)櫟<b'OF�=�-FV���o=�@e��ef��	��j�٩L#=�2���!󈈥�Z�'.B�����ާ�A���#��)~��:j�w?�#��
�'4���:|��1�J%�6�;�{]��3{Gf4Q::7<�nu*!���6Y��0��4��%d�ʙ�Z ������mcA9\Oa�nO}vfSI&�9�_�k�΀�|h��\����ݣ˶�{�)���ap�9l�_�����h�#w�t-��!*n�;G]kt��n6���9Sd�q�rí�=(z{{%�8�v\�*P��.M�q"jo��KCw����o	�K����+/�qE���.UFwv=���o<_�Σ��lg����K'�퐇a� ���Ĉ�T;gm�C�1������Wm�j�p��cmck��F\�w���xPBҾ�}�|m�3=p�;(�|���Ƴ�-=�x�0G�(+M�W4ûГW)�(����(e� *#	�#�w��:s�4��$�nԁ0��%Zfc�I$ySE�F�����NA���|N=-��s�K���+�	q+�u���`�q��Ó�*�I������_�/p��n��Zi�Km^�C�Q-ː�w�i
��)t���=nO�<n�k�ѯz��vS�� �(\�5�e	gu�!����sSH��$��(��U#>�G4����g��ADd	,��i�I���w��mc}�{�<�g}ZG�QR�{�x��f��	��^L�J�=](��'���2An�4���12�AP�$/�GxqqE-��+�8(�>kgCNe`���T�m��uX�F։���XxF���O���'� {�
爻h���ۧ,�p��j��t���e8V9���<3�|�A�c�;��Ug2�q���;�_����~d q��I�z=���HZ]��G?r(u��=�2�OKZ��׍��[�g=��|�g�>����(.�f Ǎ2��6����X�%���ioɫD��:�!�y�;db2g��F���1���{�Y		Q�_@dj�h���-WEIL��KZw0��{wﵕ��2[� ��tU���^^�`�z�y���^W޿��T��{������<���i7J6�>�/�*ܸ�M)QVJ�d��)d�����b|�'sW3�Ϟ�s��"@�ӯ��4j0�~1�!��jh:1�bh����Bi�q��d_��ʖ�(��+���@�IGy����� ���S#U��it��*�<:+;���s�a�sW�>�T�Skʖ�����2�4Ԝ�`�T�C����� �cF7�Ш6{%=q�#xŸS!�� <�#�fjU-+{�('��F��o B��+ ��Ј�C����B�)YZ(S�Z*�*�c��̓�=�kH7B8�#����G95���hS�u���/ݒ{�m��q)�VS8��Z�T�aGh�/��4{��ޥ���t��Ы�W�>��tB�8Ӎ��[����)��S=����(kF��|�IR�i3"|Se5��tzW"�]�T�Rg���������������G�򸾀8��z��Rr���}X��9
^�Bgh��)U��Q+RY#�n�{^��t4��P�O��,���X�B+
𘍽��?�*�4���]p�B��p	o��
����8G�+�(G@s�I��]8��e�����՛����A{�|�={��^��k�>��nB�a�*�[�1��uZ�K(��Ցq9�H�[��o���:;�������/�������o�ˀV�.�<���^}<����q%)U���hϿ��"�\��"��A3!�w�.��)�����������=w��w�ĝu�/1��xnm�`�jez������+;d<3ҴA�áUtW:Ĺ�|7<�걗���:�4�t�ۮn,��s�=/� �J�Cv �4�&4����]d�M�#�� V{iz=l��V�Oc/���P��V^
��,]�ha�ؿ�:e=G�2.z�2>r��Ƴz�_��!��U�(>�g��n/�4i��A�nꥡ��矷���:w�������4�ez�<K��c��#`���K�2�2����/`�p�l���\v�����g�t
?��¥l�K��)�	!3T('0��pC�q<�1��ք]��7�6�)�M�U�%�l��|������L�5ʷ:+�^����-��N:C
#L�n��H#r ��I#f|�t�G�D����U9�K���7�݉�n�_�ӊ&y�Nm/�+��J��޺N�th�h�CV��T��$ԅ��)��dA�l���p$q�����f��v�S��X����d�p�{"F�q	W�8|�K��;�W��3��6˫��hQ*��tq�w�U�}�_ҁ^��V'Ewy�����u��o��yx/��_�n�_p�������U$*T#&0�V)���h�6�p�L
�2��.7@��S��T�B���p�7Gp�©k�4u
����v���ދ�c�u��i4�f�$
�?\���]g���J�q������/�=�{<�w�z^~�"={rh���S�*�D���^R ��.��U�ͱ�*�:�;�FLod9B�P%Z�g��4��`Ùj�R��d�x���[����{�Y��j�~��J��y��ng?|�N2+EN��F�zW�ghLAk>ǰ�����_�4&�z�� LU����\d��Y�!��w|	={��1F��=#FW>H�m��l#�5P��9*h]�W��)i�ǆ�q����L��5_��� �C��rT˵:�Q�6�n�;9=�Q�;*�9�����j$�[-��`�*�3�"G��<_#�c�1��&IK�@z�4js�7K2S88�\`��@C����!Y/�߸����M�r'���ۥ{3|�Y�����M�c�u���/�z0����1b�O8${��9�����i�n߾��!����z4ȯ�w �%m0����/��g�����k�ySq�[�
�=��4��ؘ�H��@=6�6֝��_��G�T�ª��a,id���m�UJ�.�4[�9
u���4����.�(3R�8��ʡȟ���_������Y/7������m�Vܛw�z�iP8jU�{?mM�Y��I{�/R/�޽mo޼��޷����9{0v�%櫊J�����_�߿�U1���2�vv�;�i��B��E��^qd��~�#�<4xck�}�؆��N���%��>��K�����6wlYwup\k�N1��2��:/��$�����i�Ϻ!�r���	�9�4���#RbŉMiO:&Y�����s����r^�[:��@~�ؒh�H�z�>�a���TF�iP���������I/�G���@��D�laK�)ډ�_7�i[����W�-���������Y�����$J�� @�jl}�����駟�'�����+���K�����yaa��ah�A�ky�7������",~i�-?.S�O���Ň2�ܴ�z�X]�N������w&�4�ͨ����X*�),H�1Mޝv9F�1r��1q4�z#GCK�j�|2 �ȓF�4M~I��M�6qL��4:�#h�_i�&�_��l�ҏ4��%���~��5K?��w����@hd�87Lt1t�,��-t���s�a�ߔ߸QGt'141}��/��;��O����ͮ~*m��X����{I�)K�2w��H��L(�yp�x�Ѵ��;�u�U<`}��F�.:RGW7R˯��4�өo����<�O�4��\	�=��u�ݏw�*g���I���&iE�s�i��Nx��o���^���HR������2^1d/X��B�P�Z��� ���L/�^�,w�S))¥�n �����1��`ؙTanYz�eˌ*��z�*d �k�Z���?���t	xųB���A0����c���ҩ?X#��-�ROm�Y=��T����S0�� ��{� <�@��������Qr����cۓ����{2�z��1���|T�;��S�GpRO�����!��C�� �O<Yy��lL�[8�P�a���,�
�Ð(e� �#�7a֧Ǒ��L�;-1#o�����M<4�=���c,�-�M�T�3�D�Ѡ�
CO��]�����\Ik�M꧃'�j��0�9��Y��&��e䥑�"[��`hML�bh�h<\�1�!����܈��D0�NC�*��E������1�aM�P{w���s�\���k��aI����_���f����S4��{� ��?��2 F����9&�<�k�W^�?�~��;8��j)�U|�l�~�����N��@��ƽ�-GH� y �����=��(�^�CE܄�]��e7���{5��|���Cg(�Q&m���'#c�o�GI��u�i��K���zeKJ/6J������g5`���W����5����uλ]t�ȼ�d}��0���N1�0p{]��-�����՛���m�`�W�3r�H5�l�,}P��!��4S;�������-�4gw�͈4��C\[v�.��q2 �?�*��~�o��է[�?J0��R���yG¹�_�Iq{dV��z?����?�������`��+�s�~c�������]dx�;D�����r�i�n�c�L�A�����L����lGT���EYlsP���:������|\ѓ~N2�R؋�2R�������2�aL��txu�1�-��X��'��w.J��dy (۝ ?���z�T�K�7��G��_S*��#�]w�l=/����a�'���/�ӧO�˗/1�w����r{�4�/�l�՟�i�����?��?m_~�U{��af���Tyw�SR��q4�����ق��q�����WX/�@�"�U|�q%mtm�#N1�iNk�aQH8R�;d�%�;>�*}��ް��9�˚1�V'<N���R�-}�0B�̩H��N��NGY�2�Ǹ�0�1�9{���>/��}�z��k�/��K\�{����!�|�V����'���*W���0�i�� �\	�Q��!wu��K�&�Hô��_�e��*Ak�n��墬iq7�տz���4�*�*a{��UZ^��^g�/����v�8�#�'�%-���^��]^/��ڙW�����T�t�s��l|3�^��]:Q6:z�.u��җ�����W�x��>�̨�1��0��iz��]I��K��	���dT���O��dEz �0# 0cw��%����+GB�%!{S%�^߿�n�~x��dyy�ݽw�ݻ���g��&S�g��r�s:�F��hE���`�`�m�h�m��=�@Z����)����s����5)QdI�������6a{�Bp%�@��%��O12r�	yd���z� �NiR���Lg9�;�Ni/����A'����L�)����	�0d���S��M��Yp�Ҏ�>5Ax��]���a֍FM���]Q�4��B|�]A� �(�	�[0gKq��)��M٭Ņut,
s���
L'�u�/���<�a�"x���`P̣/@33��nʞ��������/~hoi����]m���!4�l������^�iv.2������v
����w;`|�t\�葸j���
���<��Z���X���T2D�L���uw��:R����43u�2{>���
a�C�]s���l���ws�Y���6?�����$�M��,i��W#ViN���ӆ&�Z����|���f�Y�(�g،^bĹ�\gd��:k6ue�u.ui�.P�U�M���PƤ��̈�1�E�4�6:.)>����H�����ˈ��C�]����<�O�SV}��:\�j�B�6~ ��4�
��yw��n��k�(/%�e� ����v��ٱ�z���|�hJ:8�+;8�"'M�����J�rS�7l�ROOɃ����=2���R2�κùFF�3^��l5O�)�#;HK0d�K�ew#3�l~1�*�1�Q�nm8߽�����8-<A}({OΝK=��`x����=Y��"[��!�����}cAeʵ[��;�w�'z��9�sw�P7��1��;��y(tBD{�����8�<�:O�)����>y#�8q��J:G���w�w�C��_���'��ͫ���w�a\��ܧ�1MNbp��m�������6.i���aC���w��;��n�q(����ap���vL�O��`��'�R,��v6�h�(ߑ��A�׶���*�Y]�L��i�z9M:�hS����V�HdxJ:*�҃�M�<���&���?i֩��ȳ��5����N/<�A#٨T�M��;49�{n��<� ʂQ���,GX=�^]\X^���a�=�	��u�e�s:o��t P^g @Q�re8�b|��K���v���l�@���kۇ�����j�cD�o��ѱ�d�6ک�K9 })k��f�1b�i��i��;w��[�i��$y��E{��Uv�"�\�I޶����9����۹������\�h��8����"��z[\Z	^�j�a5��y����qm?�;�F�t������NGt�k@!b)�+y��g[;��tͱ��v��	�@[3�併���G�ɣ[�ed��H��p6y���C��<l������:��@f�)�9@��6��܌#�KK0H�$T��揍O�C� }����87O��l�Aۜ��9�27R�<����83���6>B�D�k�V}٩����x��&�k�(iY�*�mw��D?��m'�k��{�w�92�$�C�{`$7�i+�Ľ��lR�c䨿�vY��:M��\kӉ$3�x�]�u^�Z�߻ᕧҺ��ʬ"pmW̸�Q���A\˻9V:$�r�v�;�2�6�KU���J&x��_���<�=�e�oD��P���lC�9tZ�PF��Ó�] t�v�MtfѻV�,�0J99��?��_��؎�a��& ���1�2�-' �=.��P8�1�ɀ)��"_(��u�Q�U%]��ȅq�k���$����i�T$�7o޵�/^f]��^KK���[���b�AP�K�f#Y9��We9�ă�߿�4�����}��t�T勨�e�@W5�%4���g	��]��%s�^UY�<��,T����yp3��L���l�] �&�d��WcV�ĕ�$L	��s�Z&y�SI� 8|�h�1퍝��S�mCLa�h���\���4ŷ��P��s+��VY�T�֡�8Re�K�Qa���khē�b�ʕ��
� �|΃7Nm�壄|��1��Ν�U�:0a��ei��ۻ�iX�>{��3�y�2 �R��4bG(ȇmc�(kvQ`1��ZZ?#������6�pm�K��gmM��b�+��T���M�R+i�B�:�ӛ�덬��#D��Vi!M%	�+��a�h<�`H��3�cc�ԇ� g���n�M����GF栅9�7��e]��S�%m��dL�� O�X��\޻+��W�k�
���KX^�/ك[��^!�.�o�uS#�N'�n2��H�u��\����S�4��|F���o��g��`?
�|�7��������4Z�e��S�����E��0J���,��F��C��p���'�^6�p³��E����t�<䒼������Hr�f�%��y��?A�]<�I�q��T�|��em�k��O/��^(��F��]���G|��׵YB)�Q*�K7���Sa��a|y/��uMnؠq��$"+�Ѯ��RI�����JL�  �A�>J� 
4��p��8�R�
���%�.R�]�ԓ�1��s��V{��u{����������2��P�/ol�ͭ}��a�S�l���g��Ä�
x|���8
�R����4_`��S��#�U*[�@��
d�l��1q�3�����t:�:*9�<���{�2[R�o^�i넧�~x��2BT\�"����:�?�r�� �ЦD��{�W`�EF����$��7C�I��N�(#�ju����$S�U�mG��VM���7�w�,5ãx�.�s���l��j���L#K�N���I3�@�/r�mw2�����Y�|����� g������b�aݹs�}��'�.��;�������^�z�4,�#9d<�ybjz����
~"_g} �r���OCö�Y����K��s7�2�Oq;!�y�
u�7CA!�4d��ęvFR��{O'�i�(���y4���%��jN[[�o?���k�(a�up��?<{՞?{�i�v�؉���1�a�����C�ſ3jRǕdh��QK�I:�^�e-i(�K�BX��#׫�1-/8��YG��}��x���U�+�l�<�փ��c2��Ϻ�{��|xVގ0���KKnp��)��O|_ʤ��<'+�
�i7)Gd��#YYo��旎G���\S*mc��^��脝�6Ô�� ��Q_3G�H|���e�?�^mM���>�*��T�}���^�)O���f�S��]W:j�F�o3��Ҳǹ,wz2�g�z���c^�O����Ň��4Xx�����(�)�h6sq
�Ea�8�2�,b�*~)�*T��
�bX�`r.�=5�kh����;�,Bl�j���mks+��dw۹s�v[��ܶSH"!eҗ1����ɩ�-Wi�bd햑���p�I����<�J���1���.�h��.�{z7��xC��'�FU*���S3��p�a"��%QK�c���H�MϠ�%��y��ZX�]��3�D�d��"���l�������֯DRF�,��g�e�����͎�`d�.&P�J�9�J%�j�+_1��8nCg\�lX�M�S�#�e�(����I]ڰYƚ��x����w޷��@qy�i5v\^�A�m{���?-ee?8-��.�����H�G�i�nza�*�
/F�Ʀ�0��gV!;�Vsj6|l<��}����mx�g�ПP4BZ
��N����_�M����N�NY:��,ch�i�YC�g����|܈[e��O�V%�|P W�����u���/�}�{���O�ZQ(�~�%{;r�ȲQRɣQ�*cʩz�@�u�����o{i� <���,�ʯ�C/�I��3Ô��jL�Hø��
�Z[ �������k��`:	펺9�e�<�/r���i� �¼Г�8�} _h<a����Y�z<?_xSy��!�S���%�T~��gᕩ�^IS�>*�J��@�L�'�}����{ё��/]�=�V�)�	�ߝ�5H'YG�۵;C�9�TÌrz?���PX42P�NQ���Lw'NvEQw���&�kF-%����ڲquЧE�.|�h)��r�$.�K���*��e ��99s��
�����߶�~�^�|�>��L���l��ư��)��r#��V�χ��s�U�����B��Ҫk��P��,�P�U�b]Q+�b��T����ST�,r�V"'����Ѧ���顔��Mѐ�m��#;|��� �A�Y7vҦ�$��c��'A�T@�,��T)��_���2qҽrKg���n)�>�5��$��ܞ��.A{�'���S����8��a�0��1���d��6��]��_�}����@����Q���w���V��mom6�O1�z��IYe��<�������]��wӷ^��l�����3&0x�!����A�Uh��W��1�����"�L����t�4w4U�^���Fe$3GV����2����� �6�vּ���X�{ųN�^��ёt�)L7���7E���K/_�i�}�<���]{�EE�ׯeN�P[���t��4\/��8��6I�#P-+YS�
D�r�2Ag%3(σ|ҁD���Z�S�2�4f��˒%�G�(|��H�ɂ�
c~��#�t �ވg> µ�vd��z6E	��S�1��NC۴��3;��9�K�%�eR�Š���k�#��q��*�%W�k���O�28qV[6A!��i��~��T�X�^BZ֑�O���':�`�u��çry'�_�EB+� }�KT�WF<��Lp�������.]FVMu�h
�k1:6,J��6�O����Ň�=���|����d��S�)b��%� >�X�u��+x�C���6�4����>ʊB�
�p�pF�ک	Qa��M�������W���j[Zt�L���!�L>��C�i�]l��K[6`(�� Fw����l!��#�K��x+��5��	Pq�5P�����7~�37z��{?��)�]/_9���l�<���%�D����S(���NN�x���h��e���|ޝ�9��9��8��-z�r{����r���kʕ�%
��n�d��*��.#[�3;A�!��A�S>l�K@�)<���"4l��f%*Ϯ��a٠!z��]{��U{��=��#NO�0�F1�.����� -+�BnE�]��=���S�RD���43{���7�M$\�dc�" �w'����JD�V��QJ���"d]��e�����*?i\�1�S{��0�f�ct�\w�0z~���F�<�Tck��_�� �2������zDH�Y_r�� ����y��t�Rn}R"���;Ji�@�b)�5�� Q�:�ݍQ2z��)�H�3鬌yI�����A9Dzr.0�t�Xg�=7���b;ty��m{��{s�t��߽r^��u�u�G����Vڢ\|�� x����aR�r+�)G�%�iL(k8F����1��r����r&a��b�>���?�V��J���ݻp<��paܒ�5�
G>*�� �7��5��1�j4� Cc�g�;�P��NjGԃ�S�
8�w�i:��h�-h4��ɻ�,��K�G�作�(?]y���Q��c�"G�;mc�=F���������k?��J���#�h�p;nX�w���{��nv��iu�gm�{g`�)�G*�ֻ��}:q��m�RN�1��Oeyz���LY��2�E1���s*}�'�9�Ը�bF�qD�7�ad�t�AY�AcPY�+�!~3@�8
���z��#͚��,�j�CuҚq��_��Q���SɁ*[S��y��{�[��BÁ-���6�=����>�:���8 F� �>�����Ж�fJw���=��#��gGBmR�������ի��N��J��1xQ���r�#�LvF�:0��N��37��N?9�A��5�MU���ݫ�Y�R��.l�ô��F	�1��[?V���zQ�+��4դ�����ʃ(��<i}��t��������c�ru�~���������w�?o/_�C�;H�I����܃�K��v���9�: �����չ�j;�ᡄs�GF�O�l���@R��O�`�	��O��U��FV��ޅDr�]�����'���d>�Z6�s�27�:N�&�D�J�2W����綫nQo=��d��M�P�A��y$$|�������W���ؑ�N�� l53E�{�	���2��ָ�$xPv����l��l�҅�*[��+Wᯞ�{՗�Q�D�0]_��»6~n~��/,��������l[]Y�h��,��'����֮;�ۚ���i���fޡ�	R+0UMݹ�K����k��tN�+L2̊�8�Q��gff�-,��*(B=�;�і _[]m���)n���� �F�LC�QEb�j�Ȫ�?r@�F��F�!^a!"�g�u�P��S�Tw�*�*\�����]Y׿�XOT!��R����`��&�X�W�B`Q>1��Z�i�LC�S pG�Q�nD����5��LUSS�`�%��i{1f��tz��R��mqe��h���k�q|�ɡ�0�r6��3eS���@�ꗦ�)�,ˑ�����vp�����:0f�������v{�a��}�!�kNQ�Z�Ww8�ưJx3�79��c�_Aw�ٴNd.�0c�x���v��
82�QJ�j&_��V��z��!�A�����kZ�g\�$9�X�F�zO��2x�a)8��Y��C�ӫ������3�jG�b�+0g���&p҄�5�R����yƫ�	�|1�.?)`3�ĝ�lhG���Ҧg?��ɩ����F����%��V�T��b^1�eő^K�#6i��~Ҷ��;�V���*0�^�̆
ڭ��HVa
Y���|�{�'a��?W�X5���$�c�ާd���F�&a�!���/ezJ*����z�Jㄷ:Z�
]�0�A�a��a*ݼ'^ŏ�E)��#�-�pT\�wS2Ŀ�'O���[��+��(��y�G���#��CœL�r�R�^��)3��r�Ur��*�tV�L��dO�֕9r��h@�U	,3o��nX�.=K�������޶�?���}���~׾��Xis3Bw�xNYF(��Q���a��d�(�P��;{��)��+���p�;�_d����}u������W{h�����T�(��_��2yi��EB��}�~����81��]��NM���*e;8�͹���АpV�e�&]�3`�Nm7�3p[H�R��!r���K���V��T=�9u^�7�_}�7���k*�|"��w�#�m�$�(Av}�T}y�4�G�v��8+���#{�Q���k��|S8�m�cڍwvw�ۖ�[�����Շ�M�ӫ���۶��I;wN-i��ʽ8����t� m[:�ѵ9v�ntצоV����X��g�q'����v��+�J�QBZҌ��Y7#H��J֥�o����1��b�{�Y/|������M�����v��j��q�7e�F�a{��M���i�_�i�74L�(�$8vj����NhF%�C�#}�=F���g��U22��9.:�0��p�s�Rǖ-4>/�������q��!c�t�O�1����F>�S�g�c��	$�{ë�i��z���ܗ�-�SX�~m˨�,;�m�X6����A� �4^�h�Bz�Y���:�x��w4O�Q�{����Z�L0o�����xp	C��'�2X�_���r�{U]�M�C�u�y��:��aT~f������qya[d���[OMg	�v��pjÒs������v��m��:]0���=�\ef�u2:]�U)E{u�4��@��[�!�TE�El��)#�J�IDNu��)A����Q�ԝ����g����63喡��HxI�<$s��A�(�.�l�{XG�.蔋�3Ȟ?b�8���׏���)��ه���/e�)���㑝��@�$�0�4:D..0��E�EA���Б��ۓ�I�JN/�� Y����jz#k�g��2b�1=�U� =���@!�!5��I��O�ī��ͻL^HL07��@?pR&�mf�հ�	�K�ܳ&��"L����&����컙	�~kg�ml���ť#MӔg:����'nra���a���赳!��p���������ܣSi���iH��e4˲Y\u����Yr�C?�tPxH:ꜻ=H�d�C&F�pЄ[�R�&��?����f�r$c�J�ڒ���_@��������1��Gbu�I����]�xW��?<ɧV�-w�z�fB��v���*R4�����jܸ���U:2*5~)|�t�4f�â�0�c���ܥ[�("V&~ʟ��,l�Sǡ�y�F�ۃ�F�F�Z凾�6����-��sY�{U8x�?��_չ�{Y2M88Կ>'lg����{���(��M��{�ª?����t�:~��ԇM>�[N�R�f`�JgR���K�j*�odNb6hNgO�А�ގ4�Z�>WY׈����	rƩ>u�ώ��ɦ�RS�B�-2�R(�ZwvP�.G
��Qá�ٴ<�_�q����K<te��JN�wM�;�F~�ó��?��}��w�g/Q�qfD���O4��ݰ�u+�(�*�5b��Nq�@V��z��I������0E�4�t�]����"{)���c����u*���|Lå�s�g���*�ĻrD��$��#��{�5��+��F���o��ತ�(.Y�LY�L��2/åmLl�E�G�u|�w���x6Ւ���Z�	�=��ҧr	�d�^�P�&�O7y�>�6�������{�nqF`sg�;u��p��9?�����D����5�<���tfw�q��ݽ�_9�,){w�ƴ[�(�G��6>C�z�M�T}gJ;-��^�QA&�שN�s������PZ�6U��,t�)���a���D���O��	�a����z���.��G���ng�����(��޽�О~�}{�n�t>����4����Hg=k�'i�g��)P��e�N�K�uu����[��[q0��3����c�:�����2o?䟼x���{�*ÊC�ϓ<��LO�2��<A�H�\�
�	�!`��a�Q���1�H>#[�7�*��O�>�8)~(�VVh7Lf��D����$};Lm�]7fGT`6���l"���c�H1�*�!���Ū���_��Me��;/�#�͇�ħki��\4b���3���|[t���
��:���NegϵՕ�����?��Y�ۇ��Y��u��+1lUZ�2�� ���ˢHr� >HY���9�F�*��v~���%�=������f�]xn/�|�Y���eA�s9'���0�o�
7SB�.��<����?�,�ګ��E�h��R ncX�nT������"K�����I&�.\��1�����Hc��  +3�a7]�LbO�s匄wIHa�O�S�wH(�m�lL3�of"�H�wJ"6V����/ӛ��(%B��s�>=�
Z"����_`�S�yi��i8�^�x�);�C\�GI�F�����5����k(a�1��ux|��r�v�ak�ÅO���]X��7wq���)B���[�c	&��)F���4�p�Q��0�`uZ^�f��ާ� \d#�X�<��b~�[� ��:0���u�D�HЀ���P�]}�f�5"G0���ٺȃ��ҟ�����.\>�]��g�&M��4��ݼ��3Iu� ���#p�xP1q�Q��NN9�ꖻ��\^zf��E;���1�jͨ�_���z��C�@`X{�ԡ�(ǘD�HCc�s^��n��������<Z�.ڇ���!ge��h��A�Ұ�}:�_��K����0��O�[�`\.�%��K��)��3n���Y���>�<w���?����w����A�Q`����p�T}/��	k�r��8�Y�6!.Đ�i'���4�܍.J��?�g�T�t�+3����t��#7P���1�D8�G��% ��_�y�FiX�M��Q�wpi[��:���#O��-�w�ً��o�}�~x�T�����N;�w���$�tF��Vޡ�+ϱ>e��L>�vR��������W*�JH ֘���K�Q�J��}]��������3�O�d���_��^�4&�ю�?:6��L�wsQ�U8i�'�>IC��C����*�3�{߯N�LYqQ)��4��K1�_dI���J���I�����R)�W��n�{�,��K^��cG!%"-�Q�UQu�����
A���\��F�]��?�5�*��u{��7(��Zٙ#��y��I��/�g�}�>��ݺu;��Ȫ�����5�vZ��W�O:�(��J�U�i�s5�)�S ڕ������n�� ���d9��!�v���0ƃ�����svX:j�Kqk���fq�z�߲>�0�w�����h�"`�?�	g��QAt�Q����������'��Ź���:I����/ߴ�0��v�����'�/� GQ�؀W��Z��yߩMX��3W��*�c���	�rWJ�!!�P�7٘�td5�'�>� �#^h���F��R�4��!D��n�:K~{�W�=�3�ƭ���n4�1:%����0��(!�i�����V�oҲM��H����k���;������t�(���J�vj���8�Ԃ�V㠹�S��r��<ß�"�������K�����ϕ�r�R����X֑�H�1��Sg<���ŵ�~�3|��OD�r߃�����@X۫Y��ocd�5���?���׆J��"N ���<11��3�%*�9K:�Q�r��F�$���*��w��v��:�^z��Gih�=�6=	0��)�Ư2΍
������E�����Eod�졔kd�g���%
� ���սG`�u7�C㋥�����Uo����?=ӳ"#�i�hDr�D��2jt��+0
7Eإx��%$�GV+�TJ���;^�����S�NQH\�znP@��^b�.N^�|m���r⧱d�]k��y��xC:�hY��4ȜV�W8��T���zI�PO���Ը��#<&��T ���u���a�quy�v�n�:�2C�a�ꕒa���W��;�p��f�0���\��L�5OY�
|�IA���-�����������O���-�tNJorr�1 4~-xL���#��F�ʔ)7�vM7P}Ёc�� '�3��˙\�Lv�3����3��o�����$n^:�ܸ�\��A��Lq��B>(��/��B#ŵ?�
X���`B^�#ϸ�N���ℷ�P1�(���4!�ʖ���v�֝(1��btI�g��⼵mO�2�zp�]��>}��S�I�}/٠�Q8����K|�ٽux>�n�D��²(5\�Ϣ��c�2���A�����A�p�ze�
��j������D'����,㨏cˍ?����-�4��{����7J�U��t�L���͏t�}�;Ǯ�G����5�sjag|�Q�|��aw&�ǔxwjU��<$L�?��1	.�&w�"Cwj�#P�-��y��=�}����7O۷��О���Ӷrв���(
)��#V�Ϻ�n���|����o���5��J���!AyhO�GުH(�;E���&j�W���)�Q��l*�
'����vki��_�2���ʙ�J%Tyey�Q�9|G^�{/���Pw�OZ��4���,W��K{��R_�P�|�7��-�N>I�we>24��T;�OE��?qa^^������W�v&��r&Մ; b��N�|S�FI���©YZ� �2\ՍKU�-S�V�3���Gq��6��.<���ՙn߾���Ͼh�?��thR�XvJ+�4n�w���/��`�4؝Q�t�Q�3E�'v@P&q0<4E�q�~bdMz�k{G�v�q<N"��M�5��C�M�֩�f�k:��;�C��B^_b`] �7�~�KGU�c��4h*(�[��������gO�O���k�͹-���$�v�ڛ����F���j�D�e��GB�)Q�_�����r�s�\șq�p�&h͸����7p��vN����GY�����5k��dII���<�O^��/_�o��8������NQ�WmO�W>�z��w서�t�t���LAN���� ���_��֟ƕ0���5äpX<SƖ�)x������6�T�Kgda�����b�Lų̃-��.�"�B�х�ͽ`韭�z�'�-m���	
��Q؄�����ƤtgܒQ�!M ������n�v'�ce�[{���]���V�_I�5f�����d��������z,G5\�a&5�"��"YVde1�Q +��Q�D@8��&�@��J� �����O#d$�r���₨����L_b�J��cdY��m>�B�>�6�5����|�`d�[�.G#+���B&����eȃW��r�=Wj�������ܙT��K���H%S� " X�3�S5�𓰈=<T��
����K��z�$f	Ⱥ*b
8d��0u�{������"�����{��m��uG(���	B�TK�̴H��y)#� ˠ��%���*�a"D9��`�K�tQ�9����;u:��đe~������xדI�J�F�;���i��ο� �	����Oa��.4��u'F�JUz�T,:劲���Ĥ;+�{W��4<3��^;���$��'-�T����bZJ"�Wp��_ē��OЅ.�nD�fC�8a4q�A#ˑ�ж4M=tkU�#���^��I9��H_���z֛��r�K�W����J�*и+$�/���b�F�������څ4��ڰOA�f�RR�ƤI�Y�N�8):�� �f�!�д� �C�*������޽��u�-",�Y*�NUt������f;��@Y&�6��9��S��kh����T�=�I$rN�4��g�Żᕱ�e�x�������_ڑ6�^�<��p�[�d={�?�5H�0]8�a����/�|�F�w��XҜ�<�����SF�ve=�߻?ߔ'���#G={�����h{v]O��<��QL;���`6�@�|���7u��:ȼ�:���ـ�{fo 'bP�vy����o�}x��3�^aL}�-����i��[�g���7�ݻ���{��%�Զ>U,z�O΄�+˒�v/��Ǜ��5����pVQ�j��چ_!�0䔯�N�˪=���fS�!�|!���є|iu��%��x��28�c***p*��J�_ַY�<W�=JͷR�1�R�*]�C='���N��/��J��Ҝ�Vʓ��Wh�<��H�Aw���R|� ��'m�
'p���QMd��:�<:t!=d��q����I�j���_߁!=�d��  !��saa�=|��=z�����X��͛7��۷Ƚ�L!������_��>z�u�N�����t=u+�kк�}#�M/4v,�p����;
��灅vP��`�e&A`�$������1�Dv�����.6=S!k,�<�+���w��g�-��s>�ߡ�lw��y�uiB+��gȏ{�R*ހF���������>k?��gmqv��5��u�ov�v۫�2%w<�g$����a��TLϳ�(�냓ɋ:)c���n3ʦ�����Xh��䫡�L��u4�}�X)'q<y�|l��Yt䘼^Gީ�c��%5����<6�~�\��v��2�{.ڒW�
�~U#���e9�gG��sJW���[�q�@ݹ�u����Z�tHt3��z�q�e=��l��?K�C��!�c\�S�~"Sݨ��d���]*�Q^�߲&��R�mRF�dE'��	��|q7�5כN*T}7��.�az?�VuT_)��s�]���,�n�m�kGG'�ɆYw�ܤ�)��1Fֿ��=-ޓ��2�@(�fCM�P8fؕ��AZ�S*X,u��CE�pVFh*��ݩK�Ӛ?G�9�������>��I��Q������ʬV"NV�D;5>Dz��uyXɢ����1&���S&7��v���,2FFA؄�h��F"�����;z�ӫÿ�yW8��� �|�DT���%���Ȳ�S�8�ɞƪ�Q��DlE�G�@ԻB�rK����&Di����=�.�>DY����;�"|T*�����ptr��E��1���K���sz�A���_
+�X�ՕK��@��LQ�����2^z��1㚛-KF�����N��zn�Z�<pZ#���=����8w��ۭ�����ڍ�g'�;�dd6�I?�[����ۤ;�5!d���^�ld ~��zZM���:����ோbi��~t�����fU 9���ȧ�r������!�gyod�������48����a����M�w�|��T�+�4��s� @�S4( W���O�)�i�,�S�t`��մ�ť��*�ehY�6d**�tEA2%
nC��\�|��apҟtf�:!�G3-��rgdy�ʋ��Bhz�n����o�>ʌ
5�2yY^�<a�7�����	I���'��3҅yE	��y���ݽ�w$<�OC�wy%yq�F����>y�����^m�k,%.��OA*\�|]�������4]��X՟Pq�F�t]��C^i�#��4��_�P��S�Bˤ��D3\Nſ\�6m�����?�c�����ٍ�����i}[�������{�?��>`@}@Y���F��9m�ͫ�Y����ٳ��勜y��n���={�2�_�6��B4�<�6�wcd��M��6n����:2�\9�?{�Je�SL�]��)�r�w9T~�X��#�����g�%�"��%��	�A�:�3�;m�#5Vh?��)���Q2;G[?1C���/�E��d�55�7�h��}�MO����IL`��7�(��NOCy���5�m�m)�J��P�03�W��Kd�x�P,��E�S�  �k(�DCAgcv�	��kG=�V#F<ͅI0[��#|��e�Ƽ!�L����ԓo\c���c�����"��Y�,���'ݾ�9X�e$kmm-�������7�f�a���Hz�֦_ /S�ST"%�wt״{��ds2RY�M�����	p%����m08_��ᑣ4gQ���g�>l��Yz]B�<����ᙛ��jy�Qa}P�v��4��#�v�`v~.4ggZ�;��]�����[+�g?����O�>��C���O�6:��g������vx��i���hp�Q�&v�e�p�(�	~ �躄��5�4t4�=GCK�����%�/�)22wB�k�%�,�ou Hnҽ4�N�F�5�)����)wt�AQ��1�>�w�k\���ai�ͣ��7M^�=�x:>���11	�ܿ۞<~�n�Z��x|���v�ch�@ҝ:�SPm�/�m�r�vI�-�$�p�3���#��;�0����ö\���D�.�"(xו�Ui�L�|xOX]�y�z.w�*�v*rbpU"�lW�Ӟ�OJ<믱뚫���������l���7���0��*x��݌de���G���?��������6ĸ�A��a�A�,
+�iï�-��<LM#9��Y�"m Th����g6]^xV�߮���J���O�O�����Ob-&��N�K�F�<��8SMy�{����p������8n����mWm���=��Ȟ>{m���!�V$�^���(��?yz]W*_}&+��\$|9�д���<	�Tf�i���s��+�ѐu�2��#�^pL|Ó�#�e1}�#P��K��{^�B��%��ڢ�wz(F�w��)3Ntڀ#_N�?����z�uM�yrS��a�83�@-N͑��S�YVi㉩��ڨ�sa�o��x��0�"'������.�c�a(u���4�N1��.t�`v���s���5qr��w�%e�ʢX{H��@c
�L�E�Sg`|�ا�N��On�������.���H����`���40�ʠՑ�B7֧�e�U��z*Lr�ϸv,�lH�G�zHt�(tEk8����U�L�a��ǵ�za� d査4ҹN�*��p}Z���Y��9��r�<xt��PdW.u��^h�����)0��Agy���)D�JvL�n��=���(l?X6�**���=��!��nO�b�Ӟ-4q���և��ͫL��`Zy�?\����Z5���Oy�ݺ�s�_�#���y������J/#�ٲ�mç$�j��J�S����l G{!kx�eK�;LB���*��n:2b��T[��Jx��DإM0FMy� "i[F�k$ف�s!藍��T�!�.�Z{���z�(,"}��� #y���-ᆲ��[U{>���U.�r��&�wE�������eL�x���=��sϞ����z�����m{�������A��v
�� �.��g���]�.��^w���.�8�*eo�Ӂ��~l0�0��)�ȐgXz,��:�P���6f���;��e�)'l'T�3�:��0wJ���,�Y9�3��C¦C���R	�J�IH҆�z��{�c#�U�:�L���#���]���Iځ�!����a�@Yp��РS�RL��̬�:���-MJߣ8���3�.���f&���,��Ɍ2�?��p����6d#�������Jl7Gs�K�!�����JeAJw����(�����r彅��v�ν�~�6���=rktg�g��c�a�#1�T8z��h��ͯ�ӧ�b�:,��/0�?��#QZR;�D�A^R/r$�g�u��0������,��_n�>A�:��*zR�MaD/ͯ����v"k�v�����s#G��7���u�L��:�E�]��'�U�!�=�s��C�����Se��i�NP���W���y��{mw�i@}ȵ��_���>|m;��y譵3u\�9>2і�pˡWGOQ"4��V��
Z�҂t6?��x��>�w�Ecg�:s
���Ϊ��yhz�v�e�$����7tYK��K�H��oSm�+��k$i��+�T!EH@~8��}HZ�m�y	���L�s�+�95R�=:lK��㇏���>z���ww3k��e��ٓ���3�s-���C�:��Z~!��������'=Z�+�����%}�d���$R�T
ġ�{v�������q�VD��tm�;|ɣ��vA�����J��Gi�8�i��U.��Q_�s��ν�ڝ��Eg���;�3��m�:x�Ν������v�БLg)
&]S���J	� q#1��_����<[*0
E�@�v��d..��q�["�d׺�H�!וѢ��V�)��˫`������;7������w��=s�1�gݫ�}��@������˨:åg�
uc7X��ɍ$�:d���T$Ư�bV+���|��g�G(������7����3}�{��|�^�H�y��޽�l�]����ۍ��p3�����׍x��t ���! ��J�֓=j6�s�% ��\�23����r{�ff"n1_�$�`zY�R���;�ã*�ԿJ8�����]���Py��{������t�0/L`o�����P���4\��h���NU<���C+ӷ�|����'�"����s�%��s��̰���X2>�eZ�u��7�O�?�׮K�{�}� *?C߼�/ɻ�?1~3|}��x�>� �~�S*��_p��dM���,�����\+�+�ou��k�T��A���we��b\�Q�מIx�B�8�$�-?��"���?1��낊���LF��g?�W�i��xMgV���|"3�W#A7�v�t��i��q3��`X3��'��WW=$-�ƽG�W�����O�=N�J���~�-i��]ځ�w��|+����C��{��|S6��S�ʮ�w(��B7���7ߵ�������~��}�������_�M�կ����W��������/��������Qv=����r���c/��n�����tn��t����SY'��.��r�n<�M8��򤜖\S?*	ٴ���Zi(cd{��SW�_a�9
yU
s���g��͛g�!�����C���$��32D� �J�i�G#�}�u~�NE��Aa��o�Re�kx���0����3�	8q=��a�4}V1͋G���3F'��w�jz��Ʉ;9
�*k�rh����ˉ����s>�~�%|���=[*����ى�n������������}��Wل�!�\}��7�o��1���!�N�MG�m����8;^n��eDҜŖpQ���~��)k����IDW��i�v��-�S*w6��m�-�Fi����5ț����1L�:Kx�K�pƳNQq����b�qͻ���ꜙ����=�q|�4�5�(���4�xv�b��/�������;��m�C�h0f�V�h iI�6�]Cҩ�N'ՙ�g��ay�p�m�2>�'ǆ0
G�M�(*F�z7�<	���0ZP�J�#a�QW���F��NC�������?�8k�<`���W7Cgs|gM�2B�Y�]�>�	��5@�����<Q��l���llÿ�y���7�۳��'rGN��<(Z(��~�9ַ�G�]�eNq�Z�������_�=��A#_�CknD���e	����$76�i;6ڦ#���9���(�_����D����"|�p�'�����^�\�P���,�܈'#N�|vX��c�����;X�
��M��e&����:� �y��Ue��WH�Qp�w��g��w�2�p�~�¯ǋ�q�Uj����1HШ�cd��OC��f��)�Z�UO����4��Q3�jР��z�%��B�m�7�0��y��k��ڇ����S;/�1�w���������C�t��CGh����Ѝ	읲G�h"�V��ϵ�%O�.7�0kv���oZ���&U�f]e��Y�������#���v�-�b��;�ӂT����@��pd��n}rG�eJ$�۞�i�1�2�5a8uŞa�)t$����~��]52}���\F����K.i�sծ��ݟ��3x�G��MDtߒR�|�o��#~|�.�/�ūB�Q�ho�%�r�DA<^�A	��!*N��@����4�t�:���K^�쪲���jZٌ�;���7�a=�����kϠَ0��	�Vy����䝻W�����k l��I<����r�4���U���)n*�2��+�'߂�ŤOZ�g㙰�o9:8t)��K�7v��x��N�:�.]Ջ�}=G��?�7>�$=�.g�]ڹ���-�JFu΄����S!���I���GA #w���ms[�����m����0�^��j/_oƽz��^����N{�a����u��<Bfz�i���:,�Ѭ+4;�I/#�Q9�r�(��/r��Z̺*��@ed��e'\M�ꜳ�gZpF��>!�(�<�um>�[i�^p7=G.r�!�vd9��c/L��!kDiT�C�2�)�������L�h���}�3�</}���ؚ��f���S׉��so�i��a���`��]���g��,��h�8�?��0�>��9�州���r�)���D�x�Fw�LÅ���\Es���;i�g���ّ'GL����w�ݽ{�}�q��'�d��4�����7�������?<m�;��a�LuZc<`d�~Ϳ⎺��4(x�;[�g`�
���	|y�_Z�Һ�B3ⶣ���k8��P9 V��H���GM��h��}���j2�Dݔ��K���w�7���C�ֻ~���l��ӳvX���:x���\��yq����r#�(�5�$��)��s��1\�XjKW��ը��� f\�/G>�z/\fs�Fث��vz��1��.��I���H{����NZ�;�~335֖����L֙M��-C�A|�$�K�pD�ul�WX:��i�N������uhG������jV_\\j���O>m�y{���v�ޣl�07��.>_����G1�<�*S*���~�;�+��N��ru��)�:��0��NS5�-�.�s���t�
�/�1��D�(�<�:�Iv�ȻD��=���w���$��쬰~��ǹ�)�;�G]f�@{.O��d�$~�j�`���Z���N��mnvX�3�as�%V�э�?�Q^�����>�g���ŋ�fl��9>A�!� �4|V�w�s�*V1�d�^$`���0�w"�\ߢ"��X(�yK�N|������O��{w!�J��
c���y���B�P�U����. ذnY�� �]``8U��F����{f
i��UCa�dCPMN��)�H.K�%�s�����n��/��������� Ҽ�l8�{ J ��Ɗ��G�'AQ)`2��^E"\��k':����r.W�ш�1�=w���i�����,��Ų��ld�,(F:�|�8�,  D'�B��K�YHl/)�V6]��*Z��qʕ�':	��;�t�4�Lu8C�q��s`���CK�5�A��+G���uN���%��Mp8c�M���y�3��#�,�|�C�����K�q2��fS�4V��nx���IHPD]Z�T,	W��{m���������p�Ϭ���{�xֿ�^�+m��J�%<���?���8���OeR��`7#�^�1� J�#l�iG����N%�C��W��t
���J�Ѝ�9�<w(�뽫����m)�2��K>��xW�r�J��{�ښk��fӠ����/ڳ~��z���iS��_�/8Nb<w�]C�W�ED ����'��^��2,&B/O�Stx�z�*�1���x�鍡��_���q��(N�bZ�ۄ�*9T
����TyzC�2DV�$���,^׉��ۿ��;p��!I3��r��V�+�Uv��>�7~7xQ���|�cQ���\F�/T�Z�I�]+[:����	�x��i����:@��#-��+�Q6gJ$�9���܋�vx�~��L<�Evp�w�'���4����y�]��R
W��7����]��~;�j��ګ� ������	�g
bD	[6]������}d�x^����A]AC���4Ӌ�FX��-��%���o���@��pZ�r�)е��(ū����";V<7����k*c�gz��	�pDD2=��)^\Ǜ5���I�H��Ćm���˪���K����6<��V�P1_�4�4�����ߴgϞe��rQ9�����|�q���ҕO*���� �ވ�3�5%�I�����2�N�4@��Nk}rՍ<o;-�3�RYN�׃�쓞[�S�����&�"ێR�&"�b���wJ�߭�6��a�����=����]���X��a���l����ؼ��)7rm�F7q����x[X�m�+�m~��|�m�o�,�)�z�����X�sS��JXU����N���F/+ˋmaqc��w��y��xҀRo��s��Ѱ	ڼ�Z����Yj�o��{wo�;�����<F��'nw���|,��v7����Nq_]Y�fM��_�[N��N�O�3)mr昻T~�����{��(��G��F�����G!ŭu-���T�S��et13�~v�h|#�����t��,����<&�@cZ�Yt��o��_8"����8ɣk�9ŷt�»�O����7s]�u_�4]�ﮝ�K+m=@�,;e�<����Ch�����}�n{��a�s�68��n�h���/��/^�z�^���q�)�f���S��F��0(;٥M��}�:Pp��(�-�x嚆c������\v����Ĺ `��\�����i��q��#.F���A�*�i�QF��\��(ܗm����b\mo���s����b�� )T��"�0ǫ�[���W��{���Sv[��Q�z�D��(�U^�ͫ~{%0J�@2���D�xK��r9O��7�ɻ��r��ۘ_��O�Ȯ�K|h\Y����5�гAD����I�����	
2]�9�<�Aa�0�cc���:=5�����!��G9]�w@�p��v�q�,g���p�V���P��pb/#Pi(�O�#�9o�Թk��5N�1��;�i\�XW�wYS�*����h�{3�3�	�GV:������T��N����U��SIy�W_<����uwk*�� ��j����KN��^;�z�����4�І ��>��-?���5x�!e�!���^���ɿ.�7?ס��*�`,u���Z]�TF�B����J��g�%]/n�xé�T�i4[9�o�N�����R�M �@V��-X5���TW�p����}׾�����ݻ4HI��$�º#ҕv׸�oq	�����p�o��.�����I)yJ��`��'�ރ{��ǳ�7i��0Uڕ�y��2�,�tiя�_�\��r�@��{�����b��dg��ӷ`�S���&-�ﾬ\������N\]�>a��t����K<YO������s�,+��Z�u�iTu��L��\�Pe'�jd)S͋&`ĕ "���#\��L�2��)�q�o	#�ƥ,i��6L4UZ)�w�V�^�.��Kٽ'���L5�R�#3]���3�&G���4�4l�j!+U�ٲ��k��QI�/�U����ƻʙʝuc'nFb='�|���SZv�MM��50�����ҋ_��p%�t)<�|P���]��:�)��]��Ub�����&�8ů�����g�������Z����WF��T��G[J��.���9�ύV��{���|��������W�m�MCe��S���h�����Vǌ�[r�©"�S���HΤ��	����ư�-����9�C�X��cU�k�A�H�#ԙ�9]K�9kE�_�����PpwG�%�k��|���>y�)el�5z� xD��X�@Z]] 6��i�$�Qpm�G�pݜ���r�s�v{�������Çwۣ���#���z��n0��f&1^'c̭-/�|�}g���/�U�]�d�Օ�v�t?��Q���/�g�=i�o��pZ�����h��9���-�϶����ڧ�>i?�ɗ�O���g?q�q�����o{�Iw��AKĿ{{w�|� ���O�W_~�>��K��(��͢�Ўf��w-��������s,�]s͟u$�X�Z�5=X\�8��)������%]]IWY��y�A�/�ʏ�2ꭌ�Oc��2����-Ƶ�#���Ԙ�l��#_�ZKj�U���>N#MW�.l�g8`��
�uf�Ԥ��T��v,�/a䮶��լ�t�q��z{wD>�����8K���r�7���>�Ud͡����/��ݟ�u���y�~x��v�h-\y9!�����¼QLPG�����B�Eۑ��
� ��a�4�ȴc�SQrU�]ܾ���B��A����vbY^^�N��t��<�q��^�߃��xii�ݺ����Zh8`�y��ٞ����w�ڛ����Q���a���a{��}��k��*�Xʗ�1B�yg�ĠI�BV�(JkڢR�*o=#�Sf���"suq�_��C�\��FK!�����("�t�`��fA~�Ώw�gI�j~o�8IpCT���J���<yߘ~�h�_�ڊ�0�4J�ò 0C�!QE3J.��Nw�$��]��!�A�r:��BO�m=�-̴���MYC8,#�f�eF��F���ݵ,�%�Od�=(S�niH�֎^4*�ry��;
5�s$�5|�Ũ'Ώ"|���^k����{��l����!ʀg��O������ڴ�,���%WG�T$dȡ��61=�&1ǸѰ8��z��D�q}8Jj\��`�b����H����4"��^(���P+/��(	�>G2�9���Ж�5⦟��
��x�
-�띫h��7]k�*��޽����ċ0�U0h5 qu�Co(DQl��O)�e��i]���&Ǉ��1hb2��n�k'��	mo;�tҐx���%�t��;����c�訷�)?�S���*P�h�#�N_u��W?�Y��p+Vq�����������/~�޼yENaEՌ2"*fUf�I�=�g��U� 5p�NϜ�!E|�y��K՗8vږu.U�T�3ZG�>��[���F����ec�k�e���̋<{Ó�w�2?��M\��!���_���*�/y�gQ��;�ɦc ~8���G� Y�<�'����b ��c � ޴��e+z�ܨ��@J�]z��.߄M�WY�4��~2�<&�W�5q�l�H�z�i��3�w���OD	qq�P7�%ޥ�.?$՚�\Y�y�E���^<����1����h���H3m�7�І4C:=-%���2�_��s�'m�����NHO�nq_J�!] Ӕ�����ށ��W�㤥��873��֥�Vv�C�񰼬v�Q�*ez��GܔS��Km�]eQfҭ��J��I.���G�R��d6M;ԁ�uq��A���2r���rđwD=gv:�쬍B|��
�9%^ģ���&k٣n��Q�Nuw�f�8�	�Wd�F<��h���m��n:qh��W���s���L;<�ʆg���G&�14<	���"�!u��63�E�N�=Gʀezc�T�������1�)[��i�Q*���\��e�u`ҩ��5N<�Ђv��7�(c��@�:��3��t�;+s�g?�����럶�>�ظ��f�C�������/��h;;�u:ʴ���L��o�n��^1͈/��wwFw�#�]��w;���(�:|j����q���ťL)S��x���ɚ�����5�B���˸���Pi �k��-���������v͞�`e`�(�n�3وÍ��)��nj�N�o^���3&=GS��}k�=���쁰��D\ef��w���7/1��`�?�.��[oѧv(+��L���AYY�Dnp��Q�����V���k��#j==J+�񍛙��N�5���Fr����#�:��i�2^��{��G;-]ɑቒS�#�kL�a�l�)t��,w�[�S�n��E������v�ӎ��Sb���;��G�`��-�S�]�F�_�Ȃ�����T;�0W*�E�(Ced�e�sv�Y�J|�da[H
	 2��G�����;����_~ھ�=��^�{ûNgxXA��v ���^��߾F)����ѽ�ѣ���,�9,fxW��x�^F� ��>�ng=jO�﷧/���Gm�Q1�)���/=�b��QN��R�,Gj-t	��'��ĩP@���B'�Mh�+L?��������"�]�(:�d��qw�.~�>nW�*��jh� ajd)�F���۹�ed�Se�-�s3H�!,�S�)}��m,~���<��rw�V��@\b�ȶ����lF&�V��!��6;KE�X����!���itm�C����=k�v�R�v�rv��,�$�l��)u���?���w�0��lf�D1�=^*�ZN������V��S7��a�615��1�Fa�+���(��Q��p7�l���*]���Ti��w����m���u�O�;qg�M���@*$���+E�7�����ԍ{�y^�8��LE�x'�gR(~�v^���{e�:4��x��S�˕BT��F����c�d�ny�Kq`oϤ�#N����܎)hS�<9ޣ��n[�[1��#+ u��U�9�2�.��r�x3\�ߩ4� ���N�(n����'O�����Obd�,�QWV���c�,���ܶ�4cP�4�f)-�%���g�{��2��y���'�p�ow�o���R�������O��$3�Q�3]{5��_�%�44�aĩЈ?�L� �^~��ß����^~�Y6rB~wJ����]yzg$� �+��z����+߭�"�x+Hťt��1c˛�#͊gL5��������\�v�7.aKR����Ti۰�c�q�u����O����e��q=:z#�(^Bj8�C�7��
�������;!�[ꢫ�j�;�U~�|�lؤ�_��� >�� :(��������)_��'W���aC�(U=�����Ӻm^��\E{��>?�w�*9%�W�+`-���Q:�ݲ��,��G�S3�p(Z��z��;v$c��<�Rxh��;ιk`9e������L�]�����.�W�q7FwJ�`���m��qQE�Mw<��z�#�2r�Qv˔�&�|p����ʹk��b��ԑUQ6��jD�#k~��it%��c�Y;	�zG�#3l�&��F(��� ��iS5��'i+�Y��L��]��<��g�HB��!'���#�F��3N�wɂ�(��N��3������ۧ��o��|�~����٧1>����347޿k[���Nٛ����uD6�s�:-��
����g�i���7X����)�/uGs��7#8Nw�N�[�8ګc�h���ꨐ��%/ʯ�f�L��S��m�%	�wch�����&�C������d�鴞uv��X����o;Ur��z1�)t:�y��(���oS�_֕3�hk�7��wI�>g�}����?���(��	_P!�_�ᴣ�І�8�&��<C|zNV�;�wu��-���Ҩm�9�C]��H�Pg�.ț�q�Ç6�4ҥw�	�r)��BHW�v�5;킳~��i�� I0��L!I�iK��ʻkf�A�'f�P;����$�mu=xy��Y�7F�N|��}{�&���<2��qGX�����-.s�ӭ����p�Xn"�˻J���֬�����}��� oC �t�j8ĿCe��w��C����tA�L��,�e�]Q��+��@�[s驟L!�?�t���Ӷ��u� ��cdXp5m
���L��?�~\�J;��Յ���}�{]�a$�z��N�_��&�I7=�6Z�+j�/|�Z&%|Ot��-�]�*�
#�����k�ɆQg�&c��;4Ous�a�.⡿nx�&S^���d��Q�aMF�,
i��L�j�B�嶠�S����s�E�����)�kj�e�^����v��vxp�P���jt�]l��y�
�n%ﰸSJ���16:#+nbCC���"�e�
�N�E��9,����R.�럾z�'V��3��o��Ɉ�8��z(5��Գ9�����w�r��s�K~�$r�>�NpU���.L�/��5W9�%���#�U��W����4-|��kѣ2,�Oy�s�z��봜#t�W�7 ƴ���Y��D���<N= �v<�U<Rq4Z�󋛳,��fz���md\��yI{����@=S|�&�{�X呺�^ ��7�I���TXc�C/���<�ʧ~���6`��a�JSe"Yqy��,�E!.Ϣ�7y�V�K�]��^L�2o",�	�+Ʀ��k�U��_x�{���R�M?.A�c7������p;��p��#���̳����Ʃ e������(;	�y5���<�^�z��K�L�v�N�RV�p�~��;�S"D*X��#)P����Ea�qEG��A��˂K��6?o�$�ş��Q�Ы��R�����|��IG?��-�64cT�e=�u\�'�|�ē�4�t_�S(����i��U>��q���� 5��+!���^�� ��L�Buz�����xҳ�H�w��jȇ��/�&�&7����ty�k�l���$kE��G��+�dvD�J�24�&�=�]�3�a�6�ۣ����������!�H�3L�.�2�\#&�Y���aƋ+�Nё��D*�����M�ܰ�d���`�wM���F��L=X�%�K��Ļy���R�hk��bE�aݐ*i�F��4��+L�:<�;ީu��#��U�@'ԁ�e���J���r�¥�N^k���.1��xfv�o�m�2�M�����4J4ǒ#9HΘo3��rf��|[Z^h+n�W�:�o���*�|sf�*���`�.��z��U��:���Y��w�ޭԫg0�VVWR���1�5�Gǭ���&�/��wV��{�������x����j|��/:��t;e�8F���r&��ȗk�t��mN��_��Y���xG���<fZ�N49i>�U�њ����I�����oS�|��F��ML௑�R��^83��(e'��]Ù#F0�n0�KN���� ��	�[xQ~t���3k�0�W� t�'�NN(ץi]m�#ܺZ2�����3�����\�a;�5�g���J�[��>h�<j�����kK𣆮Sx�`�i�35ꈻF��7ڻ���d� y�����ꄌ�[��$�3m�L$��9�C%F�E�?���\��p���G!�� �	��G'mk{��z��}��7�w��C{��-�d��ݻ.�P�W��K~�Q H�
�C�霌d
���i��=ˮO�K\V6�荬�n�!9�m�r�Wʫ����n
�z�e��[��p�[~!k�x�p�o�pN���-a�6����:��P��]y��K�n^sEYT�*���w�o��
7�����*�1�g����>a�,\��^O{2T�u�+�xa�i��@ѵ��(=����a�./���4�.�<w������F�a\����+V�x�Ѓ�a��4
a�	}t�鈝�E�.^���YN��������.�w�HC����EIY����t�C�(M\�R^�����C��FO�
�����/W�?�Y��7�.��ԗ|��Dr<	T��%?���2ͮ׊_B��tN��V��S#�S��V�^�Zd��T����&�W��W���u�oj�_�U@��\��d#�D���������iu
���tly�f��1˟�잓����i]��O��ϳ>�+�$�~E#�\�����+�$H޽2u���O�q�W}����/P�1�rWnW��)x2Z�3��+<
OM�"A��DyJ���_5�2˃[��'D��y3�w��q�iY��R'?��/��9Gy�i�ȢZ�c�B{�=0��xi��wϽ_�����W���r6�\jCʭ�n}PW���K$�~�%�>t�g�_��VrFA���t��+t@|�H<�^�+�*\��7���)?�=0��pyλaBbN߽���L�J��KT�@;��6��'F��'�IzWɗ�{���{E�8����='դ_��QQpm����)�	�C�?5�X?r�>x�Y�sy�6�W<��е��hT�	�҆!����Vd�|b8��!Y���>���v��������F;N��:e���I�N9eۛ�����(��b}{�]��Z$��;f��D�Ri#�Q�R�-;���A�S�h\�x�f��n��q���P6��qA�q�X7�ig{��ۺpʜ���c��p�q��F��g�/qַ���N)_C|��n�Ri�8���U���e����wÌb��Am����e����4a�5��1��;�}zf�ͺtb�)�v�bH�^9�3���IWҏ�I��A�mġ-�~=��z ���O�C7��q�r;�/����9��<����ؙ��Ø~�DTpV�r���=Z�?�H:��sT��B?v�Q����+m	�5Xas�kaa)nye���i�k��ާ0@4��29�!2O��9Ϙ�&�g���*��Ḋ[ɳk�&1�4�zy�Ƞq�xb��z�z��DiZZ-� �����Z�N�W�X�k����&&1
1�&1�4u����Q���B��5��w��:w�WV׳f�Fͭi���)�	  ��IDATL��� ��g�ÿ��+����1�Pp���Bj�J�F�?���D��,�f������Hs��Qa
�L��"����.�޽ݖB�{{mg�!�W���߶o��}����p�4|�޽�+~m}�-�k�X�r)V;�@��0wt��}2\F���<��y��V��$Df�@ˏe��ս�B�%x����l�ޯJjy�u����/r���:� �K9���[�����g��`Jp}S���.�
�� %��Q����J�A�:wN�	7���c��Y�x��Y�j��F�(8�������ҵ3��h`��$[� ưGL�Z�!6rvZ'���J!}y9-^`d����Q;��:=Q��d|��:"=o�@~%hۛ���0�[��LG�+�l�s����"n,���P���~u�#�o�?��A�w))wn1�(���'ϩ.>枰����o��wWh���k~�ʻ��h.���<n$���;C��L
���2\�%��ˊӅ!�kZ4A�xG$-�jh�kR)9W��~��L���
V�2�4�2%�3myû�̦�!uu��D^�e�tn���z��򳼲BC3p��;z6M�K�*�ֽI�̲W.*?��?��/5�#`�{�j��t����>�/�᧌��/Tz�kPa�oy���I?W�/����Z���;�R;M�^D��0�|sz�0!��˨Vw�F��~t��Ge�>/�1��~����/��~��M�|Vy���.�3_� ���J��4|��p_���0�����Ye�߅��C��'-�8���iE��,��]��ܓR�XTi*AC��ܠ#^���:�&4�.�WC�<&e>]��7��x{�*���o�4^�%j#�H�����8=�(d�條�M6�\E�"~�EE�����!��� ����[OwɌ��o;T��w��$
�:�&cT������A{��'��3	�K^�'pj9z$N�ė툺��1�Y��ˋ(��/�?o���ߴ�����5������Q�gG�7 @�>���y�p?<��}�;A�q��5�Nks��[�{wGH����BYG��v�Y.��h�@C�޶=x�#Xe����t���N�R�pI�g�#�9X��b`�cB���J.
����j����Μ���9>>�f1�n�G9��2�5l�K$7�q�0 �C1���;{�ر۳�N�^��^hG�3&T��d�2/�	C`q���5p�!�5:nc��Ņ�N�"K��
�����1��#���
c��9��4Fn�."�.�9e^1����C�ɍ�N�m�]Kw䎟����FQe,�����D1���E����H�0;,��.�A�;u޵FC�Xkk�r��F���h\i e��D�JC�{����53����C�];VF���J�p�K��:���64��0��;7Gv�cSv4 ���Ю�i���h�u;g@��z�t�NH�Q�W��uƔ�$�����9��s}�$F��y1,Wo�i��}iy}]�YP]�puH\ �j+�q~&=�2������kY<d{�@�������a}�j�Gƞ7��I���,I�:�ŗo$����f�Q�m�^�� ��z+�M`�ĝ�ͭ��o���mm춹�嶾fo��R|�����6��,$o�%��:v�ֺ�r�?k[;�B�������q���b��.RL!��@�Rϟ���Ռ���!�
���"�I 8���s}Ux{��G�t�¯ �`�0��1����������Y(�M�ll���`����#O��&�,R �@�)�����z|Jݝ��#��:*���6N�N���v��c}������8��h�U;��6���Ãd�X��^�|�e��H�>,*���F����i�&0�hZ"L��Is�����)�|�A�6����4���z|��L̶ቹ�!��|�n���ێ���P`Y?�κ�9�һP9�Y�SDԏ�
�7-�w��H����k�j��xI���u���ƨ{��K��#����а��<gD��?N�S�]>q^u�xJ]�-NO�HQU��Lm����e�_�s���?9C8;�}�NhH���&S>�U��o]AU���b�=�Nŭ�3q붿�����6��p����:��o�5�O:٘��F�f��V���O�ֆQmn>+�Ҡ_֪	�饀5�-XU�J1�q�Q�ş�sQ����F���UڻnO��F�h��4eCp=�^̠��_$Qs�sϓ;u�]����縲��͞|�{`��iٛm+x�~���:��a�,��?J�����aDs�f(ah'���)^	l��DY�h�*,� �#c����2�9Lv�(Kó�K'���BiQ~ʁ�[[GyIݩ ���F�#`"/ 'w�Խ�j���2�m��)	RF��|�*Ul���t7d�
�g��-s��%e�\ߓ*��N�&*����N�~��miHz��Tz�O*i�D��>�.�;Ҷ7��y���N�x�K���9�'��ԕ0Q7֕pRje�� =�Px݀�j���4�O�]��0�ܜN��ҫ;F���u��pdW>��!��)�=���݁�[��3��f#���%�� �%�I������� ��yg�#��2K�KC+�
�r�"��{�4j�mS��s��N_��4NYa�#�1����n¢⨑���NOVQt���{�޿{���5�[mg��*�G٬�/׼��̷Ut�ed���\����Y�,�.�A�:hQ���,��0��z�Vf&�ܥ{�
BU��F6�)�\�XS9��z�`�'G_,�9T'_�Zm�����X�ּZ��8S%2�:�o�~� m��H�$0LO�Q/�-�`�!���h;:n��0{Gn�^�Nۇͣ���n{�j��|�:�md�a{�r���߶7O�UH�q<F�3�{k;���8i�q��?��˝����ޥ��������~A�GGnr�^��j/^l�7ov1���;j�?�c����m;�\Gmg� �ھ��}ʲ�y�>��m���w�}�ў?}�^>����=����ƅ�,^��ׄ��]{��]{�n�mf:�?�\��쀍�p;En�y7�<�y4G��?:n{��
���Oa�mנ�G�0�=��#ä1���t�f���D�45�]�;;{)���v��B'N,څPh�N0��v\o&��e��^�E��ص���=�����3i�q#苎�-.�a�-�1h��v�|;C��@���K�0d�;��Ɩ�d�,=�nv�sk��}��mo�oe��a֋_d=��8��9����_\��_����o�6!L���+{o%X�!�E=?7��]ܫ��Y���K-��$�f4Y�`Ȩ� �_\6��z{}�}�ɓ����h�|��a䞶�����߷_��ߵ_���������=�������/�|�=�����FA"��H?*��8p�6�����Q�`�}�l�={3A�[�SE�ե�HE�������
P�Q�m?��+�Ў7��A�_���`�{]��=V�<�w6nCE��_Dè3�B���<�w�lxl��ԃ����~��(���tX�A!���g��K�֨����;��x�9J�?³��@��Ɂt�g8��Q*;�,;g|��@�oS�����6e<j3��Z[jw﮷��Y�O��.����[�M�����l�(����>n��b���؋�|��y�j#����b��2��C�i8T2z��0� ��9�v�΅N!�L��.j�n��F�@���.w�=ਜ
2�o��#��h ��uYF �b���F���1"O[ʒ��,��nży��w��34,����%�rſ�ҫ��Ŀ�Sy����+%�YWW�Ћ�=.��&����u7K"���w(
�mwycpd:���b�"���:e���A��~dyEɂ�b� �
��7�m��7y��W�M?��gȚ/��Og#����_�_��l�W�i�^�D�ٯE���5���Ȭ��l}id���ha-�L�w4�]x����]Q�'���W_�E��«�7�xOGXG#^�e�q?r�l���TȈ|�� �Ft��*b�yow/
��a썷<�l萻����FF�T�䓔��:�i]��R�u��b(�|�C�m��9�ho�F���9���rm�0�J�0Jz��H�o�
Wr����ر�(��;��Nie���g�K2��K�iv�v�l�N�N�0�]�F�mw�. `@�*[���7�ŰλƎ|[��t2��"�巌
���:�X	�U��-���+�)_: ȯ����L��.��B_���"��I�w��D��E�9~�9�̙�����+d/�����^��R�v8���q�����4j��g�`o0HN������[#��s�J�80/G(�[�\;�$rOew[��C�5�n�#�1�9Y�̓�6>��;~�������,7���r��W_���?�G���;(����o��˿l�߿O��G>)�J]Q�֣���<��}���IC�կ~��������O����y���D�fy����|;��̹?��(�v�Q�a{��ؙ*���sN�ՖVֳ���[mw��xn"h���Lv�t<O (�R���� 2}H�$���C�Sc�K�t�����4R�ǆ�"��
����l�{o-�fݺ��3�A���kV�����q��3;kЭ��1����H9g�Z���ui���Ñ���FK�#��Ÿ�/�Ƙ�u'�I�=y�Q6!q�BeG�`���n�.��v����D��Yc���z-;�\Fa8�[8�q��1e��1��4��层�2@/���w���K�Ӱx?:���ʳ�Ņ���T�1�?;F,��Ce���0*,�k�R"G:��fYz�S�1F���G�`���`�p�mb�3���Θ�U ��K��	0�n����Z��Y:0��6׎��0���v�P@޸���_\�(Jl:����K8*G�g�j-� ����D��F�to�hY��g�ݵ��ȣn�:� �O������˫��߷���Y{���s�0�X����X:�2i��?9
uF�1��s5��D#K� a�$_��@B�P�sa��b��v��ӏcd�Z_��W�t5��������_����^�(B���?m�}�F��nM�ֵ���C0��c����7F��X������#kb?D�\�Iĥ�BHcg�S&]�0?w}�����+eX�_B�&N�K�
�Gn��:�LR����j���فA��5�m��f�!04��x�='�#��?��p�XWF�bX�PEH
��*h	��N�! ����@J�:��1�@`�u��,{��0��i昛ǠmSc
P��A�=�.r�n-�������\z-�N����}x��}x��mn}�Xޅi�T������''<�x�̷���i�����ًms�p�q��p��4D�.9$<22���1{)��#�LW�m�Q�����2k�;�f�k*�︆h$��Tš�uT�C�^�qod�?f����
��+�A�g��L��"?����F��7$��s���ĺ���>^��u��� ~�f�Jѫ��ywβ�A>��(�<�3I�fldmo����{�;� �e�O����3Jш|�T\�M�8�^x�w�[Ӌ�����t�P���۞ݱ��Ծ����K�+y�)�*�O�~�~��?O��e�{T�4�A\(�E��O�鋡~8Q���r�Uufݡ���ed�+?�x�~�����ec�� �8������_��MyӇ��, ��˝�&'����rU�mhyZ�Fͼ�z��ЃPwww###��H TB8�FGr�]Yb�n�1����g;f�Y���,
����Ju])��l�#�Ux,�����4h���dʵ$���0�-GI���H�o���Ȳ\��g����GKD�O�o�:�'|�_#�
Pi�����'��,�t^�w�D
[x��M��o�U0�6�4}���C�.�P�e �}4�^1^i����Ż��*.��<�C��2�-7� }2ç�� ��w�β&�������p������ﵩA��({��z(�n8�|T��TŉayN;D�*C��e�$��G(����o*TYS�+:|�.~�Y�M9�1V��A���H�p�Đm��Ҍ��b`�È���5;����v�������Y{p�~��)~O�>�9f�	kop�?�S��G������(������S�n/_�M�.��3p�zC��-,#74����6�s�D���4nT���ǉ63�ؖ�o��r;w����-�m���;�u�����Vѝ8�,^;*6偑�cd��h�92o�Jk5�ڒ���0��ڬ�����y��Z[����4M�:�պ���j�ҥ��MYp>+w#�����ͧ�I�5�2]��Zdk7M��[F]�E��` )��7e�F�k��'�5�2�HOZ��G�"Ҝ�d���OBU|Y�a�10)�D�z����=:/�:ER*�)���,����P���2�hcuy90�;�G�X�2��A�ǰҸ�����v�uT�%Y��cB8"�����i�ē�,�ޮ�p��5M;�=�`v��c�v�\���F���S����>��є&��YϹ����B���X���Y�O$|��Ä�w��<��6+2MـSV�D����������j_}����+�G����0﷡����?ad�#�9F�v�=��0�N�1�H�,FA8:v��H�1�<�HB�3�$�!��?�JY6t+���z��<�2V�G��G��tKǇ��gh��տo�2�Yw����|�>��S���ݕ��<B�2�������<�#Y�;���#Yed�v$�$F�=6n�ݏd] kz���r��[g6o��J?�QY%��˻e�@�Oc�_$^� ǨG6\Z�$�*��f�R��7�!dG�0<Ψ@G�N5��:���4�.Ҙ#<�ꍫr*�Z�y�D�)�46�9��^�/u�a1;�&;�PaQ�l����gi���F�̤sS�*��mn��z��W������[�ޭUf�����\}��C_�����>妁4w���P z��~��ԇ1����-u��}�ڃ���P׍�ݦ�T�v#�e4k��*��� O���ž�
�&�5�w/� �w\Q�Զ3N
��c��R쌬(г�et�ϡ�vT��a�{�HO��/i�3�� L^H�x��ݥM��Y~�#Y�����������p�R��F�	����w��,G7�f5�T�54��ף���mon��=���2��Ȃht7�,�+]��+(21�"NU|y�J�. @e���V�A����O����eA�k�<s�/~����?�O������}�1q�ҋ�`)I?�%.#�9���I�I��0���]�C�˺��:�F�����k��<��J�E��q�nQ�֢ xLB/}��}�؀���F}H����Ҫq��]��f!�[od�_�(߼}o�Kc�Y2����W������x�aC�UHJ���;�De�����;w�^��#1��p����4�I��5�r��4i��6�6�S1�Y���IG'��B<��K�r�T�4��׏JON��!M^Ґ���ftF<��ߍ�l�����s4 _��h�#l�M �4m�	�=��*_( �/ͯ���_�ˇ���U'[m�-�+2� �?}�ճE^�A��'FG{�����X�&L*�*�^}Z�oZ��[�Zv�^���q�I�Ê�L��[�sE�ƻ���#ܥX�/��Y�r��Y�P9
>�(tk��_ڗ�~���r]�R�F7+�N��pE�Y�mu�#G�ܺ�Ό��K���jSSc�<���ɱ2��*8�jd��wG��D�=��kdM�..�|�Ѥ�,$��EeN>�9^^�U��$������t9�иc�k�/�h�����]hWB���1ʫʳ|'�1z1���uA{h�i�E�$��n��Ȋ)���n+���2�:+5pP��! *��P�wm����O�bq&e�>H�7�}XI���C�f�Kck�����?���GM����6;?_�F���h������Ӏ�mc�o��ƨ&oq�ugԋ��tX�I��/��2o;��O424����:�Or>�['� ��'=Fz�t����Tyu�2��=V�:�h�G ��K8�آ��p�']�*����\ʓsp%���F|�_�"+Ȳ(g������3����C\e �4M��s��t�(����C&:��m����
G���(p�v�i�n�b����a}�^� ��Z���9��i��C)Z6��U�x��mΩ���W��v4��X��HV�:����H�*;�M�C�g�M;�"�<��].?}����?�I�����ۗ�<hWǛ��n���?����HFJ�F��4�OB�Xy���։�����k$��!���B�PQ*�
�pMo��`]]YðZ�)�k++���J�w��,���u�����.�O�/���5]p�A{�H#��-�;Kmu����Ù���Ȣ� � ���}���0�����,��n��y?]�B#K,�J����p�*b�����-�4�Rl�杴���_�r��8��v><F��V��W͉2��><N5��Ⱥ��v��*Q#����ͅQ�]�	B��)6���B��8�#AI\~/!���gc�8ai�z#W�eB�T������<C�g(�m
�76|B���9F�y��m��K���{���{���[cXY �!k��?�~�^�~��c��:�+�h�G8��@����i�;��՛����71��m��#�Q��ˉ�nz�s�݁�ؑ�a{�\�(Ө(� �PV=e�� ɕQ�����R�J�ideT������4"�Q�af�$.w�I�V�Ɨ���]z�t�?��^t�c=k��0�qM?u�����U�HZy��%߇������+��)�|Iy2�Țls3
��Ȳ���m�m;4�{{�M��Q�R~�ЊqmF�bd����7�$s�i���# T�ʘ=����>����g?k����]����ݛ�W���Y�7ݶ߾E��9�1N�2�+�u�Uh{���-�!��u-ųgOQ��u
�
v��B�N���H@�q'�4RIsa�^��S���O�|;��������W�j����yRm,S�j�-g�PN��=�O<��+�����Zz�̯oLTZ}���̖����(N����?m[��L>�XI���Up�5*#^*;�u�����}���)�p9���.�)Z6����lo�{��kl�C*:ȧ*�2�*��,K��0qp����P��g���h��s�3�E}[+��N����]%Oe��J���hKO:�nM#�2�P ?�c��_����k���rҙ�\D���'�^���v��`��x��������@}x�Iҡ���WST��^YN>u�1{�5��o�mnn�����/?��rc q���K��q3��m�m��%>���x�S3�U�TrTZ5�,�#��=�81��C[�^���h�.��KC�TH��{�6tw;��߼~��K���,�Z������2#�I'kU�qQ��]>���H���.�E'bd�]Zt��3��G����۷o��9�!�j�:9:>
�ϡ;S�{�{#_'�y`��W���o?����L���4�hA�8��ƹ��c�����Q,��S�02(�$�Z87X��Z]����3mkg�mP�Җӷ��%*3��Վ"��1�C*#mH�;r�B�ď���O�͎��i�gG=	��/yR_;;�G��(�n40FQO�ɭ\wv�u�!��(�eqx����?���ҍ<+�젰-�����Վ�^NE/ ��`m�3�[md�K���\��\�[9����9��H�L{֣��7��G5�k�g������<�z�&0I+���%ϙ�q<�W��8�Sk��TZ-^(XI�gyO�vic�(�b9���Q��29*l�c��G��,Ҙ�x:���u�<�\u���3vJ���V�>bg� �F�ĻF�Ɨ�H��uy�&����Ì �������:��N��J�C_Og��?�\�������I���ß���?���9����p�����/j��m'_H� �0>H,*w�Nt�/�i���XSQVxz�B<-uY i`�(-z�R(Dp��g���{wrx��'&��%Ij���m�?:<&�4�q��R▐�z�(6�ƒ�� 8{A�?�1-���L�.��OE_f�#nݎ��40�h�B��%�_�˫�N��_�wUB>�9W���/?���0�p��T0�w6\ρ3�  �#:�;f�)~�Afyd`��0��ޒf��;�7&"�g���T"���nM�) QF0Vj���#i���|�.ңi���W���g�
���1؀ź0�!��g�����
h���Uc�C3up|�l�����s��$�����C��#4���IƳ�0�28�:�]�|e$���w�}U��{����DsрL��;��8�����P(0�����N�_�_�#��a�4-M�L:���U��{�yUZ7?X�*ݤ�[�ܿ��3.~�{}|�.��Q��iD
h{��U�� n�O(�m(�(�8�鵁��W��Yȥ\�H^U���M]ʃ�@��RIX[[o���F;���X)�%�$|G�N�}i���Y.�*�0
/��F��m��O��?)c�����[�zE�獟�
7�W�	����}��g���?�� d��=��h��(O�E�w�t���������(�kQ���<z�͆ٻu���ѩq��T���+�U���Ic�s�Hg�O��l�5:�����I�<Zӂ-��;U��F8����K�n�\q���\Ca��vΪ">�XӉ�L��!Q�.,W^?vE��Z�~�[�F1
'ևr���B%~������}������r��]���$�V)�P�S��J[��yὤ�����>�8똿���/�(�����@++���7RxH�'��Ǐ�Ym�bZ
���g(���w��j�*��~㬕�/���}��'I�5ԟ�q���s���}����l�}�=y���yL�?j���#ܧ�|��E���~�_�f�aL�ɝh����{����4"�|��~f�|D^���p�z��#O�u$�Q
2���Q)ͦ![G�Zj������������.�<ks�����7�\��h�r~�ɵ������r=Ոm��]��ȅ4�s�K����B���"4�r6�Ƈ��'O;j쨭S�\c㈲�k{v�v�}sk3S}w�N@3�U��N;ʻF��]8�Fm{)�d�E.:�����д=�*ol���2$R�VJk�{^=��c¦������4�W�+7R�_e։��6�!��ͳ��?/�j3��zrj��wZ�����s�:Թ�9�,�]N��;¢������Ⲃ,-��c��n��S%ů[�_D�1m�����v�:Z��av����wu�������d��5Z��a���!�F�F�X��e:eJ����/�`�\v4���t`\��>��e��P�-x1|�,ՙ_��uL���R߂C35�$Q�ťv:�Ô2z8����?E�B���'���R^U瑻z>��M~p桬���Ъ�v��	0h@� ���2W�Zz�lև����gj�<gk�����Q|i�x�C�1��-/.���%������_�z���ox�'3�L.�s: ��XȬ�,Z��P�ӛ�E,5�d�<�d���vĉ��J�n��y���9�ݔ�
��]����B���8�&�H�q����5ųV�B�hb�d��kX`�����F�)N#�ww���-�{#�ћ.,����g{~&>���>�7���A�=���8�	���. ��ޙ  l1�����s�&B"[�CL�ՙ~z[|7ip�_�M�*rJOX���Sx^�ĝ��m��O�~S�
c�)�7�2FV�F֥��Ĥ��0{>�n�8s�@�,�T=�Ɯa�se��r��5Q��ջ��1��2JӉ �1` ¹IA�+�g�����X�L��gFmăw�)<�8w��M��/:������������L����5-�/���t�t��w.i�g�7���p	ׇ��]���s�w��C��o��Kᯄ`�
����'S�0<�J7����B\�$J�X?�pRʧX��/��	��J0G�d����ԗ'����� ����(��Q����:���7�����۷��`S~��=k5Z\0�H�SGn�kD|��io�#o1ؔq5W�FGP�����V0-{Msjѝ�wbtx֎���x����A)�&~p���k��{~��}��1(�^wrj���Ý�\�y�w/w����|C���E�c���
�#"*���ũ���<����#đ�>j��TE{��4�#��i�e荗��T��U2L��D���iP�J�oGǇ|W��ϝbV��=/�'/��MŸ��:��v�J�W9g�,��f?��ӯ�4Ck}m�G�۹����J�<��H"�V�Q�>Ao��2���u��?�H��/1��P�ݲ\�07K�bd����x`�'���!r<���8==~;/0��+ʩ���^ه�����j�}�$Ӄwc�yV���~�Ϲm�k�],�ʷ;�^{��]�~��K�����r�����jF?q>&Ku�۷V���_~�	4�qרG;N��mh���e,��)�y�It��R���v7��v��J��۟���v��b��<:����ll!np�U%;dD4!��u"��ÐO���:�ΰ|*�KK��Ҋ|L�S�2�#�v �w�SvH_�a:�����v�{2�w��9:�a ]����=t��0I�v���(u�Z�e����E���N?�	ڴh1���b�ql;���2��f"�C��Wn���{'G�/��8��H_d�b��ɉ0�O����e, N-��Q�tF�O��VX[9l;����y'c���O~��.���t��@������И������3L�1�S��^�Yw}��o�c��·N|����W�����R�C+��i� �4h� $/GZ���w|�]����~�OC&������/��/N	cw�ݲgs5��h8>hXil�ͺ�G�C��y�Xq4T�Oö6�pj����k�F�š�W�b�J1������Zi�I��y���蔖M�p�>��:۳N�zu���N�c�L=�h���I��j���<lG��8���B�A�'���?����/^���Ȃ)�1�Pp{#ˊK:�(A+��k�0�Ȅs]��TXS!�Տd��@��iO�ʈ�V��Ѳ��<)sM�F����PB���tfr����}y�n�c��j�B�C�Yn�yp0��:<q$놑�m�U�E�=��$]���g����Sf�󮇕�ӧ���ߺ0n����7�gRȿu���R����U�0�7�`�P��\� �؈3A�H�إ�����3\`�XK����^g��H$��,8�^Z{���rq���zf5 ���GE����N\|{z��,i�0�(���4�<W���f���<�o��C1�v0�\�{
�hd���v��ĳ���d����Q��5JCC���/�u$R7Ћx�Iv�������_��ͺ\U`.�z/��;H�~�H��ӧק���q�a+^����ş�����=]$��ܺ�?����8�=������Y����SJ�tJS{V�)���4$�$��&����M��>U�(���\��� ��#}#vJ��n������&g�<ko^���N`v8���x�tL�ڼT��b�|�ѣ�r��:����7mssEh/
J複��+�g��3My�z�iN�]�4H����������F���޽�>z��-,w�q��G��}�3a��r��k�5(�U�2��֬?��k��(����#	:�e��p�HVh$x �G����դ+��TA��+N��'�9�ȓ���ࡡ���idy���S��x�`esDT��w6$z�h�g啛<eӦNi˴ 噊"qc�\%2���FΝ;���������0�Pλ��0�fZ�wo2��uX��Kd\����u/YG�_��8��	F���Յ����=���67��Ӎh��Yck��RF'ő�#b��~�W'.x/�ؾ{���}��������O?y��4��,��9�XU�WI�cd���C�G������
�,b���^|���z�9�\��tN�������b���o?���k��G��2�ܾy�ml~h�Ч� ���?���Q�j��R��c\c h��Όc쭵��x�~����p.=�NO��q�����.�Q5j9z��v��=���*�e:�0HgWY^�467��?F�m�0�����9�5�y^XN�k�K��C��Z��K]j�q .���sD�((NK�����{Y��,���ed�X�~ζ�"�6��b��+%Q�Se��Ve\�u�5Sų�W��{��#S�(o��_i ;�o�w�
͍2�n�NG�}���@g��)Y���pyF�N}�rq����2Wu���;�9'\��઻|�����CaDؤ	�.q�+i�4��Y.�:�J#�,�a�<0��H�e`(�����$L:�`�g�|E����b�� ��W�M�j@��ah:��Q|�Rfu�
u��s�뢟eV�Ằ�!P�x��74h��t�������`$�P�	��tFE�{�B��b�aJ��^�ݎ�P�Ƙ�%������9�����;��D�HS7T���*�l��3�9iY�aK_v/#w��Z�[�����:��_��_�y�H�^�Z9���J�� �"I�ѵ����6xQ��X`J�I�U���޸l� �[# d#�N%Ɨ�D���4�C�+2���F�����7���W�Zxۓ�W�I�WGE�ds��"�Y�GG��du�-F��X*�*!�蝤l�D��)'���O�^eӅ}��ׂ�߹W��.�˳�^��O\�H���9�1��8�N/b�Xt������cf���x$bqkY-Z塑U�F1t������.aLp�D��
����Y�
Q�+�)����[s��/�L�,��z�81��Sy�X�@r�ݝc`�Oc<��ge���!}v�Ȓ�(!.�͐/#���~5*�[f�����P�7��c�S/UGQ��E�(q���)��?�	��߿p�c���uN��y�x&b��'��D������iyu�U�¾^����Ž�/i��n�
+��=d��z8�����L��ɑ6�O����T�Y��Hc�F�J$uqg�+9Y/���
���=�t�y�9�uW�q�ȭ[���Q��N|��eF���s�Ɓ�˂��b����&�$?x�=��Q���&��S[(B�V�ƥP*����GZ�˼L;=���R+�*h���C�t�ӆ667����������_|�>�������;w�����7.,�+moofTK��2f�O�[�+�P�0J���ᨁ*�<�+J<w�^��eAq����G��YG�L뜶��K��wtd�t�=h�����PAp#�9}f����7g�${�X$2�DH ��*]եZ�;wfw��]#�_���,iF�"mf��w"��-�K��\��եEj�	-3�<?��Yݷ�,�Gĉ����=$B����w,�d��9��B!?�=�3�$��X��wxX��5���e���3R�/�'�9}�-��ws8�
�
��|F��Ke�Ux����_.lO�
l�:��u������o�������=e�������� �v��8X15=I�P�fm
!}ҕ#(<ԕ�Z*�*X�6�sV�������[���(X�}�)�y��˒ܸ�`B�e��\+ ��3S�H��&�a�אs�KJH9aк>H]� `��̵�����ѣ���ö�b??7�>x������^�=�p���z��*<}�$��m�p�$�D��6�I\��RD'3��.�����.�Gg
=m:u�z��m{�['x���DZ���ߢr!���e,���]�RFс`P�����7�v�L�8����L)����R�U,R��mo��Q��e�Q�Ia��W�}�A����5�Uˮ�P�t����/:t9����!��Pw�H؇��U�K�����\PpdK���]ɣ#���|j6�K�Rq���iͰ4�,�nZޫ�aZ#�ܒ{����L���=�rf�ȃ8�uPJo"'��I;��ŹyJ=�s([�8��w�#^�Y���z��.�W?A)�ޙ��o��<گ��T�w�Yt��V)�����Iʳ�-��̷�̓<VZ�t���^�~���<�K2P���DY6�r��7`��J���s��U��w5��wռ�%�*��d�vyw��囖1� e`�G޳�b��`
�{�)����x�	��8�lW�"K�*�I3f��)��#�Uvp��{jU���/Ϝ>���'�d����������Q��/��d��y��PV�Y��KɂD��(Yh�"�Ġ�f-�*�ȿ� ���t$�v�Ւ�����h���$����J��r�>}q9�3a�����ر92gӄ�aU�d=��R�ʞ�M��&����;�(V�z%��VY31�=��'�nJH�H{x�}����7��Y;�����~t*sx�\
�	�
����jڄ4q![E��F���7�J��g�3�kJqǢ��ϼ�E$d<����A@V��c�=�ۤl��0A���D��8[%˓�r�a�T��6.�v��Z�3���o?�ի\B\3Y�1�s˥�P�s����x���Q���剒e��X�,O2�qc#���?�3�u>Իn��ԇG�o���x��G��vn7|�҇qH����a����T������}������B��G.��Tj�%��R|�/��:b��fMZ�5�f絵я�����dh(�
XKY���G�Gjv��ɎԎ�Jb�FQ���ה'��rG�Ϝ=�._����Y���#�	��}Oz��僎K���H�

H��*,���[�D�q���'���1g�\vCAO�O��S4��Q� �s��<�Dk.KǼ�`�B5o��@�̔��KUl>��s��ۥ����c�"'�"x׆y���j�����t���l'i]�'���w��6��Sk<Q������}��/�?�r8���}��	*�5���˕/��V�y���^���:ra��N�w�N @�{��q��b)�P'҆{S�9�D�(��A��k�9 �q���/�u�_q}�2�������>�l�K�܇�b���|����ݻ��u�-.8h�`H�*;��j
�m�ą3}*9��Y�8�����$�J������d�q?W	/ҳ^��)����q��R��	��Κ�ߺ�v�8��S'���s�Vq���b�x MG���{���N�^�j�#�r9���o���S�Ch�XY^oW�ڮ��C�{�&�b)�n>��}gﴓ'��6މ�Y�U��y{�H�!���g}�h$���: %wvv
�8��}��P��&^�moMD!w�����%S �l!.���LL�U%H'��3�]C�I� ��1-�e��B��d���2s�L���������]Qr��=Y΄>�@��<~�(~�qy���O���؃P�!0$�h�WH�����L����U����u��Й���#*�>�:�픒WK+Uvj)�� ؞l+�l~�Ua��>!n��X� ^��Y,�C؍(t��F���Y)z���<�X���G��J��4r��+��'M��m�i��eo�
���Ǜo�dF�0|������d�V^�*t������LZ��� �1?Ɠ4���
���&o͡�7y+
/���,��/�����9��������N9��@*���<X�釼��<�-g�?��U��S�HGFa������-q(�o8(@����̪���%ܼ�x4(��9Εp␷q�����2;�錗�x��9��sp&��`�DrX�ȸ����¿ռvƥ�ϟΉ�'�ηC㴽}���������'�ړg�ma�Nt�!��'��W�� �h��� 4��H8�K*�'�?�~��6FG��h �&�p�e'��f��`�L��C���ܳ1�@p
a�T;��87?�pP�LA<�I�V����H_��[�Q����`q�-��h�  6Ϻ����t�_����8b��`%ֳ�M���0�_�qIU�K�(��S�*�Xy�#y0���o[=
�ˈ�Ӝ9��{���4�'!$׌NBk.�d�CQN���+B��c�����q��0Tde�,H�)�0�_�)� 1LQ�6�m��M�� ��t4���m{����c�4
�t�:6N9Lcw9�0˷�~�8^�a&/�7ڋE:(L��u78���$Q���0e�Nv
���IzI�|�O��R�AtQ�2�d?�u�P���]��� �)�e3֎@��'��b���{��	�O���V�t��(=> ?��y�4e��痸��t���f�ZT˒)D�'����o٪��G��h$�>%-�;���X��Ў��e����~2^����G����a�O�\X�$�XKt��Z:�WkЇ��%}���Rr�o���ݿ���~�Sv��'��IA�9�Ճ�w���
�]�5B)��Ѧ30f�����P�.]�@|Wڹ���a� #����z[Y|�^>ܖ^>��6 ێ4FG
��r���_�s�u��,ۙ3��� q��I�p;�W��#��'iK�Ϝn�)��G�왳m��:{�B����,.����>j�֖^.��~U�3I��'\���I+=�!8�^�c�3��ϙ��O��Ǐ�(�^���G����y��/��饩u��Km�>��Ν��֭k����������/���s�ަ�t����=vTZ���<�E��%3
L�(4�U�mK+eO��/�wK1�w� #���y�;t� f�`�Qy�0���y�r����J�/r��ѣ��R��U���!y!' ޼y���!X��y��9r�������0��߼�>��;����v�$J(��
�esm��-!��7�ʱ��>V��M��U�`�u/Ħw����65������۱#sm�»�hu	e|�E���M>�����*8�v9V5yt��u��7���I�.�7ͥ��;4�y$�����붲� �2�ۄ<ܬ-�������l_���(Y߶Ǵ���U����/~�q{��K��TX���Q�Vr��˗�P�A/�.�;�/���>_�mg0��QW�~����_��CM�P�u���?��j��e�}�z[A�q��8�es��Bh3�pB�ٔ�H�iG&K���Ѝ����9�0=����ڴC@��|� �P���������gO������B�'�(X(\�'��N�{�ه|�/�ϲ]�q5���rۖ�Ll'N�m'O_hS�G�1'�u�ryI��l P�,ɲ�����l�T��Y�Dр譫��25��nH/G׿Vqݡ���>y��9~);0:;��\�u�@��	��!�}��~�z�Q<����ۆ�l�2��.�"V�=;���)�B^�O�9�d �/*��՞��>y���`���'�Oy�gx���=X�x��?q����R�N��k(�7�H��wRee��>AX�X��\ 8�*�.�/��Ea���UJk�G҂6)�O)F�K�_�ޣ4W8(�DF�"��"7��K7�_M ;@{*3����>Z��e�
��R��(u��CX=�P^�B�N�zY:����j�|x]��-�-x~��]Elb�P�Pn�!*eu �x�5�Oq�̳��
f(@�M�'�i2cƻ}=��6a��a=.�>{�D���L'm�_���6_<z�e�#�!"
���U�����KԚj������%d��4}���O�u"�Y�E��k%��:�u���,u����C3��17����8d�M� =܎�N i[h+�7�w�����,��邮ϔy� (����n��gч��2yHj�S���{|�h�e�?����&���=�~�ɂ��k4�����m�ؠ!	A����p=n�G������w�w��4{6�,�We�~�NC���;�+����{T��w�^(Z�ZdV�t�
�+�T�\�����#
0�m}sEz�-.�`��/.m�r�ut�mO
$,͕�Pφ�Q����I�g�J��8�����k-���=O��閌 �y2�tK��֍I�Q��_�㻮ɤN�+��/q4����˼��ߍ��^�n����V���}�]O?�Wn��-t,���j|�}0]�,�����/gI�������.&�&>mt$
5�������܊�
��(qxs�Q?q�yA�,U�<�u�=�/��.E�-:tG��[k)Bvی�\��s⸇h�ޘ��_��e�AJ���1%�Kb�b�w>��%FG�k�1岿�0s8�u�ٽ�{��$�v���K�'3%�vOYF{��J�#�w���E˷ny,�����zFן<N�ͷ�۶�W��4j� ������%g��0��Τ�\�=Y���m�����D>X�{�N�~�Z���Xv���
�Ϟ�Q����l[�.Gk��w$�^!g[,�K⤃��dc� �v�b�ɣ�G���ts��,�/��\/���e�ҭt��ɃB��۷sw�J�x��{�����H�*�.����E�q��}�UO�\R(�\���S.U���K���2�08Ea�y,�7k<X#�5 @����,��ӧN�+�.e�ީ�����%��@��B^�6��r������l���y�tJs���/ql�.§��_�v�}��ڗ_~Eb��hޡ螰��B����(9��2�*gv�V\��<�~�%@�)��=�KF=�^�ʥ��o��8�|��ܻ�_ͽRɇ���%OO�V�!�fX�śm���+����>����1�N\9Z��D UxW1	�I�^t��%�*�\�l���.�\Z�DA�3:�5�GJ\�1�(���:��Uj�Iaߺ/~�#����a<�O��]Y�Nk���jK��>�Y�8D�l�2�H�,�쀃J��_�+mg�A�*3�����P�����F����N�6�3�/V����@�_~!E���'C']b ��H�<'�k�����ӵ�y���"P�����0��E����͸H����rx8Y�||K�P����]bZ3�������C�J�4f�K�2����Th=�V�
{p���ǟ�@�O�c!6�l�5�6�+g�����Pu��z2>��wە�k��O�x��&Cx�uD|5;Ez���GLF��Y���|ۀo��;�����B~�'�� x�G?֧3o�r� 떾��y����'�+�b�?}���?�綗���?�o��_�{�=|���*Y��tG%+�����E�5%i��Ւ`�a���.Q���%2㑘e۟QX���%st>�����,֑#GӱMN��N��X?��%:L�H?+ي��ڕ�%��������+O!�
rmo=�7�ŉm�y
Vv�H�\��k��M������mh÷01�O�n%Cq夏�g�f�)���k]���� ����pAE�f7���򥱓�������O╏�Ҋ�$�u��[��yu&7�M\�����%~�`�{i�斍�3���[��ci�u��ō,���T��������;@f�p˨�ʖ��.�������;��`��<rϻ��7��Q�����>;���x
cFQ`|�{7^b�f�����I�݇F��-aF.�ĭi}�}�u+��E0d��K�-�J�'��_jd:��
�kk��r����ҍt%�1����Js�n�Wɪ�>��gl�yM~��.<z�Df���Zt9�x�E�*!��'��d��Egۙ�)Ќ�{��̷9����:��Qe2������=xx/K���@:4z�§����� �S��Q�>`^����^{��n������n,J�S�~�lϟ>F����y��D�z�B��RGC{�#�(Zvl9�[�����[6>ӎ<p�����0-� ��O��z����W�lл�l����Ig���W	{��'}��^x�%ɥa�Ϊ!�~�b��[�*�u:��I*4.�[F�o�9�������)��-imM�V����<��u���.���ӏ����#�
<K�V�#�D���딋2�d�H{�\N�v���NM氌�?������9!p~�EtQ��}М{�\6�*�=h�C��e��=V�Է�R�5�N{طk4��^!ۛʨ��[�vz���i�P�ϣ@�;{|J�J�v[YZiϞ<�Rt��-������D3��T��O�8q��I�~w)�~o���~��������[�V8������(���Y6��W����@��Q����e���וJ7Yʐ�϶h٬?��y��) OOTH�_,����ݼu�]��S��)4yeM��Z���(Y�
��*�&u�Ll͔ �����^1�e�2�t�����[���~F�%�gC��(�U�)�y��w7ݦ���^{�@��_�@� �{\\��o�&M����8�'=Iq|x��|�i�Sfd%ڡJ�ǲ�~)ۘh�_�/�_�����ހݾ�fT��|�m�U�ӈ�a�B@STп<��2�R(l?�xǯ~��z�~��~�TB�Q�/��'�)�;�=/�R�ec)��P�(�>cJy�g��s��e�4l��̯yx��(��_��S+&T�<yR�Sq7-Ö<�{��Rw�6�Ǵte�;����օ��J��5�B����H>�vO�4y�G�|I�=��).����3Dp�闟}'o.�N�A~ķ9Ȏ���P�(
���f���wZ2��;��ж�!V;�@�}�Ka�'�
 É��m�6,=Gn酫���~d�M.�/O^�]h��[�1*Y�3�ml�cg����_�}�=z��2�%˙��v0���J�Kx`F��L�:�.*���.�%�܈}�)5W78��8{��Y��9Cm䕑x��̴��x�c����L�FD��EshP�Й�U�,��µ�U�<_8ӡ����$���~01_�7|)Kl��k������;q�V��[�[��_�;3Oz�mܘJ����_JU1�Ҽ]��	DB�����W	"���y���a��S5���a��)��<6�AyJ���n��V�Q�r���gy�&v"4h�8k��5�K������ٺ<bA�J@�^曳X[ێ{\��cg����َu��,��p��7<ûN�z�����o���(�DwM?��'��D귻�@\%�|�1��$�I�1�S��L�X����N�4��]���i���g]ů����1����#l����@���5�X%k�}��)����^�2��W�*�5�$�>�î�m=`C��5-���D�QC)PXQPqɂ�h�����¤�)��Q�"W�V��xC���6�ó�(n.u����P�L��G��ܸ�B>(Ax5O��d�~�'�Ӂ'��~,�p�8�
�*9�n_�,��ܹ���/4ޠ��^�u��-��kٓ��у��R�Q�* �޸�������N�=]�F�C����L�oW���Y�.^��.z�����e���Y>U��A���#��@8����~�=�����1��@ݒ�<n8a�CT4T��޹KynG��f��rn�y��@�=�#�h?��2I��~�_|�~���s���S�)
�T�r�ϙ��o���}��W��S���Y��|���CA9��ԉ������do���\<0���͙���ٍk7���۝[w۝�w���(�+�/�Y.���mr���۾$S�z|��w���������\�x|�+�'����OPn�_�������o�j��m����f�SZ����\�� �{�j����Q���c�C�8S�޿֒�����=����Y��y�"x��6V�(�K¹'���*m�
S�W��Q
�)���: ��dMR0���{�6�����tۧJ�3�Q.��?'_"�6��c�4Iٖr�&���A�N���OLσY�����P�O8�;���<���Q�;������{���gO��0��NW�d{��\�|���a8'Q�=����WG"OM������G)�!��`8c&�bûSfqI��	�7.�SIQJh8*��5C: f��]��W���]�)'V�/k�މo4K�i;4^sCȤ�{�n�G�i�)GQ$M�/Ţ~�dz����qu�\2(X��'}B�d1ͫ�ȉC���9�2q߇Y�a�O{�,�E�"�V�.t
e�c��7�!�3����R���(�nS����P�S��-}K�o���x���!|,d ��4�.������?�捴��Q���^2�dA=��	�;p�A?t���>N�=�U��2��|D�u ��;ʻ�:WwxM�+��8XDZ5`��_�%���
�Ű��PUvq	X���O*z�*�rx��3Y��O�'�dec�������������4�E�dQa�}�7An�J�Q(��E�� 4�VbEP���e�!��Qr����(px����
�����G|&䲋�O&��b>r�3l���0��m��u�@�3[A��d��{��>�-`���J�:HV�u��pZ
@����(�At���9o���{}ޭ�"�d6��p	;Tj^}ׂ7s7PR�+���Q���%���������؋ibIX<c�qK̕~܆���t*o��q�Q����o2X����W~�/��8�@���<3XcmcyE%�N�\�\\t	h)YKK*]ֵoݫ`с�`9���ڇ��Y.�R�Q�{���>)���^^��<�黼�����MRr��"g�>�ݟ�̲���x�_f�����z��L��{�Ȑ����+��Vn���K�������=a|�!xn��	@���,��R�e���#�
?��Zv��|,�K!�,��qɌ'Oը����V������6n��T�:<�	��~$�̎���D�hpep�7#�H�Q,���xp���8>��5������
;*(�~T��!�M�>�n;��H�$�&����d��w���@<{x�MM�;Y^w�ް��Z��,��#|�3�`r��مkWD��ʣ��
b)~��aW sمxS)P��]�d��=/AU��zեW(k4H��^	����gf&��D��Voݾ�Y�����d?	?˭PP��٤���,M��
7�Б�0���~�)B�K�2�M�5�  ��TZ-�qaqi�^�x��j��Q���~��l���g���٥J���")��/����������^1,�"n�IǄ�:�?�0=3��8y�:u������!��ɧ��d����}�M%�.
V=��S�v>o/<��)�^�`��#�g���Y�.�}UQSV��,�mo�lgP�U$=��%��Ab�{(�?|�e�]���o�<y
�ʣ�R�}	CylS�K��}�V�7�(uQ���m��#��PXϝ?��Eɘ�2��.�ٞ������������p�B�E]�*��#N�]�9";��S�QR:{�8�vdNe�)�����z���e�u��$9�L��{C�==ҏ4∼��P���,3i��~���5��Ǐ�˴�w�}����{ЏG�_�*����FxHN�/]l��x���	��;�f�~�~�p�8� /8�p�7�{8Μ�Jj��3�Wޭ6��l���K(X�s� �%����! |]e+���^�=ئ�}�`�ԥg��n㰁a�ْ.��3�-�K-���(�v�$�YK~�c~H��'9�C�6�Y�P^���K�0��X�;�RI*�e�3��Q�I��̣De|��]��+�����H�Z}�~��V&d:|�RͮR%͹�?iG�6>�{����\)�%�x�O����/uvK�U�Q���Gf��c�����i�3확þ�����j�N�w�r���D>É�,�Y,Kg!l�*>Q���cZrdF}A���L�-3���.gmU�,�H�B���k�����4�L�X�7q1�'v�`��[��;(�L���G���'�Yy7}���t�
%������=z�(����q��;d�V��tTW��,7�)=#q&z2Xy
��z���,+��Q<�
�V���>�� �+���2�u�͌� �5�x����T���F$Wg+�.]VVJ��Z�J������p<��F����>!m1�
X˃��>�I���?���UY	{5�J���/��(����я�&�_K�����!4�gzy�	E:�h
XAf���_K���`7����K�]��P�%���n�����x\��,V�������ke��z��:\v�g�"X�Ձ(Vk�+~�Q�<�+
Vf��~��R�͋��y��#ʄz{�ɇ]xEW�z�?w�պ�}�$`,�)8��v����Ć)��vic�7�F΋��oeK섉b/EC�Ƀr�u��z�;�U�����[��w��o��w��Q�v~!_���>{���E�����̅(��G�`t���
�L���v:ָ݆L�x�x�A�*;��aU!�R[g���d��63=�Ia��}9���3��{�d֖�x�k���7��{{��	g/>~�xf���W�x��af��=�ig4�va��z�㌀h�Qy��&+��
��*ϟ?A��Ѯ�4=�8
�#ޞ|w���ٺ�J�k�|��O����U��;�&n���$�~�`�.sfE�L��捛Y:v���v�ǥ?��w��wG���dN�������[7nD)���������a��S?v���9!V�S�vV�q���̊3b���"ߤq�  >š����:���=@OX����_���"(����׿�e���O��o_A���	-n��{w������w(X?�ݿ���zX��۩� bb���/:��������.�{�l!8v���5���D�~������{!�:�X��}Z�Q��={�|ml��ό�?}\Xd�8��=DA��oQ�o�'o���y���ʕK�B58�bF%D�׏UW��ɿ��[�W���}���9�������ܷ������9��̚��g?�m�r[~i���r�d����(�Ҋ{#��/�/�w��G�v	�*�@� ����Y�B�p�r��޽�>� E�W)�!#�+�lw���೜h�9����.�i?�&����wX�:|�f�]�IQ_��f�����c�����8J�����J�E/wF�:s�l�ʈYp�i��ۦ�]�%ʙ��^}�����~N�:�ȝ�rf�Y+�#.�q�E��9�p*<��?�P�����K�a� _m�\A���:�M�\YU"��fl��,,�K+���3\�+ዦ�[���M��P�-i�������$��}�U)k�+���Ѝv3�(͕�>�_�B�fC,�e���j,���Yb�	��MzCyRꉟ�-{����P{���6�>�S]��ݞ��K�	�r+>��V��Yz����8�(]>�1���A�Rڌ�|%^�r�ʮ������!���O��R�6�<
(m���F�˾���t�hm%I�5m��2]��Ym�I"�r[�QfEN�͞^.Ͼ�t���KLk��qeN��L(o�NyŃ�G�4t3��7�d�⠄���s�3��Ç��A�������Jփ�(Y98�=/f�վ�\�
��N�-+hP��q#!��s4f�,�?�x�
֡��`�od�7��:�	s#MOV�;���a�n��:���m���J�G3Y Ĭخl]C�Z^ߗ�:�
��.;�B� >|��d:8�,������C[�O\�T�aԻ�O��=a|5�X�)N{n��f�%�{�n��1�N��J�kL!�]d�0u�?�le��:������E1a��,�w��i���@� ������R�BԒE���ۤC�[��h�<��j��rF�%���Tmnz�a8j�`�!�)���/���M�Y����v{l�h�ZvaB�����wQ�zL��������phC�W�)f�71��<���_"�Sԕ˶�i��[���e�ko�ʣ�
7��x!�aث�/�?n����Q�����%���[V��#�2��𢌜^��t�mҳ3� >� �����C�n���*8�ɛ�P�N�:�N�<� t�yw��:ꮰ����R�VW��;��J�S6�G^]����~q���ctTb�������k9$�����x%��Sa�?r,ˇ."|�=w��Iמoe����\��Q�*9.3z���(���%k��Ir�K�\�5,稽O
<.�B��b=�O�}\�_DpFN�������\�� j�]"�%�}�����ٕ:�ɋzK)�q�y$#�����oJN>��s�Q���`��w�ܷ��A	xˑ�ڠ,��V�,2t�p�JH�a�E���$��6B��~]ʄ
��cs�k��'�QX���������7훯�'�Q�k�����Wx�o:k[�N�;K?�����K��{(�����Qfo%ޚ	� *< .M�`.-��g��l����)|ۙ�����y�v�F�����km�G��}f�ߺ%I��k�͓ˎ�Cqy���o~���_�3��I.gVU��"�O�x�k	��Π:�#��/���%�΂�@H��cIyE�D�^r��
�k(��'(YK�*4������و�2hq�'B=2���N��ﵷߺ؎�M�i��竡�����/�c�Bp�/J}��˸�Qg�]~�/�F��A��m�*eE��ˡO�8�٬#�#�=?q2�.GQ��K�Mۉ�{H\&����?g���<�3���~��:��9ܼ7�po�U��{S�_���L�����G�ס�,)Y��\j��;��$�� �= _�vmG��G�K�<6��ãz�I[y��Ct��2\!�U��<"ڸ �2ͤ��Q�ʿ2�p��p�!���>҄$7�Siv6M�~�N�{嶒Y��q%݄3o
��8�_�'xĭR�p�7�U��#�Gb nx���f�~�iZL�o���SN��/~�����8}*���d��?��)����C��z�~�����J�h�3�$�et鶇��������	į��[d^����>�'-�`VyVZW����xp��\�P���*��y��ɤ�q$ʐ���|���4���,�`;ql>3��d��i�S�L^maam#ę�����s��$ <C�*ҝzT����T#�^��~3�w:ܾs�}����w�������}����tXW �L�J��>��!�Ϟ?��z̝Y�:��Ϟ�]��5|�I��Ǳ�F�=�6D�+%�B���0��r��E}�;|F����=M���$2:�1�%�v�f ���K�g���|��!�̶���m��y�9��Y��� q�� �z����$�
�:�v@���7�4����"_����Fk/�����v{��ݞ-l��/���AI�i��j�x�C��������	��v�-��2�0P�^إ�P0�م�w=��ݟ�'u��������Lǎ��V�F�Mod'_����s1������,��7ؓ~b�� !��W�O�>����3�{�ѡ�arCǗR���ϱ$_e��	�W&��
�n��iZV��Z%,��#�Jk�n�/��F+}�Rk��2��_�؁�l������)�}�O�=��f��Ēokxd�	a�D���G�ʌ`<�V�̻�f���3�,��X$&��4d���g�]�7��(�)pyהy-a�N���X��2�q087��~��ʯ�����y��(�U\��`�j��p��L,�l�L��l�vg�Y'�=EGw�2�8��{���=Q��SaOٳ�v҆5m��YЏ����ˆ���w7o���P�)�
��E��b��v�hS<�@�u��$C�߼�E�to��˗��k��\D���l���3�ŗ��������kWo��G	��]H�7:sO�s�C�Tl��zѾ������;���o���m_|�u���P���hx���IK'����(���#�7v������tig��ff�0<�[����"� Qʈ�c�8�N�F�m���1���J��������_������Kh�r�Yգ�ԩ#�ĉ#��E�:��}������_�����+�/~�v��9�	�@�*ڼu.-�\��s* �sH�|@w/��'ϟ�'/��EO.�������d�[ɡ�Z����@z9&Z�ᙩvR��g�ċ�=}Й�&�h�ꬺ��6��)�:�mrΆg�&q��sx�0��x;v�M�sawT�z��2�H;wt� a���i����U=�f�0����i� ����.*��d��G�W�V9s��3��sG����;��>:yF�t�O��R6�N�`�?�����˽�v�=��e�,җ9�E�hH���]���|p�
C���Sʖ�j������~
$gÔA�+����Q=Y��#+Y�Ȩ(�?<ǆ�F_%O�<P>(h'^�Z��L<�Ŏ�w��e�ivU�ꔁx���|Ԍa�����#�i���-���m��Ϟz��f���>�a�j~_�>����(��-?��?�B��T�������>-�uJ�!+�t"�������Ly�n�Ï��uO��O
τ�_��d���ψp��|��� �:~5-Od�4_)W��'}�}r��xi��#O������I, �Md@v�3O8�6��0��2���Qȯ����=
�ߡh}��W�;F<�Ƚ)�q�2X���^' ��
�+`����W��a��N�QH�[w�=��[���V&����N�Â�#?=�|�'i�Ê��O��`���H�� �Hf�T����Ql�P���(��0M<�V���]�B��:�	�l��|��p��l�D	#L��S�0�I;�0wa|r*�1s˾~U�\8NP�^�;�Ƀ-�Wk�jiy�-��n�u[�����m�\��լ��l��)D�Ș����������g(AI�s���ۊ�ۺ���k ���t�O-�'a��k��F�<F։@chԁД3���<��覔��*z�[��$�{�z�h�<|��9�������V��khg<E��,������b�Uv�G�]��r������%B�e/ތ�P: ��$O��̼V�����K{T�5v�D��w�o���J���2]�H�H���Y�Y�6G�MCԚ~�l��_1�q��)+�=w�e������L�p��K��=i�Y���<���\����t��{�ϙ�\Ψ2 ��6
�8S'X�ި�T�&޽�p�w��"�QN��9�%
�u��]7�Q��z,~W�:���'���1����G�7�6Q0pKQ�{�����a�U���.xdv��8�R�s?�BY�W�]>4g�=@��W'Nk3�ĉ�N�O--G���ru������p��M�G�����]9��8�R��_;c/c��}ii�������������}�ۏ�{(ɽ���ټ���B�~�v�l�����)����ę��̅�(<�b�<�#6E�[[����y��x�H����r����ז8��=����3�O?����a�t�<4L_!�A�r۠H�'��9�h���/����7������蟷��{����f���{}�S���s�\w&m-���z^^]n�P�Q�W�ۆ�74��%4���]���{כ��!����h�PzI��c'�W�Ee��Df������@,۔#���/����Uh�7G�W"�O8��5'��DљOې?�A2^� ���ܘ���5����ݎ��t�#w��LA��?��.��*/���#T�\2,�Uhm��p��Ye�TFAYJ�A#*�ڊm��7�����������?�̲?�\�X�JE>�2�ϙN�E�͖����<��{J1���$A��'�/:�#�\֙�g�@�����'�(;N���Tکx�y��Rg��_{�IG?�ҏ
X�����2�+�1��-�����7�!�4���'��qi�m S���,��.r�ni3q#O�5�t�=�*����F��})�T�d�K7ІA%<iW6�>�J��K@�՞&`wTru���Ĕ��O��B��,��	k$�	(��_�U��~ހݴ��Ζ��{��y��N,�m���d-h;QZ�Ql{�J�?�e�f�)B���� P�鬬D3h(�2�v���֟�?vf�Fu���,]p]�M�I?{FlA�;�yN����N~O���`�[�B��Vnه
߭����O�Խ�����SX��`a�M�0�h��#n0�ė|`v�b��7!`!{�ͯq� %<;i��U�@FF��h�Dpf��8y��J�M���3[��b5�Y �>�_`��m ?�~SY����cz���Y�~�d��on!!m��o��������9v�J��B��=`����SJUWnp�n��zz�`���D�h���~v��;�Ô9�W�)ŧ3��n=���_�K�n���
z|=��~J����ӊR*����|��L{����fP�e��$�B��ҶtY�3o�!�/�v�B��2a�M;l��s���(��B�f���[P��b���}PԆ��t�f-7�H^��)t�\�P�Z�� �JyOGa�
���2���'�)���(;���ȋB��9zm��P�h�'��j��j�o
>�����⡢ �U��e
�}�k7us��S�^.�̱�����'�μ8���o��w)��u�C(V�4���`P���̷E�z,�S�g}s�y��K���WU�~�-@Z
L�O�B�v���͏Jd\�UH໠��L��4��W	`uxG?�-��8rT/²}�3�.�R�&�f�שX.���ǟ�����nݺC�V���|pzf.��*Q�&�j�|S�q���Ż�<=}��ݹs�ݼu7��?���&�~�|�Di��e2#�<��ޝ!={�l{����{~�N�9�#�-�t$���:�:���Y��Ne���Z�-��&������Q�����ӧO���ٔD!F�t�h'zﴜCas���'�G]�Ɍ.5��B�{U�\�;d|ԠC�p��F�b	�]D�ZE�P`����t�z�F�I�Jh0"�ù�T$��َ��"�Qz8��s9+��Ӝ����8�Ʉ nے���਄Ey�|���H��0���IO�N���I[�ʥGW��uګ<��b^.�L����Zʌ�˗�����u�W,P�S,{�~��B?�U�T��g���I8P������.{x�m�S@��=rOx�m��fJ�	���屠\�j�I���)_�G��<bۺs��=��(%��-�]�5>�����m�'�1@{�-C��lf@��䕖� @⿸S_�!��dWS:0��6&؆G OJZ~w�q��G3��R`d7΢�!�(tЯq�]7�˻��'��C �?�1���9���R�}/~j�U�O�R?�=����TX�m�w�0q�M~/�WځK���F��/�U�-�	�$O#:ѯ2���Y�(����?̞7͡�M��!��5���F���Rkd�la�� �OYT�\��D�h�v�M �*���������>kO��8W6ڪZ&D����3yp4�!���x�v��rDKRٗ� �ps�B�*�䈮��T��8��ĸB78�r,%�����:�>~�kj�MOxZ	��tPP�.���X��ޝ��W0���ve����Z��^�G�S�݇ !�c�3�f�ʾ�&�� !��(��"F3"6�j�0�u�=S��턷	�mԙ�g�Q�0z*�h��W�u���ӱ4��R�/�q����|�f�,1�/qmc2�����1�����0Z:�A0��7;�(F�K�bό�v��?�{ �R�����6���,Yt4x��ڋe܎'�RN�����.��=W��:pd+ߠY�uG6]R�咄?5�%SCC%��CS�3�I�E���ţ��!��J�a����n�9~^���Έ;���O������e 5�W��(<�k��H	���s�ʬ[��߉[�W�4�op�v��e~��W`���mx�6��	�W�mL�[c��PM#�:�#q�[ #��pE{�OP��n���j
�+���
|�
aoFd��)�a=���+�������f�w[!�4����7�,��L�I=�	M�Az���y�.G��E���G����ۃ���e�GG��s)*��;A�v��v��Y�cIC!�G=���ֽ�ʑkis��v����2oˡ0䬕��s��h묊{�܏3N�qO���<��Ν�m�����.\n��]@��O�l�m׮_�)xf)�����"|ɋ�W���x����4Hk����>BE����y��M ,%�'��'����O{~՞<Yh?�t��b�@ۅ#O�7P�"��]� �#h'�5��u�q͞�K"��|���F
�Y�	�@X�N��\f�c�(So�P�2�w�����"i�ʉ�gϜG��Ц�ͧ��]{�=������u��/�����_�w</˦��}���J�8QȲ�E��B��D\f���(���
�}"B?�ʛJY�R�=���m�y����[�_�տh}�q�	�!�,��	/}��~�������������w�������:9��V���,�q�����-�����u���4�q7N�T��`�yj���V[Z�]�6�')�J���D;v�p���Y�Z%�[А�leu�]��?hO/�7�l]Ӟ
`�O���#h�6x�ĩv��=O�h�N�lG�GgP��)K���ŵv���v��#����j�RQ�ڗ�-�K���m�]l'��}� ��e�?.W?�"���ﷷ/]i�N����о<�l�}n�T9���<���i�ʸ�T����躵"�QLR�󊃍ug��)B�3�t���򑧸BOS�|S>�~�U/=���.��N��۝�x��q��kdy��K�3Ét
���O�j��#�bc�j�����/���� �ρ�Aچw���b�&1� �pWA<D��K�����5m�����A[L�.x��nQ>��x Q���y�ȓ�<��z	-A��`�]9��{�Y����3�~�+������үf��rTx�m�0�>�Ez-%�x�hF���'yX�ˌ�򡛼D%0�f��I?���y �ˁ���w��g�(9��0ʋt>ԋ�(�
�����v��Op&c�=��k���W;n���z:*p���vh���(y�q���k. �U���3������E���ɸv��kշXF�I�8�Y��nw���d$�x���d;���G���3�~���L��)p	��S"#��K�F��h��Z���װA����a�����A�[�o.w����c'	@A�w�r*�Q'���(�$y��/*�J�
�l����d	�v,��&�+H[�+��C���w���;/y/�E���w������ppמr7@^�����������[�V܌ ���#(J�6Z��Q�װǪ��)0)LL8��v��>|��Ax�e��������\�r���^�Wl�C{�E�"��LW^#"�5UJ��|C1�h,x�P
�Px*�D��i��
��˯׿&u�����,�t ��0���PgמǴ��;|3�n\IOz0͑]���(?��c�#P�Ը��?���I�1Ņ��6�q"���=�Π Nf��Dᚤ�c�R:�+|H��Y��#>��V���lٰ�!���#����93����D/r���zr�}Sy���#��pɗ�1\~�Ye/^�����Q�ZE�qt�x���t$z~�fyȏ�xjp��u@���v���M�4��q
=���a��"����G��?~��=����lZ
Y22�'� W��~�e��s���JޝEqt|4�E���J>=�{1b�|Ѯ�jt~uu��,5�嬺uT��V�U���B�:P���m
Q����4`��M�S�*��ԭK�$�w`(�n�C����
�9�^g���kye������v���v���v��m��g�vr����HţN"���)O�o�J�Uiw�3�(Z��}A
B�Cƥ�`yr�>t�
��O�P\��V�r��v�����F )�ŅU�����A1�����s�i�l ��"�%>"��2�!B�X_՞>_i��h7n?n�o��wQ���~��n�}�2m��I����������/�>����a�S.x���g�s�Ҙ�,��Ki?
5�H�u�^z;��@G�^�Wo҇��ϟ�l�z2������ΐ����5�Ryw�����%�.iA�?(��h�(~��M��xf]"h�9��!%�<x�=x��v�(���cr�wϑ�j��0�W�%헶⬔�Ҷi���Y��xy���Q~�)s��̠�j6ݣ�;� �Ɲ<q������ӏ?n~�Q�t�r�qF+˪�g�m%�%ګY`��n�G���Cg7��ĺ�q��ݨ[�<�g�\J�	�lR�I^��п2���3��>A�Z8@�,�[f��,���9(PGok~7ny�x�,ɘ@�q�{ ���k�7�$ ��_�!��t���!^�|�N^F�LQԺB6ę�
��: O�y7�2�q�K�e�r�ڻ?�^�I�' ��0� ��?�$���O�f�eHs�����	����,r��)�_��M�ػ�?*���{Cx��I;���]ARiu�(L9��*�o�_�ѿ��{�e�} ���HE)z�YQt��ϐ������X�ȷ2{�0!����B�3��+7��R�
�(;l;��hO^{��������` В�I��@��2����T�a��Nk)��U�\��&�I�Fn�+��=|�∛��{��p���n�˾j�CYb&�J�{�c}@蘊^��՛�@�Iz�hǑ�{�f�����|�48B�����>�f92ٚ':�Q�be���AGRs�ǰ��}XƔW�,:_b���[w���{�>��{�ud� ��L����c�ײ���`��0	1
��^ ��_e'�ʡ� �n��?�O�a�nq��!�b�0�|� ���Fi5.Î:蘎CE+e౎��I6B��[���m����*�=�����"<���x�'vh��N��A�.�y��q�q�F��;w� �,��%d
X�)K�i�C��^!Yw�m�@`��֧p�<~���	t�X�NA�)�4���4��]�2O*h�KƽU��o���^T��]N�0�S����dh
^@�R*�Z<��i�IDW��{�\��x*���D�i�r�hgN��ۼFɢܹ�Ve�<������T�S0�X3K����F`^�+�a�5ʋx#���N#�`�'~���^��P��:4pTXe��(��,oe����(X����D��t$�t��#g6�����VVi�t}W �rM�c緎8+�+Ļ�����%KY	)�-��!�S'P�.�`��N?�0;��:�i�<m_~�m�w����o��v�֭����ﾂ>���ӈ��I��w�O��k��E���������l�_��������E����۽���
J�ֲ�'��w�m���/�'����:s2u�������Xr��|-,.���%?�WuE�����.�Yφ��Wxo�{z�A�g�⋞/���-��[iK�(��ߤ3�A���%3��Lу%�w�0�d���)z�|�������?��C����׏9._��6�Ld
���H�ҭ{��Cp`CE�m�k�}̏�3�3Q9�=�?�J�Aq����/rł<��S'O�\]�E��?t�|8Qڼy
����?A\^�x�;�8�X��ON�'T���OB��v���ȿ�]F�<QN0��١��u�R��<���_d���ٞ��euP�a���b��R���?u�Aؽ�=�.������L5Ph����w��4�4|mdH?��ۏ�B�ڿ'oo�0hs'nev;���Vi�P`���5�x����L����3ēv	�|wߒ���0�t��wM�o��qv��`��n?g~ę��ք��@�Z��f�Z�7��3ƥܖ�5{�Y��粛��e��cP
F�=v#��q�x|�]#�EPe�
�~����d����<�j#_�V��2f�Lc����ŏ��Y:K�R�iՓ"�J05Z�����*�R�,��0�(^�u�G'AI�"�hZ���^�F��=ӭ̡�J��������;�������[�FaH�4{L�?t�v YR�R%Jծ)�.;�F�����|�C�_����C�i',P
��r^�\���[Ձ�hm�(���@������A'6`�ey�U�E��*)	���� �؍��7���u7��P���!�G�PzͿ7>ŵ�'��8��Щ���.0�}׭�+��$�4����I�\v�3.�ف���S�U��&�-��T���)i�K¨��0kR����F�*�:��{ap�c�s�eF�IG�*a�_�Q��3���3���+�4;O��ʔ�IaW>g$*�5#挄B�T�AX��!�<}�,�֪le���y�"UJV��:4�À�����0�e�%�Ǵ�Oe��B��WC,��6$��C�P'>�bx� �v-'a ��G�;��X�.��+��ʞG�����$nq-.	��3O*�|J�}�������xQæ %J�U�@2�`��ŃiU8���wM��e��͵�YO�<��<�י���z9��vE����/��O�?�S;��,����� ��^ޢq�.� ]��� �g#�zX��Q������Ց�����Ï>h~�A��z:�xY_{��ӥv�Σ��?�?|�u���P��oV0�kk��f�KX��[~���W(k(+/����kw�W_��r�U������������}����j_|�m�v�&4�l�3F5`�L��8�������ˉ���L�d=y�e �j�%q��q  �9��4M��rZi�IW�C�Z���+$WE����F��(n�*OĹ�Ay^��������ʊXXE#*y�[� �qɮ3��J�Ҕʏ�����ޢ��moOP�T��G����ﳤ���[��Z@����8���=�ovV��0�9?��?�ƫ��U��9�r?Ҏ��Tlq8<@��N<0cyi9
�;�w/�~��1��xށ���I�@L|0˯,'v,eJ%��4����0��܇w���v���F9=�J�2�v�����K�k?�$i(gȻ��ʅ������
�}DܪI��!� �H3�	�����s؄H��������|�xh���G�k��q'�������w�i����k����	���F��e�>BY�d�:0z'��)�ߊ7%l��nk��пʇ��7ݩ��Mt+��������4z��}\��@�f�<�����Ǵ�~�!�/�K�@H��\�o�r�#Q�$n��tބ!�x�Y�K�U�R�}���2w#I���M�������DZip�A�*(ƨ+ê)m���N�oN�~�J�!S�d��h�k�m_&k:�({�	��U���Ά�N�Hh�vf�����Pn)s�x;vͲ�.�H�w��y�0OQ�b����L����O�)��=e���q�/��*:m@�H�����U�]o["K�4�b��G�Q��0��=���f���(UQ�T�����DL��n>��r�����:�:��w���v~�z��-���F�qo�r����~걮m��y4{�i��/�n~����������i���������x~��`��C���=� ��t�' ��}��T�2�I���M|�[�o��3�]�_-g(F����]���M���_l��=��4J��Ie��n(�/�/�/��e<v��_x|-���J�3��Z�5�N?�N�<�S�.d�.�q_��I9���C
�<X�@+7߼�mXB4l0������L���D�:
�J��F� �V]֢��C+`H��*�>��� � ����U�_Pv\�g�*zK�����&�����C����(VF9�ҡC��<�f�IS���kQ ��aF[(2*Q�p��쥥��gI �J̢��=8�/�3D������v4s�J�ѣ'$ϵ'O5Ot�n����P��ً�P* �$����b�U���Ż�\�P�f�����i�L#e��*���6�c�8�&��D���c����i�����տ�g��N�:E=O��x��f{�d��>i7�ߋ���b���B���e_��� ]�Q�|ãݟ���"��C��k��/�o_}�C������ͷװc~}�}���R�k�����u���(2O�t��\�|�p;u�T;r�hh`�����Kj]���n����fa��e{��T읝]�ֱ�R�N� ?����>>�@��R�l�ݻ��r=h/^�b']Y7��'}�7����(0.���۱m\<Ef	�Ԍ����ǧ��ݻws���;�Q�d���p���"�P�#NBc���J���c��v��:}��<q*'!;����;u��?w�]8!w���R���p��RT.�ޤ�_�h=m�<l�ߏ�u��m�w�=|p��x�����?p�\Ar�Ţ�9-����(X�h����%�^�|%k�|8�
m��Jz��:D���2*v�4�-�tTr�L&�G�ь�6Fl	�/G��!���7 n��Z��>�WΡ��^��Ⱦ�wd�����y1΂�CS��΁ �0 2����q+;a���O���@�Ye�{/s#���w�)4=�?c�����R��{������	��8�ݟ�](�$��|���Ώv�A����)?�aZY��#yM��?�L>�/����?=������=�Tږ��,�T<�0����������`��>ՙ	�B�@F�3Ed�8%�������t�%���e�$#=a�O�'H6t���YYH���A/� qO�> ���y�+l:m�{\�H���בM<��� i�Vq��Fe��	Ĕ9r�{����>���l=ͤ!�"S��HF��eʗ���증w�DJXd��{�sxO]nԩ�rx�h���_���q�w��g�T�2��t���*�*~�c���x,���������� �L���;���(#�m<��RPv�S�H��Bs���vR��p1��×�N���4m����c�8�Ƙ#�] @@Z�,4�N1��Y "����3H��Ҋ�Q�$�k`���Ifg�`�Ly���G0�S&(���.�,1�7�O"N�J��yh��'�����=!����.�QQ�.�*O���u����TB&�(B�K��1㲬���;�s^$:�K��o�#e�#GֽJ�0Z �Rˮ?�C*
z�%s	M�S�h
W�w�JEL�J�Q���$���ómҽ8(�֝m��̪�N���ŎSڭ���4?��M��@���=|�BR�Z���w�es"X%o|L�����z�>
a�W P�TB�'o�i��Xv�#�Q��6}��T��������� ��f{��&���픋�mmAO�ħ��m�Om�G��t��:
�R���ˡ.ԧ'���iğ�����_!�i������3�~&TYo�o��ﲏ��ЖK�>����[���?k��\�����Q�<�����w�������myŻ����(V;���J{���������n_w�}���v���v���v������o��������������?��7�m�~{�ݺ���#�ݻO�-8�b=x����{�~��z��_������Qf���t�ԡ��.!�]Y�.��p���!�Ʀi��g��2s�������Uv���Y�rEt��;��_<�N�=�=S���/Q �Ǐ�6O�T93^���u;�B�����厰O>��]�p>��l��|j/ʃK�ȗ�!��.�V֖�������((*E��=Z��Ss9�F^a��j9�r(xR�a�a�K�K�l�;�2c�~������A��ߌW	�ߌ����!.��^��O�۷oQGwړ'��Ң�l[9��G�*���Bۡ�6�9�ڙ�g��PO���V�wGfH�#��*�.�t=&�<��K�r9g�+���E�(]]�-�t���B2���������Ю*����Z�(���`����80o�	:.ē���K���=0�1�[e��=�q+�����x	�
*�1)� �Ue�/q�R��'R����0�?~;����99�M��a���׀i����z��%����+?� y�N��;��J�~7?��nZ��i�J9*anX�w���/Tp��#��:ؓR��,b<�2Τ���^R�����K��;���n��A-Q�̤���t�6(��;�m�$���L��_�R��&'&k�����:����Ξ::��h��N�@w��3~/s����^{��i%��3(�D�ݸ�7���r��%��?�+�=�n�pV"F����iT'�o�%+?�	=�� �W"��e�{�d�] ����~�5G��m��M����NNa��[k���P�wÔ�x�2 �O�*�ho�+܁��g��'@��0z��)N�/��S��M5D!�]7�u�Z�ȇ�r�u%�!�ݰo@�e�[wH��tw��R�ڥ���O�xP�)�p#�t�4�ЄvpSI���&Nx�2�B}�Sߞz4�ݓ�<1�S�G���-
�B։�yD�, {�_�7О���Z�� ����gaF �w�!��ȓj��=*\%�B����]˃jy�3%
o�e��m��]|gF^��qτK���r� ���͛��2�i�
G*s(~��K��ᢨ�dWu�~+eBA�y0��ʌ��4�b�:���wx;`]`�ʔx� �&�x�/�]�P�P!�d����I��(z�#�
���4���\���r���ʶ}�]��榇)���f7
�7y.I��K���)��RН!/�#�vμ�筶��,l���}����e�(�
�Y��i�_	Uҕ��e�h����S����v��i����ԛ��Ba�6���}fj�ռ�Z�<������;���s��D�"����*J����7߷/��U���۳�D,΢p�C����~�m��'�_~����Ͽo������~�e����w�]m_�d�����e�޼u'qm�8gy��\���6���ŵv�����?|K�ߠ��m�(�VV����b�� �e�%MF�P~!J he*J��aOt�u��ע���Y ���%
�&0~p��ε3�N���q��+g^���k�a[�Ez?��"��������_}�"���/�����ߎB!n@6�v]� ��((�����4m~�y��sgQJN� ��=y��#"�_3��|���{�l��*@���
B/�S5K�rL�;r���l�\y�䧟|�>|���S��}���g����r������#�IB�t�
�����zY���r�G����`u8h�k���u-�מThO(�cАe2��=-;|���k�����N
ec�����#��_H�r�3?z���kbPf����U�v����{�e�1�B\� e��|#��κ�n��9���HF�տ`�?��]�7����7�5����� a��8{C������*��+H<�!T{���m�W2i�,i�L�G���Tڲ�J<��ȵ��,���}˾1��?�zL��� _�O|��h�|������C^��q3\A	gء��x@%�#0R0�3;�괻���oZ�q�h�C���1z|�'�8��R��3 �@#Kȋ���7� ��������w�ۉ����|�A(/V8v��=����w��&���oA�t"ޓF�ͼ�4*Ϩ|��=O0���ü���7��|t��D@7���X��</��OCL�
ON� u�s �C��W�6~:Vb�8b��P�W����p^0�_?�&��^ʩi���}/��I�û�i���[��7�y��3��=&`{)�����7�џ�����_`�^��,CǕv�@N��)���`�{!���aϻ߉?�	]ws��'J���� �"�.�X�L<��(X�Kޣx�7އ�I�ա@/���Xw���#O���붍��=N.��u�]�+yP,�ǐ���d})`G�ϲ0g� �v!���|:�(��S��ŋ���5�	w ����'�3g1����UJ�;��`*h33ӡ���B.$��-e�1N;�����l�w�lY&;$�b��B�qJTp�8UZ���e�H��JeR3�?
���P!RLt���T^�W�?�e�S�)��I*�*�x��%�^'���H�文�tᎢ$έ&f=���8x�}M�Dr�YO֥K7[��Z]BhO0�F�>�ߙ RB	SyT��U�L��{�\h�ڧI�5�D��)���&�/�w�m<o4�;��3�δ+o�UG�c��sh�ayy3Ko޸Ӿ�����ڵk׳l���-x&��M�ء��o~h��������ߵ�����b�?�$}��u����������s�E��+G�]^Y'łSy�������Ki��9Jk�K/۳gR�
�5q/��d9r_�'Ν�����=6y��Q�깴U�+> ΢��ڌ` %k��l��#�(Xp%D�ؖ���Ժ-D��Y�lfv
e�h�|�|{��+���|�]���p*�*�ҧ������-ۤY�.�Q�Tt��u��z;��.]�����e;�t)� �.:�w��Ј�	�&�K�uPm_��Dg=w�3f.5<w�\{�w�g�~�>��3����4��/��y:w0[�C�r�;��;�(�,z��0�9��9�De�.�Ď�['�G�:��/il�I��-�6���^��C���`g�;��{}&z_R�n���y���_�i�)�Q�~�1�w%OSa'�����:�u������=P��է����K���W��7���_2�ɗ0C��'����i�/�*]���x�<��v ��`~�·U��la��V�a "a�;�{����%e4>�|ׯm�x�y.>���Un×���;^#��������@�y��G3��"�g*������@��*����C��,��m2����C�vy�0�h
/*Z

&��r�c9�|e�Ub�u�2աZ��n�;=�{��Ћ����x��N�G�0û�<��;�/��
��������I0o
�2� 2��ih��i�1�
�Ʒ[��CA���p�ﯱ�C���7���+��N��a�o׽~�L�������dt�;j7�Wy����-�f|�L�R֢3�����w7���`��6u����;H~`7h*�rILڻ[�W�63�I�k�u�(���7A��^nD{�Ð�l��y/��Rq'~��Q��?i�oU�o��jJ�r6�N��t���JD�� �0@`�8`+xFu�� jCT����E3
l/�eIxڅKgR6�(�xD���\jfZQ�6�T�8|轟�Qj��5��0�/=G��3��Bˣ�uV���w�ލ��P��LZ�k,��
������yO;Ζ�����0�h�>/Os/�T��A u)�mͲ�T��#!/m�zt�34*xVHǵ<��O���Z*P
�~ρ��̊u�A�@|eOT���N��R`]:���f��+]���.�Q�D�ՙ#5 ��}�.v�/��·�J�=�]�j(S���"��xz�J�R[Z����䛬�ó��6���2���l��hͼbtR�ch���pn~�t�q���G�X
�u�Dgu�`�D��}����ʕ+9�"�յ�}F�o���_~�^��~��Xx�83�~/���&M���Ä�߼�������o���}��w�˯�AI��ݹ� {�Ro��|���S�M���_��yQ>��*0�P���:�N�u�m�p6��+V��FT��q�n.�	u�U�Zd*�4��
��!�,M�L��i�F�e01>y�����:T�Fy����QfO�:�Μ9N{;J��v��\f���6A�E�(Y�㬷ǚ��A�'���ѧ��O>�8�s��g��x��H��*[�ӑ������Q�z�����O.؞�S	=���%W)w?v<{�T�>x�}�+Q���O�sJ%m8�J�%���}Bf�i+�+y }��C�eɂG�+Wx����8(bX'������]^]Π��|�SV�%�	��^���!3W)9iY~�E��Y�Gq�i�!o����o����>l��`v��7u�^30��L�e*����m���}P����CKC��.(��|G7*.I�]w-�M�2�Q��!�v�$�t���zO��3��I�X�d�0ţ���Q_��0h��/�����C�$��D�{���ߞ��!��=}v�I�#{e*������}�)�C����`4vj>.�I���}���8���4���8rU_P��E�6]�T4o!�n�x1_
硕�a�xL�����Nv3{ �'5G�����NƼ�W�״�ҥL�d��5��'��c̡�G��:�"w(ek�;~��:���o�v����N�)�M��"��� �7~�vթ�����?@��7n�M�vt����!R�C=��A��v~�Ž�*h��F��a�k���|�|�4��q�~�M⨇o���o���6��tt롍n~O<q���o�o�ߑ}�۞�ާ�:��\Gt�F�S
>� 3.��dw�_����8,'�˝�[$hL�t�/��cQ��r�o4�0ۄ/����PEQ2%�.��.x[&�;G�rd�ĸ6������~��P���̉�ئ��Gf=�f�B*�'k��Y}O�z����CP~;Ky�G:~���E!B�r��e?�._i/\�贊���
.O�<ɩe��e�� ��g�Y&	�Q�w��aW�2�fĻI��9� I�(g������wȈǥN����>����J�d�:����Ε%���P��@y��b��$�q�o?}XE��c�|��I^�z䈳
��1�����G�U?$�JV�p1�i:=��I��o����R��mu}%եz-3*�t���,���쑸�C ��6�{�8�R�c��Me"���z�ql����E�
����Q��b���h�Mx�4��y�&���������~�E޽�̴�9�g̒3N^����BY��y'������ɳv�^]���3���������/yo*�SN�����I9u�l;v�(�G�K��3qK{x��[�=�>�(�@�/h3nʟ���=A�(���?b.t�ezl���}��
���<�N��N7���u�����~hs�_h�z��cm����\�M��oܞt�r̓ԉ��>�Y��l��m�ȼ�޻(�5OS<w�\��'��>ZK����9<�[�;L�d���)HW�f�8�]g_��#x)�Gќ�.�P�~NL��.Av9�p8;>A�����yP��zx���(gy��\�<ޥz�f�ܨhѴh�E�k�.�Eɂ'�L3�Dm������n?PP}B�σ]e�o��wQn�����pv�uPQ�Di*w�W Hct+{�=�߈�g�I4|�J��}�;���0���Oށ�C�L2f�u�&q��m��{���ԝ8JyR�������Cw�%~t/��zv��y�O��4m��(��?Fʝ_�����.��;��#?���*5��0���H[������*�|��t�$�&�V�>�BwD����m�U��W!�i%6����̀�1�U��F�r��6>'^gTp&q f��Nt|�8&7۫�����!��>�I�S�<�{sM�MV)�����&�&y�v���J�L��}�|�߶i��n�}�)~܃�:�1���a.�˱��:N���0���|���{%����-Y���Բ���a���r�<ID�e�vo�V�W�گ���ܺ�������7�@�^�q
*� �!Ա� a�`�H� ��L��C���M�6&"r����1����[����q���v2H��'3l�ٙ`/�FNGM�j����t�T��ד�0ELt쯁W ��%g4p�o��/�7��`*ݍ�i�@p
.�PLp�{��UQت�\WA��0����p��{��T\�J��K�q�����ٗ4)����{�%�2��s?e�g�S?�M�m���^&�oӎ��O]rA�Q?�xȁ�0����W��V�W&5ME�S��R�H{Z2���p�����<�5� <��ש����84<n���(E㑑�~PV�8��$�uy��l���ew*>���[k缿��v�a��6�������Ѷ��rt��fp�
j�S�����/�#����F[APx��	��"�|	�@����JH����f�ˬO��l"8xB���3/��������v���v�������ҕ���p؍��O!��R@�}���>7׷�SQs(�޾�>�������S��B���>i_��=%��<l�o\o�n�Dp]"|՝Kж��{T�ӶI��}Cy�P9A��7��6	��:8֦��]����X�.֨w�D<��i <��_�e�����~���x�r͐�mA�����c*"����e�ޝ�9�̽ ��=F���Q��n�I�W�%42�����a��;6�ViO�H�df^O�=�=;��,c� ��	�CzT�.�}�"�=|H��Wg�<$#ˠ��$�˝|�%;�6�S:Vᙝ=��{�����~��v�ܕ�ۯ_������A��Cڶ�KiD�c\.*���X��5�#�CGY6�f�lc���sgڻo]h�/Ϸ�'��mkǏ�x�|�]�z��ዯ��_}��?�ߖW�{���C�H~&P~<`�M�[�eus�-#�nPn�&:��,�|lЮV���Fl��W�cx�8���g��j�^ZESC�����MS�ơ�#����6=G�'�'���Ĺ��wpM�*|�K[����
�a+U��v��v�⥜H8;?C���m��}m���.n��֗hC���z{����٧��޺���CC�z�xm߂�thn�M�җ��֡.�d�fjj�d�?9ێ�8mɒ\���h�;�f�t������������3�w��2�r3M;8@A �����'OҌ�]@��@��`�{����q�d�o�}�+d�B�y������Ǖ����v^���h7�ߞ>}����8�����Q�'i_�q����=@e}My-��O��1+�c��ޑ��w<��0=?S�4�J��)ڮ��F>��ϋ(���ۆ��Oߡ\�!��_~� ��l���jiqG�£�_y�������� N�
�Vg�i*m��?���"���S
���O�!��w�_	)m���jHP����4�JL~T-C�XS��|�6�]MF����x��e�绲�^�1���Ol� ���O�$Pe�}����e��2�E�tC"��)����~����#��@qd ZB�a��/��jp8_YZ�6y2�l@�O(���x��	��R%3aS�Y�Kt�� �6neM^gd��w�p�q��h��=��X�܆��2��N��mp��݌(�[�L�4ꌠ�$��nm��
C0����F#������)o�f4�C� u��P��$�Zr���[�%�K�*?3*������w���T^��Q�.Q !@޿*v�Q,��z�~��q�7��uԵ*N�������@.��'�
�`�=�)�n�H���3 t�@�1�QZU7�3a�ګ���B�N{���.a#�"�+p�/D���e��V�t/0�rK:I�
�O��,�H����o��:$�n� 锽����w �1�O�e&���+~�=��w���^u0��J��;`]��ǐ�*�E�Ug�f��o7�(��E<�ҷay-"�w�V�\�^I�S��|{��\���
��x�]���Nx��ޞ�� �C���d��}8���؞@�������L�a�my�[z�v�Mۖ#��gg�lWB��tf;(��Y9��6�z&]��%��U�害B��_�v-�^�~=���#��N9��ҡ3��d���gQ�<��X�n�p�b{�w�G��}��g���9��28Kv�����՟���G�����)�[� ����TYK�m���N(��[��>�%�F�����H��d����i�x?��s������?m��?���_���={�zP�nI˲��l.ut��x=�)¨��*DΚٱ)�(8�o4g��Lp���8U�)w���w�i��������c��Ge9Va�?ʧ�$�����尬��l����?�Gg
�c���^<_h�K��T��D����>m����(����t�.�\ݓ� �3#�;�R���Nڛ`�ձ�w7l+t�4���v��9��C��q{��w)��зeYY�i���k?��c�����U��{ݜ���Ӗ�04�i3}4�`B�|��Yۍ{w�}y�=������[�>6�w�W�K/T�,p�efVE��P�l���8��*%����a��<o�_,�U�{����g��Y����~����(�����=z�rhr��<~:��~��Oۯ~��v��9�g�l�ֳ3�;ԥ�)��~g��yā���g|�ɣa���N�!|��h\ҳ���i�33Sy�u�����m��K`1�'�;m��΍%pݩL�����{(�CC�&may�%<`�������z��{�6���Z��Ç�sO�7�|Ӿ����ӏ?�79/ﳞ$�dJg��҅K2�e�U����Kl7�S���hf���l���4a|���,�<iDJ=֏`�o��/L���K�@	�����޸�.+΂r�]{���cT�K*Ƙ̇e�_�6��A�ƫ�lӃ�|�R�0���׼ǉ�YF^ﻼ�M0\��� =�<{>�(��y���8��?��Y폾+�F��3z�=����2x��f٫����O�x�o����>�C�gx�o��'8̗�<Y����#3��俊���]��Ĺ���o��_�{�=|��^,��u�<���	,�X�������8\,s0�}� -FHSA \^�S���ݎf������ W��]� r���v���v���v�X��P��X�4\U%l��6�8q�-��	F+��0�Wm���c��^�I�&�(�i�����H����������RXf��/� d���¤�@;�R����o)(ƫoҫL��~�SH�
����B�ݸʍ�ߍ�<����'�{>���+����^{�V��\�~�N�܀{ ��3�ݴ�~���00��9���n��7��8��F��z1��i����ͼT|��0���~*������ˤ��.����� $w_e7=/ �@&V����y3����K�3��mP؍+���;�X5���v�{f�F�`/ba�6?�M�i��C��t,OaZa6K��O|� �~�	��,�}�[�����cS���S`��d��a��Ky|W�p��ĉ�(��Y7�=r$���?�;e>z�^.�-�����Wک��)�ʛ��w<mp��F)��U�� g��g�M�e�Æ���4����Q�i�ҥ�mfz.q���������([��/K�B���o.R�;���a*�*^.�\�b�'���g�*���lއ�}W8r�{Y\y�I��W.�?��[g
ފ����r��\¨"����"�Վ�8�:R�{A^��p." �@E؄V.3�	��}�t�bJ�Yd|*u� .\���47GƢ������ٱR�}�%!u�;�g�n��ޠO�0�K�;
ݡ�	��ʛt5���cs��R�O�>��+�5��栁K�ܷf��o�y���d���m .��2�Ai�{��	p�v�쳏�/>� ���F0�|��Q���o��_�~��j{p�8Uq��h��G����
ޑ`�ַ��8���o_i��V;s�T��� �
�mZ�/:��{����B��G�=��z�q^��g�q�x�%`�ݿ��ݹ�={�D��n=����i˚��:k�&.�t��3�V��m����c���o��.>��%��O5y���A�Yo��=�^�o�kO���I2�S��I��6x��1��P��M��@fz��I�p_�xuU��N���65��:}�P�iy��u_��M��B��������J��tV%���r<�����.�P�t���o8=U�e�ڣ��#��{�n޸�nܼ����>B�y�]/�����w��=y����K����uE}dN�#�����mzf��:y<�8��"|�*3�Y�|�A��5�/�re˘KB�Ļ�H���4^�Gk9���6�G�<(��
���}!�!��h�S3�/_��f�Zq����*�����x�w,#�[܇�R����~+��3\��>a_�(����>���|��8FL�=�o�V�޸����a7-���Ob��3HX�w|a���u>|+{�gߋ[b5���0��88�=~���WPq�/ȯxT�H��g�Q�~�ߦ����o�?27�N�8�Ξ:ގ=����m�������݇�v�,�\��r�R�2�0.iW�A;�%+Ģ��Y �ҁ3O��A��5s��&JL��[!Ŏ8'F���P�Bu�ıv&��6h�N>,���bu�B�J�&J���k�wT�C�Q�`��[
"2�!��ݮ�!�ש �͟��C������123�G�"���}���4�6��n��`�(�Q2��9�Gy�fi��A���V]�x�i5��?f)A]�a�GBy�@�0�Î^<tsH/��;de��s�O�:ÌB�)��=i����Y���<�H�s�L���y�R��0�iP)6���-��0�$����O�/���ӧXmٌ"��?�F�[O3���D�x����K,q��_�
��z5.3\�f�S�J^?u�~�c>Wu�/f��s�*���l��5�O6�!��Mcz�(
�!x�̡�g?����(�P&��ٳE�N�Y�3��9�5y��xh��|E�Q�r�����Q�Uq��
�����Oڽ�w��x���=�F��;���2��w��aXe�2�7b��8a
�������q�|�;!'��<u�L�'���u��{�����
a�F�=��ZS�"}�Y�hY�3gϦ��W�kޤ��OU���|��+���e�b�#�]�t�]�|%ʕ�9'Nz$�!�����у�e���"u�?�}���R����/��@ ����ٶ}K�\>�".n=<�6�|z���u���}י�������8���9��Pጲ�8�ag�:�"�6�/Mk��ZN����*Z�i������h���NU�S�����(Y��*�����d�)�^�s�no�T�d��6�.^�Ǐ�>|�}�ه(X�K��#������r������w�?��<�>�	K?��(X�`�h����(n�a�����g���O>��m�0*1ɫ�-��x����2����v�I�*��{�]�t.���'����1���ݸ���(
�a?ʾ��8{<�ջ�����q�{
�A�ϊ���z��J�����������>���u�4�1
�y_Y�h�<kׯ�m�}w�]��F���.1ևeA�:��v�J���57q9b��"�<E���g�qP�}Z�P�����Uق=Q���D�'�҉��e�*G��5k��{�{5����˄��� *P5p�B}/g�ʁ�+�z�� �z���������^���,�Gt��[�?���<��������={�B{���P��'\(&���mR?�(kgϝξ5�<�м9�*�|���b�b���d����2\f	�Kd�'�Rr�)���ӷ�a<��^�x.�=xڻ�3���wQ 1�="��g<C|��w�V@�U�������.�ߐ��נ I����[N;� ���
S��q`p�U`��]0��f�=O�1��+�LC{O�<��G�P���47�)�e��"�^OT&���_d$+Cs@h��䡊�D����JɪA]WD�ͺspRoտ�S���@��7�d�9u��86�!�������������O�ç/ۋ��R�\��
N�3T�'����VFT��r&���g���LR ;�*�_	3V�rĥ`��^���Yz��G�i��;�{��	������ѫ����|QfS���T�ྸ;���������:�(Y[m%�۶��K��ku�Y��2�:ũ**�ĎwM��z��@=���(�d�S��ɠ��:k�S�.K+���Ž��|�3������o���`h�!�$�ᦿ�ծ�n��+ T��r��aI�F�+xi0�(��#T�*S��%��cʞ2��^�!��0�R�_��e��R��ۘ�K��k8�9��G�7�*�,�^��e�ғu7�K')WL��r�W�A��UO�@xBe=n�p ��5����ػ[���x�O�-�(�p B7���a��|7|W8��|G(�[�Ǆ)���f��H4�ψ��(Tҡ$�K(S�r�q4������՞�;��S��&���Ħ��۹�g���ۙ�'�g^�[A��)�(g�T\<�O%�2
�n�;#�B�r������}C�n݌а̻������,�m>d¦��J�-Z�&�1sH���].ݺ�&�珴c(x�Q$N�g�p���#���r�WV�<���/��`�C�(Gǥ�X����U���Q�Ӯ��e�,.D(�xm
����G�ϱ��y�p�و��|�x�b��q��2��s��}��{����K��u�6zY�ʖv�}A�}M.CS�VYqT��yM�XY�]3�.�<�ru���a_x���Q<''�7��ʧK�AW�SɊ�	~�8Kᥬ��43����D��R��Џ:\��l�W��i�Q�)�����N�U�ө�nm��挎����Z�EI?١-�����$�=G�����~��O�8\�p�Qalm}u'�C����?�����_�{�}����� �+O<$�V������mU�w������g��%��	�Ñy���UOĵ�4𱶺J���`����#(W�Ϟ�R���(§�GirY�`�6u�]�z�=}�|�~�G�0��+~rj��i2�j�_�e��=�~Q�p��)��?B!�X�h{��̐��>�P:ڷ�\m��_�?|�M�z�f{��m��"�A����T�:{�,�ө��쓋�uZG�z�Rm�/��d!x�LM�����p����]��K]a�d��b��˗y���
�~����(�GQf�]��(zB.=��z��Ax��e˙�Eں��Q���n��r�������ť�����v���v����Ue.<���m��j6���S�ڹ�dy��3��A^Y�R�/���ۉ)�*%K��s��m�!H��Z��|�єq$�����E�ݾ&.�$�j�	Q��G�ݝ 	���Է|�� y��V=�}�}��r<��w�q+����G�E������û�gx���6��'Q���g�[=#�?��Oi��I�gd�fw.��� �.s���Xq�񻟌K���b����q������ȫIO,�k8He,����n4�?y�H;��u��� R�����տ�뻎X<��.���M�c̑�QI�Do'#�0?N]g�/H��Q)|�J��dx3f'��ú��f�\?M�O;�Hc+/�T�rY�&O�q٠G��!`��<XEώM�sSk)Yn|��hmem���\�����(W��HP���A����ur�[�T����'�B�t@�0��pv*�w�nu�e*P?Ɲ�_̓�2�
��Ox޳�5��+@cV�P�2n�4B��?$�*��{����x'J�7�R6	���n#+�����������,̧zO�q����{�L[��v5��{OC�;(��@����{��{���ޓh qZ>̚Q����^�\U�(��ow����v&��(�-߆r���%sI^H7f�{�/ܪHE���Y�ҭ�/nU�=��;�?=L��aP�Rf�<�6�7�T����@��<�m�ƅ��¡@��޳�x7�U�U����슴%�����y��S
�.]�7�hթ|�Ξ�R�>"O�;��u��%����P	A�Q���\z�]>�ݸ~��eX�G!�fRFx��*�휲�k�d�V<��y�|�~�WJe���9��l��0JeK�t8��&�2C��0�<��o�`=~�8���%)�IL_C>�3I\�Y!
��L�݂�GP&QV�n.�W!���/��;���{��J]�l��w���K�έ;��@��gG�8ሹK#]��a/m��`GJ�'
@��̒����E%X�����G����S�,VW7�=��~�ھ�����ի����iY�?mP�QQ؃,m�ࣀe���2�=$���J��jw9�Y�j~޺m�Ay �!���{�VQHd<��:���ɶI�d�<`���-�K͎�Q_�x����~��Oۇ���}<ʎm���B�ķn�,\��Zh��'C�^��ʓ�P���O,��&B���Z8�D�c�/���\�rt��>�h���G�4��,[Z^���e��(t�ё�<����{;J��E<ua�iy�~��:�|�=}����fP��*cX�	p�C� -YT
�yr�Y�H�@��0�K��%�Sm� <�"*',,,��?�n�7_��}�m�����ZY^��`�;V�qp�vJ���r��6GU�����/����d=*%�r��N�f�Q�Y/�Ea�Omm:C����!;O��x �v��-�haJk*Y��\	O���~|��r�ʺ��`�����#�B�l!ˀ���������1iN�(�<�Rf�N�'N�g/�=�t����G�%���9�80S3�������,�<{�6z���e��^k��y:䗋��ey�!�$�/l����6���d�m��dk��z�w�گ�=v������_��aj�
�[�_��5���ݬ��Bb~Pp��߄�;�3}'�=������-�(~�K��>���޼�[����<ũr:z�睧����^y���WFbO!R`Ͳ'f���~��>��"��3�`H/�t���~*��Ğp�я��i���O}�R~\�� uy�����]S���1�өv��|�xf����].�������G���%�ā���=Y���Ͱ'�%�޶��X�?Wɲ���n����M2"�T��r>+2��	7�*Hx�E)Y�&g��1:h��
���d�6R�0�R�L��/��k�VQ��\�ȜHB�>"R�&G3c:ZPGJ[���1HEXP�����~�$l�K�i�Tu������վ->:ZJX;t:)o���ݽl�S�	��zw)��`"DSE�q����i%O�=Lf�d~x'z
PE	/���z$iA@�/r�=�λi�ȿ�������H��Z���7��_���ၤ]y @�!��40�r�I�")��>�+���u�~��w��C����U~��w-|.%eG���42ԉ��Xm>�^i����bO`�+bK��{�5̀9BS�Q3�gR�~ �wp�b���ɏ�%�R��58|/3��I붻����uS
U-1�YA�'}�Q8pψ���T��p���W��*����l6GY�nzfP&�?�٬�O"�����.s�Rރ� Ð�ďЌ�����M���w�dI��Q�&|2�����7�v��h�2�.�Vys$�%>vn.�sY���{~
/��#�U�\/�ri�ݽ{�}����{�+��~�p�"�"*~���^ �&�
��ˀ
���\�73������&^Tl�wɃ6\��e�*��U;}����(>�RQsf��{s�~�m���~�n���
O*��������%���!S(�.����p��ԽʆJ�iZ���(�$q����֕�P�.�3g<
�X�i�=�����9��͛����ν�����R=�#M�V7���q�o�'u��S՝�].�@��)m9C�L��d���ޯ�Y�>��������U�#�X�:�.j[ѽi8𸾹�������S�a����PoA����J�x����{���w�+�c-��Gg{\*���=eGQ�=}���>(��eӴmy��3��O8{9׎ 4���D\ui��t5m߅gsrߙ3�h�ҞlShg���+��[�^io����p|xb�'	{��Rs��U���s�m?�hW�=������yL����tV�� ��̤\�r�]�t���ܷ��:���������o�M���~}��,�F�ٿ:�nr��K9�?t�,95u���8�8�r��U䥧�Pbg&�ْ���PhS(Z'��gt�(�����S�x���9+�]eJp�T�X]��)ʖ��TV��r�ji��0J��7�U����F]j(�r&,3W
J �Y��>^m�uG��?r<<��p��v��
]Bo�<L}�]��\�(Fy<}�4�j����IҠ�H߽�κ�@.��9��r�Emڇ����ٖ̜-U/�\��=����6�ǴȀ��Lk��9�|�O�����D$�ov��wdv;q�w������Q�ǟ�e�����2��w0�s��#J��ӓ��d~��{��`���S����aO����'�Cd&��LS���wh }j��Va;�Ry~J�|��m�ۘ����)e��)?����A�~V}C��ϜW?���jʳ�Y�(Y��S��v�4z˱�65�B�ɺ7ړ�rA8��f�Q\�GH��Fs���W�f�G���#P v ɘ
����^^�7tnG���
_vLnH<����	�"�8�������EgEX���>�zW�6Q��,���:��6�9�bǐ�p����P�c0��q܅��"�h���1�^�
S��;�`F!1�/S��Q%ܝ�B���)L�.�s�v��1�9�7R�H�U�����O5��{��D�##Q�Fy+.�+7�K��n$B�ԓ����Nq���	���9��#����R���Dy(K>�?�'>��<��oډ��a7�x��}���S�kbi��%}�o<�{�G��ɿ�i�>����G�Q�z�IK��Y�0I6�t7\��h#7����(�0z��W��aV��^��Uyح���M��Vfa�[�^��{ 
����/��x�c�K�&��pW�MZ�)�2s���4bg=�	�Y�C��x��m�\o�s�˲����U.%�VFІ%c������s�9bM!Gah)�z\��l��N��X�����������i����}��x��±wg��b�|��
���:��#������`�믿i�|�us	г����ViO�~޴j���,m�96�MeK�i��e��s�T��e��2����Lj>
�»����Mަ"����(7_C޾���a[�ҏ˹,��T!|��E��B�l�3X�@O��5�8חt:{�L��]"9z4K&U�ŗ]��xɮ#�?�t5
֝۷����CA^��K�/�5�>y/��o�рn�l&�ڲ?�}Z�(�Kշ��D;Jg{��ցCwp)�˅U�Ut���[/�:<��稇�(X|�~���_d�C��5�~Ӗ��W��Ӷ'�zٳ{^^5��=v�:;�YYg�ٽp�<��9�u����5�i��_|y��$iY'3ч�o��C(Z�f� uv����ͣ�=��zrfϙ.3/̾�rxE�����u�d�Y���������B��i���n��T�Uְ��P�+gw=t�-hT��;H���/C�'��ǥ�c(���e�z���k��_�}n�A�JMQ�S�a��Ӯg����B~<�b��#��G&�v����v{F�޻���v�rC�� �f
�8}�X;w�d;q�8;��^�k���O�D�FaR!��A������\r�=U�G�~�RJx��YYJ��љ+��zȅ3���	�.'�,�:VY���ٿr��,T��@!wf�{�nݹ�n�6��mu!��鸟�~F޼����'P�ϟ?�.BW��2�M��h}icf~W63�m�������"O�˭L�#�Կ�ms��0������sP|�`�W����В�z<y*T*�[���������R}q�O��L�W��	_΁^���F�%"��2 ���;�6�{)�䧿w���6����
�t��<��E��o��z/����'��X��* &P��Wю�~�@�%�d�{O���-�����P�)dʲ���զ#HG�����Odfg����P��ǜ�P����5J��G�ۣ�(YK4�~�E�g�MBT��#h.��Dɢ�ڈ�ɪb�G��x��J��T�)D@f�|E�!v��/�����LjX:�{	��-�o�k��r�M��E�r�{�b!��<
�;�]�+"�襋��>�[4x׏���3������5U�r�k ?t�e2�I~��H�6��Ȭ�D���&n;�?X�V�/^QT-?Q�����zѣ��$�VMx�7�de��πՑp�Ks�"#��:ȯ�XDX3E�{�*w�=~	?E���c��:1�0<j���r��v~�T��hL�n��C�ȸq������[bK�z�QY����^���{�k��J���˪Ŵ��Ѭ�(��0�9vʜvRI%��/��n~���Sy䯘�
����(��/~���\�8�:�ި3��)`WAf���2��~8KpP�4{�QD��{�[taZ�SPpP`t?�J��갱[�ǁOӎr���6P�<����<����a@!��4%�JT�eYn/^,d/�����C-�q���ϞD�Q�r�Y6p#�;��~�y/W���
��ݍ'V�n�(�g�;7���iʎ�V�W�2��$ۍ�7W�^m_~�B�U��4������?iTj�g��{�s�2�5�J]A�69�hq��|��	�=�������7�p�K˜r��N����wߵ�ׯgF+����*����t#��7>��y(���������ʗ����8�Re~ff< �eF��H���8Uܜݻ~���E�)u�)k�Kj@���ށ��0w鿻�hi�a��xy��+͚�ֆK�\F��xd�����I��8���;��C�Ϩ��$U�	��1���.�|�����﷏>�����ۙ�q/r��� �'��w�5��S�~���j��S.�=y!�|f�<���[W�:��n9�	c?�>.G�P o�������Y�З�e���8�x�%-O!t��
���\f]��ȋW.��9���o�:H���?�p�����v���������J�jZ<�@Z�*1
6Ό�6<�Σ��3�9���(�'N�f��>ys��{�F���k��v���,_s@��8q)�`�F�����#_C�kQގ�͑�'OΖ�����§�_R��۽����� ?o����Ȟ;�NK�(7.u���A�R6ڥ���U�2�Dyu׮��z���y�Q)��F�g�t�h�u|�ʚK8�
(Jҙr��>=��ҥ�����x;���o���(��P�oSG�0�����~8+0>g�Ϝ>�e��(���}���[x)߄�³l����l�G���;�&�/�q�>�n_��^� ���+>���7�_$P�啴\M�(���U���gc�ϟ���o��ߞp%�T������O=l��2����0;�[�������p���}/Ƚ�_����}d�%)i������}���;���C�����7�×6`�/�2L�Њ�L�S�~�S�q�I:�`��&�~�p�G��t�	'�;�#�*����v�ӇN�#��9���j��k�P�z�����%"R`�W��v*���;C;�,k�!zQ��N��?;L��P�(�>��IfS�Y䩐��2��������E��K
f:� T�`�Ƒ��j=w_x��#u(^���U!$B�3Aө�9U8�Z9z��'��
�A��:E��|� +��������T����$M�L�,/���Ly�L��{���Ф���PѠP\f�k�2R6+?8���wA]"�U���-	S����M�A|�t0�C�|�%��
0��|3�SH)�:M퐮u�^6X�6�y��p�kf6�đ�B��YqT�����=�� ~�W���?�>�٠����i�?��:�u3�G��wq<h�؝�.lM�X��a"�f��jg�|'����r3�Ą=y�b�8�\��JV1���ed�u��6�C'I��Y�4���� C��*�6J�
Vu����/s�@)I*L��8���PhE��X���O����,�q����s:z��<|���a��~s��͛�r2�]��5������ɓ�����B^A�ӽ�TR�ߒ��U�t�ûe�Y����l��N���Ic�[���p�0Fh��Gp�DP|��<ܸ���72:��2f�� ���D2 a�QWҎ'���[.����)�iW�r����i��+�pO�c�Žql�W\
q*��S��˯��=`�ZA0��|e�e�$Yѡ�as�,���3�S��r-g��m�ڀ쌼���e}�.|V��LG���������Y6�>�Foz����z���.|z}��'��ʹYM�L�n?X�*��H�s8��VW׳L����9.�;����S�hE��rQg�>�����+W��(8���-|�T�U����i�.?�.�����+�w����[o_�2���ɓ�T1w?���@�i�]W�8S��5��e�b��k�@�2˘�Q����X�UG����h�=|��˼nn:����'�,��o�3�N�4ytz� �3<)���Đ^�����:��%v**�s�|v�>�>մ�"2��8ܿ��}������]#���+�Q����襶��i�^��cm��e��P��uϟE�<ю�O�dN���W���v�0�G����6��r������ʥ��4
�a��j����T)��V�GMiºt	����&�;H$>�]U9kɨ<c#�-z���Y=��0�/�ص��(�q��C?4�R@� �m�� z�y�~�s�a{��ef�<�b�O]�����Y*x��ɜ�:77C~PQ ]����u������aO���*��X91��ч����ه�]�W�߸��}�GR�H��W~S ����S�!6�F���p���wO$���-y@�x�D�=`|���$s�?%�`"�4���i����f���0��Ra�ɛ?���=O�՟���!��������{��}�[�S�T?Zv��M�z�ң�[:ȯ�F&�n���O�|E�$���M�p��� �	;�"�J����;u<�θ2mm�_����_�{��/��d��17����#��6J`6���U '�@��5 �h<a�(?����^!GP]�25	��D�bn���Y<v ���3�2��U��~7	�.B	���*~�_#��T_�4o�_ZDP[q���"a�мfP�).�k�-��k̶�� ��{������n�tj��@��m��Qt�E�-��d�B0���J�>`���}<&��f����*iM9c51�&���.��ԑ}m;.]42��t�}��7���&�o�q	���O �8����4,��
С$͜j����kAE�w�M$O�QGF�ﺊeB��Zp��P�(����[�"�N�<A8�s�x��qG���&B�~�"��*C��c�9K�0]�y q�W� �!i�ka?i�q�%���?a����c���cϥ�B�B�	S~��t��mc���Q��Dc~�Gwgm5�&H���x/
��s:&:�I���hw2Z:�����%4Y�*>d
��2�$�F@��蒮aE��0e$��m���E����C�5�S�b���@Յu�L�4�(x�/�[G~k��B<�x	����U1~�5y��2m���m{s���m��8�����G���'���O��0U���()�mw��l���@��� �ߧ���P�L=QI{����ٓg�y��yF�U4�jJf�:��X�����������Dq�N 7����^dy��$x=����{m~�����w� �_�	b���/�@A�t�!w�H�,8�"^�GI#�ܰ��Qә���WV�ڋ�_g.�Q1}a�����B�S�{�^N6�T��?]��j�͏��r@�[��w��V�p��S��XQ,���VW<�|x>^��'���G+/ϟ/�O��m���������߶���ݺq�0ҍmJE�%��  }�t���P�G#��!�0
R�HmD	�^]b>��k���9�uv"u�W˱�I�/�(W�Y�DϞ=lt_���:��┙ڢ��b�O?o�{%�x��;Hߦb�Aq�k�_u�������ٞ�r��iO�<s��?���l;yb�?�B�@)<�Hrf�P�b�D��εP+(�=ӯ)�g������c��;+����gИq��N�#G�4Nt�Y|��������~���ؾ��t�i.��O�7{ҽyu�RV��>rq?J�+3�|���E�|�=Y Ƀ(�.;u9۾ܑ�E;X]ބ�_�^\^���4z�I�<��0J�4�~EeYŒ>	��28��)ʶyg�<�Y��<v��:�rat�,K;s
�Z]s�}\�w�}�����w�BY��rϔ�r�h#�#ؤR<Y�A�~���R�j6Z���),n*Y�?^���:ϑ�p��+_T������
���	�Y䫱��Cy���;c~�n�q�^{ \\��I'�t�{���f~��L7D��(w���k��2u�H,���ǲW�.��'�Ki�=l�����G��@wڢL�~�6�)�J'��j�
�"(	؆���=�n{��]���G%W\�$��72��.��$�7���<+���F�W��7���	�5��ӡ_+��ɢ�x�§�{���x#�)�a���k ڱ�x��s�� �;��v\��|�:����Vo  ĴIDAT��81��
����T���W��H̖� �p��WL�A�����t�ᇴ�e3<PuG��IVYMϙ����K[���k������Ə�CN���峧Om'�ε�䉶��?����z���tAc'�jػ��R���6�itg�ҩ�P}H�i�f��a]�'�yҗ����=�i���ˆ�؊iW''Q��e������fl"�������E:c�����A\����A%�LMe��7"�,��-7���<;�t��Mn	�P$q��Q��K����� �\ɽ���
cX"*?�t�n�0��=<dܡDQ�3Ssi�wl�+���~���I���pO:I�o`)�HNk�����3�^�����I)!�B	�*\�|��P9��!�!4V@GqP���/g��t�e	��S��=B8񍡘d�μ�^�>×���7�;rlC���Xt���\��8N�hd�1������2x��?����V)F�N�t����Ow߆�$\�g���w�frp���2f�uz�|��&�i�4��N�������V�c{r&���uf�wE�n��\n�?���a���m�i�Z��l�N3v�O|��Y��Y���"Ĩ��hq���g���q�Љ�^��p��{͇���A�Q|x�B��WKKG�yC瞁�@,"��}ˋY��l��<2C#��DHfn\z� #qy�M���������W>�0��3JW"�G%�Qi�:8z�2������rq+B��t8 eGb��a�|����˿��`���1~�,���pxj��;wr���[��-Ҽ}��Ӷ�,��n�n~~��'�ֻY~�ި��)3F�[�@>�S��ג#��I�.𭏗ԑ�ڝ�(�����1yP _L]��Ӌ�M��������ŉ�Lڅ��s��͌�`=��
� �?�P��g�_�q�.�Q���P�O-.-&�?|�c����s
�
�xs6 JC4�N�̋�^�|���vd~6����o�C�+��i�\Xo/�/��p��l2=�%�.�(ȫ@ll��ӭm���J3gN���7iց<�e��	]�M8sI�C�:ۨ4q�� �SE�%}.w5,܇�*��"�[& $@ۿ�^ܫ��,֭���+�(�of�t��>��HW�{ۙU�v�N:ӭgєK\ƻ�esk���(s�����о���,[��������
0�ٛMG&�x��ǐ+�8�w�d�؜9u2����(z���w�f������ٿsgO��޹�._>�f��m�d>��V�?�~��;�X�-_)vbXv���7ͣ��%�������ʷ'�j��ҁ����"��tXA� }�t�U
+k�=�x�}���[Fyw�K�|�~��ɢ.	� �З�����w2k��U��R{_X�����tv?��c"��ɯy���PF�Qmq�M~���R�_�
Wv�ѯ!E\x⡇�����n�)'��n�Q�j�7yL��ޡǳ�|������Փf��7x����4����O=?�/N����S�!Ϻ�W~�Wn�V_���y؍�?IW�.O�xU݇�e�o-��h�G?֛m0^���e=��BB�OÃ��:Ǐ���{g{��|;w�X;u�H����2�����������ŏwڵ�/ڋ��0�6	�t�i[9��y�����((�/`�K���Ȁ v�a2BA�#D��� x{4�a������m��4a��9Ҩ`�KaNS0�g�mjf��z�~`(�h��`��`���@��c0l;�5/�1�;R��8���I�� �eZ�0=+�N�NSSw�"ah�uV���QMAF��g?�٠�U���$yFU-��ܢ�ԯ�g2���9�wH��a�fo���W(�b�gH�p��A+\�ǝVˁ���Wi�
q82���"�+�!�סE{tn��2��~��&��}L��d�U΄'GM�S+��xJ�������I��xU��>XN�ոM����,�F�K�T~�����5�\e-o4�ġ���@b����|2£ɻ�%
"���|M���v��hG�U�ܟ�}4*�~�w|�'<u���sJ ��vZ!�H���(� �*����X��w�e|������=~0�V�K�ON��3Jn�(��Rn���q<�\m�-B�/���M�y��M��2>��ZYz��V��:|d�)<:��������m�-·@!=�g?�Nϫ��"\m�<E��݉�zU����8��������`Ғ�����P/��x��Ġ��eW���+�Ԟ4�(aܽ$&��ym�O�'���G87=����|���[.e>����r_�N��썋�!���ˡ`�iv��`yZ�JZ�g�&-���Ꮤ�64��x�C����Ig'��ʲg�4SW�}`�>� A�Д{��@Q�<MPS��:�poI�#�=��>R?U�g����)fF�[ ���+���ȇ�ɀ�4C��7Rҷ������>H�?�jG�m��#��6ys82��#T�m+.����Oۯ~�^N��ɍh1h�Fp+~��9[t��K�Q=�}1�A�������0��0n��`_��=x��]�q�]�v5�ڻ��[�Ҏ8���Ի�?��޻���N�t����I�*
��P�=J�a��Ν������7ߡ|��NgY��MiD��.2�@����>p�Z��Q��O����ގ#+���<��t�=�;��Ls	�̭cc���[!�KfD���ω(y.�t���&��+W.P�������?hǡ��{����/�n_~�m�v�n���eʲӎӞ>x�J���y���w	3�z�n������ȟ��e=K��qL��S�Q�*���y@���Q����0��e�
���������c<*�қe=q�t;z�d;��9u���������ﯷ7�/���9�o\������ydn�]8{�����v�vhB�mf������������my�>yj�|��d��U��3�?���{���gm�Y
�I�'8�~�����~O�����^r[�x��_^�[=���������{�,�_���=r��h���V�ݝ�$�����^~���7����'e��o)I��<��n��>{��e��i����l�B�Ѓ�x��F��Iچ�&䣴}s2/���ޓ�x�n�e7u�=g
sm�dp�輒azr�]8s�}�����O�k�{����Ӷ���?��w]ɺ����=_V�B�o�¸���Y�,�z���@��r��>(X���tT�%:�F�z�F���D�Z��~��I��xll6�+P8*����t��s�0��Y��>,GgM{��7��T�@�̗���a��T���W�:Lal�c(^�9qhs��
r9�4����6����H�,t���4i6qÄKX����J\�����N�T��A��,���c���{���߹w��u�'��QVG#��f��Qa�8�b��k���ҿ��ba$$��q�Ybf��c�O���t8����Y&*�ӫ����x͔����-3Qx-��@�i*�\f	�.H�v���0I�+Y��M:�#,�g�(k�O�ݺ�f�z~z����]�8�S0�LA��Q7�K�:�6�Q���w��nO5�6̀�n<~{M�y9#cݫTd�2
V	ĥd��bQh�4)���������|�$�~���r����њ�ִ�+\9���z�=>���\��S�s���duz�l4��+�͍,��Ō�Z~4���Y0���x��㶂����#>�}�&U�q�A+/�:����c��CTBбh��+́�(Y�q��QJ����+�O�<K�3_,rϬ}��nl4�!y�!)������V�Lҕ��|�#3�̤7zqMw��+@,���ꪬ��3+������OfUWcL��Ȉ������~�H�:O0�CF��A��X��x��V�%S�e��d�)��,=�A���"��XO����S�dN6Y8��ixf��q��fÖ[Gчp�
��s#�Ǧ���a���96R\Y:��oY�Chj�~6v��0>9�I���pyQ /��d��tD�`��K�Ve�q��]��E���;���n�����U�rQ��14����!rʉ��.��T�����N2���U8%j�1��dC�I!���'ԧ��<s��m�mZ�<#�m���|�B�S���rb^{���ߔ�uAr�(|����Z�]!�D���8k�C_z�oZ=+��[���O��em�5�����q�����=9,\m��ggn����?�/;�ꫣh2�K���ŗ^�.\���^x�o��\=��Io�ݿ�q��m�3>��9����|J6�'t�eɀ��Wh�G�:��G���|�뙛���*�{���]?�����Y�C�r��8W+l��hi��W�x�>�y@�P�^�-�Y����w�9~�_}o���o���ؔ]���'��`��_���Ɵȑ�T{�M;�|Y{��}��ַ�>������-�+��3�x��
֖_ �|���q��O���O�pU�z�K�{y�'�z�X\�|�3�0�Ǳe�d'Urb�|s�,oE��Hc�!�c�B��i��$�֋{r?�sw���_�k����q�����Ɉ�HH������]��V�K�?3�|����W_��=�;<�y��x�W�_����+�����4o�׷|����0�<����<Ϙ�%eN�*2�PR�6�>TE�I
�rH��X���t	�Ăq���ѥ��w^��u}���B����,�m-��<Q0U<ў���Y����}9	3z�>N��6��0���tt�QY��yѲ<�7�먙�'�0�@�*%ض+���q̺�k����Ӽm�<Ny���X���W�7W�+/?;���k�Goc�������8Y��?����,'�︒���qgG��e��MMJ1'���r��d-����W{>G|�����,�_1�̀���e��Z@.ʨ�Pm���~�[�"g�s�V��ǻ�C�ׯ�
���<��q(���T���c%GZ<�_��fmpBx~�!g�93��`d��<h+__ݐa��(c�I�b��X$���&ys+�ĳ`c� �:�ona$mG˛I��yཉsW3h2�88u8E�,�݋���J�<$��ld������s��'<r��o�A�Ph-&���M6vj�΂� ��%O��O|�o�����y66� �+,`�nB�dT:8��<|���^��㍸d@�d�no�:�C�j�6�0�#�:%ʙ<���c&"?��I�Q��F���4N~��C-;o�UD��8pzLzCc����ڰa����WE#�fy_'�C�m��x8�����1/{1e�5ϼ o\'߹˕'X,Y�M�V?Չ���0�����oO��%8o�\"�ZzA��?���ĉo��q�-]Q��q�x������ʦlk��P�?�|�.�j6�`WN֝�n���w''K��oS��[��\q5�P���J^�`���	�)x���Bg�D#�8<X��۫,}t�T�Ҝ�	�c&=�c2M�b3����RXG�$�W�x�m�nb
Z\�-�@�}]���%�ǜ��%���!�⍙q��A�E6D���%��
�6N�uUeЊ�@籍�rk�o��-@J,����%�J�J��l1'ø���KX0�s��*g�H3Fl��9WïǈX�*c}�86�9�3��9�D�N�W���ģG�j'8o޹=��>k�+2��-Rd��gn��,W
p�\�3<~v�H��-1�}c�g����~������ݻw��{w�����/ə��|gjߎN�!p���o���Π#<�e��3gQ���?��9P���׻��t�3�q��^��!g�,��Av�g���=Ș�n��!�!�˪\r�'[a�z�q��\��`C�1a|�lަ'�q�A9+�5��qR���לaC�ȸpR[}6M��W̵���->���`���`��_��6c|��G�o��oǟ���w�0�������s�;˭�7�]/�pSNȵq������8H� 7��J2W��/�����/�A�1u�>rX�vӏ?�<q�x��f���g�R�{��W������'o�+�[��� �om�ۺ(]]�썏n����c�w�l=�>���I2^�$�r����Dr�4>|d�������k��8K���so[�ڇ㗿~_��a{�[Jk�̞h�H��43�y&K��s��)����O�Y�2?5�-�X�E�-��	�#���-B�|�?��ǀ��\�>d�+_�|��	��6�}0�l`�j������% s����\�X�5�������DD��b�K�tBd
�6�Ӱ\�����)$�T�z�4�},��/R�v�L�̚c�o;N.�`�x&�5���K�xy�v��aV[�=��1(rR�������x�kύ�����������_��e�������]�z��!�$'��Lp{�D��C^,���s�.�pr�9�N=X,W�0~(�
�kA�26��`��f1��ھ{W^ ߸ѦGD�}�Bƭ.�a�z���&���{�6Z�e�E|�b�͆�#����2t�u	Iܽ��7�Ψ��U��1U�L86��]���M����-
9O�l�9�;��A�������Y
?Oa���r�2��T`$���4�,���@�m�քae���bx�k�u��0��R ����؛)����ʭQDգ��������f� x�_̫d�F�#�����ݫg	1J&#9��p����A?����SX���x��V���6}H��r|o���3n��o��h�gBorR�I#��_;YW��"�٧���U�!��۷;�W������ly>�M��d-�9�d��j�7�HJy[振6"�1a0:�<���x!$�qKL��(ZN)cl��1�"?�]��I;Y1*��2�訆���o6h�)W�|�:�Ng��vGtK;ތu �j�����
���يl6#��a��՝۟���z�AR��z�;�d#v��-�{�����/��k%r�y�.�qD݋��d�'t�M���R����`�iS�t��8��fi���$%ܲ��[���8�l��͓�����1���O`�o��G/�S�r `ː%��?��1�Y9v�1�^tD'z�:6�<�6O�=�/��rP���4�S�MP���,�����3Z��1��g��:⇰ݿ�	�>�������=*;I9j8��'�)�s��ܡa�"OFש�j�\�>�F{�s��ڠ�)�9vcS�l�}�ƠǄ�c�2!ߐsƳU� ~�>'%�[���e��q���b���ig[4��//��^^�8����op��Ø��<�6��'j��f]f֛/�'@7����/���5��W�>��];q�s ��uz��2H�$��M>�̳zr�5����dbڲ�Z��C���c��/����Ǹ��H�c�A����1gZ�:N�p��Y�wĭȲ�W�l��_xf����h���3���7�K/�T����������t��?����y������rx���ǵK㦜���>^}�%9]ύ�����~p"�g.��w�'}4lo��W�xc����Gr�x*�%�,n�e� �<_y��U_�j��+��V��W_�Q�_�H�އ���'�]����v�Y9�����n���������pg��fƣ������W��؈�������y��x�/�o���W��GG�"p_N��}2~%'�W|8>��=�����g�y��Ԃ��I#�Y��oZ���X�\�8`����j��1dl+�=52��$��`<C�p����wN8��c/2��SIcG��`K|zN࡝��u�$����Z���˂���~I`B��q�l��\`�S��Ά.3�⯩gl36���O�4)�����������41_�0����j/A��g�ȝ��X�=�1K�r��]�����x���o��⸼r�+Yv���g�������8Y��$<le�p>�w���������pr�'�+Y�)���F���-J��J�Í��jóX�t�E��9o�+�S٨q5�"gʹ���h�sVeG8֢�c�1�����l��|s�L��|x��/]�a�%�n�EW�m��s�8miqBt�����y��3x��%��p�'?
��c��(X����1� D�͆���㿩&g�y^6����js�[�(Sc��
l��P~u�q+��E�_����y�4�~��8Ŏ(�t����%�ci�S#�;�
����'u�G�ha85�q�pZ5.�Iu�-8H�B�w�'����S�1����SXY�Og̓�$RI'��Q��`�zcǜp7U=�F��͙҄}6Z��'�㶔v�$�W�q�y�M.r��B ��^?i�e`��{6�	񊌈����<��J��[��=�\I %��-�2%u����y�Q��0h�_z �l�9'K��T9X�>�q���7��]��X�y(9�&��1'y#�%�r����� pf�vi���������{c�o�̎/���6lR٠�!����0:�@�@������K�郝cE��fy�0����@[���E��M�������r�)��c��`#E����pK8�ɧ�>���n�2�-�lrDD3Ϥ����I`��N:"�ܼD��ӤJ���MNz���a��<��dN`�c��pƞ�d1�#�dq�ou��QD��	�y���s��p+Yqe&t4����w�]���n����i�M��oMe�.=��i&;�m
/�~���|���F��Y?��Q����Z\�?�T���5B�'�Þ�!��W����́T'ݕcJt�����>
�b¤���(�"x�I�JN#�!'>γ7v�Ԃ�l��vBmx�>'
Z�bC�D��Bg}�o�i��8 �����G��p��2��?t�7��799��5��� k� '��,�`;f;�����9�W�$='��w������;����x�ŋ�]�{c���?��O�t�����8�V��3%'�/���[�Ǹ��j��o�6~�������/��.�����?xߟ��-��q��0��4�n}�����!N�_�7ރIf\�ř��w�^�(���+r�؇���_����v�.l]�x�[��W��}���������o������ϳ�xY2�J���3�s�9ߐ}����7����uQ�63�}g�h|��m;Y?��I9ye�����4��$��A��Q���<����SA]��?Et��<�b��L��tX���hJ�����yjp��Q��:D;xm�3�(�>���	�V�����|�@�h������D�L&������"g�>DN�����Ewi[E���IJ�ؓ)p�(:G嶛B�ڍ��.;n�g|q��)�r����e�,prrpr�TȘ�ɺ�1�x��������ʋ���va���.8w���HYV��xC�Ncԟ�d��g�Pd���R�6VT�������W�l&����5~6c(1_gXe�mT�wyu}����,���?)/'���EE�Pɑ�1�&�#z(�{��z�rmGI�����9�/��/�}�	��W�AaÆ��I`aBD�뇵}�[��u�P(��3J���'<�����B%��l�h�F\(��?�-Š�7�|W�����[�sL�B�,��c-�8Ɓ�'/�dQU���h�?-��]�:�tu��J<[�Ǝ�U����x>	.�jX�w[Qb'�^����h����2�۸�K�I��!L�Y�þ��<����g,8�
dE�A4�(di��"o�L�d��K��dƆ��n4~]�1�X�����q�J��/��I���5�L�#����4�-x���T�`~(�#Ԙ���W���^�+��(��։�r�d�v*��u8��k�c�<D���f�o��1�l$��3śÐ��"�R�6�߿3��|l߻=>�sk<ؾ-���o
�D?�?%3F��T��=�?�I9�φ[���H[o��s��l���A��)>�����t���f9:����܃��|Sۖ�
�lB	������w�1�{��W����v�^����♑w�3���uA�\:N��`S/�/�\Ǌٌ�/�W/ؠ�yD��+��+'��'t\����gɉ�N�-}oۙW���ņ��%�n���C�ܯ�x6��_�$�	�|;��x�c��E��:�Z�ӱ�3��+�c��8Y�8��8YP��	�TS������3Z�8�s6���u��C�q����:n�S�-�^���~�M�ñAVq��N��׸��!F�~Δy_��ZH���MA��Z��\2��6�J�^��]먢�!���Ȇy�k��	:��S`�͜,�窚�_8�?Ą��$Ƃ9Ɖ��w�ď$\�~i��G������o}{|�+�ޜˇ����������?���7��sl?�WvoI�sz���d\��>���K�������v�._��>,����ƻ�xw��?�>��'�x�)r�#r�y*ߜ"�7A��Ň�y��?�f"G����VD^�j�#�_�_�b���W�\���5���ۚ㽏n�������w���w�`-i�%����R��C1~�P*}��5��[㕯�4��η�[���(��@����[�����{�r�>��ָ'�|�1[o�Z/9x��dѸ2����"���Q?�)Tv��)�ƙ��i�!̓��\���u�����s��E���I9�y -ژ	��|r��s&L�UFI�Yx��}���I�6���o�Z����3�É]�Y�y�>�l8&�;$�a�|��?wj�{�r�T�*�/��R���{h�ƕg[y���S����Wޱ�q���Ut���.]?��/o��zi��{r�������؍��_�d���������]	teKNo�3ڲ���vAM��7lx� /�8��4����i��X)h�N���,������HZ�eyEv�7�  ���
ޔ�֑6b|/�C�Ω{��������
.�ŗ��(Rv��o���-q%�'��8�ϕ6�Ŕ���<�d���(v�4��g�a� ��ԉ����B�B�EM�I(��J����ucR��R=Ox���+6ꋯ� 'N�B3�������3/�1Dp�d�o���J���M9�v�b�˽�.�?�g>h�H(~�~i�4�?�>~/��.mI��V��h�^��:����v]A~q���G�7~�N�&lo�hg�%�g�|��a�BW�	�U�l��ϲ����T֤�-����%z�h�W�2���9	�N�o��.��e��ڦ��y>Uqu�<�z�C������Ju�O{M�9��j%�Eʘ���Q����cm���dqK��qж6�o4�����,W�_�;:�~:n�d�w?�T�gr�������'�W��a$`,�o���r"�8�O��
��U�3f�e���"`�*���uL�m���~)R��l�UI��.��I���{�a��9C;T��v/��x<)סK�'���Yo~���1tXp�߾� ���<�-|��� <�b��[hF}���7��v�	����=v.�C�e�M_s�&��t!c�s�@h�~M�7(��\l`ih�����j�8���������^���t�\=�4%pD'���cNrHz�A��%<rb�s�֒'6Ѭ
90_�ܲdA[� n��؈O-|7>��_�=�؀��26���$;��"���=��N/�2�MW���uO1���F�Ð�l�rN/��X�D��3��D��ʐ�/�����gҌ�"��!i{U��<'^���|���}N������
�7 &�����xê�Oȟ���f���C���/���;ߓC�[���}k��կ�����;Y��/�b������ǲ��_�μ��8>ܕ��}K�w�����?���_����{V�7�L�;���'~�+^�K6���M���}g����m?�����(�����l]��<�������+^���M�ʶ{)]��C�<�������?����K�֝�����Wr�>������q�{M�a]����a���z�~.���_{�����;���w�d��� ;�Oo������ͭO�]^⥹��/�ʢ�@�m�����{���%0o�?����L���Y@�a�9�<���*+4�:��ʃ�o��E�RҴ&�+� '�h�?�s�O��~��GJCF�J�6T�s���h�?��,�,��7�ӌ~پ:NfA�eq�ɪ��#�8�����"0�F�3L��|2/{�Oc��lx�B�Ʊ�O.��Vq{3W~�a�x��t�����g�,P�fY�Z�C�rU�����k\�z�W�����r�v4{�d�?��?�����}0~����d���a��MM�˗0\8Y4������~o���J{]�����/,p'՞��X�(�0��j;J��l�d��9�r�#�f��*_��=����8X<���P@�+WVJm\y�ƪ���B���X���z�� g���� !�3O6h�#��O���KHz"ΐr����R��� ؄��"�r�'jI͙M)�F�E��\�Kɣ7ɾ$za%��,q�2��Nn��F"�&�麪��Qw6 ��
27:�����e	�	~ƚF�����b3 n�K9m5� #p1��Q��y���$}U�|?hE��hƹ7^�S�6���l��?!#τ���c�N�"*�s�=�,�v2�O6 |6�g�S��o�n�}��Xf�A�`���o�O��Qz�f@��g޸ʶ�<8���"d���%n��������@�1z��"u�5n��K68Y��ŝ�q"+XQk"�E�[9�bp�8�ĭ$\�~d�3)8p�6�q�℧�#9Yw�΃<�u���q_�֎�,��!W�oW�a�~H�70�L��K���9�	���t�z.�_e;p(�ˀ�̇ ��\�})'S����Y��U�>�g<������;���,vz���7�O:+\�_'$��r�8g�G�Fv�/��`�>�)WUT�P����#;x�;d<=W�ek'�P釪��}3O:F;	�_����� 1}&�?RxA� ���q�88��ͷp�����$�a��g�
�e��]?�X���Y�ʹ���鏝c<���'�j?�%}
o�/s��g�8a�1�ȉM������F2�|m�9�Q��O��#�jLX�q2�'��m��[j��C27��ȇ��rg̠�[����g�Va�����<�Ov��<��&���Vzp�S�X�.�|��5��n�u��M���+�q��ߓ��I�N�N?�y�S�ȱ��,�8�rQռ�y�[OZ�ON�p�A��Z�{�;��[�o�=^�Y�]y8~��_���˿.G�'rP66�]3�ғ�=�.���>������5���`\�|Y�[��;��x�!�_���r�x���l���'\�����w��G>�Ҳ���kr�.��Ꮚ�qE�c�/�f�_:��{�����������;?��q�򸳭��������c^!/{|��,oH��7�K����h)yoɾ���K������=9Y[�7/T9v�'�ޑ���x���'wn�{8��U?�Bcb�3p/�[��4��`����E~�<9�o8���2�� �)[9R�����Sp�-�H>l����Se�_�M���DhC����i�s��� �����+9R��@k��[�w�C�/��b�&X��B0�e��&A>X�8P8��!�sX�=�(Z6r��Vt�'�;Ȓ+��^�t�
&�=�����&���Õ�V�o'K�+E��%\'���ﵓ�+����������l��O>��h{����l��g�$W�r�Υ-m��H��8����n��%|Cm�$�G��U����J���A&�12�N0�dZyX�Q�R\�-�x���Pm9�N�l X��A���� ��/�������#�6�����Qx򼘂�l6��`�l����J���?�B�ء�@;G�٘) C�Y�#�>m���ތ�G���d��"/X���X�	�)旳46��6�*̲���8���LưC�`�%����gI����iA}3�E��P2m��W�:T,`|f����9��e*Y���}�hH�|˗`��e�IZN���z�UI���an�Ks�MgVu�> ����8�/�*h/��l=hyL�@3�]�&)����#������r*����`��r��6�,%���x�\�����Hs��Ù�C�=n���n���p|��>F.ȍ�R7y�\_�s?���cW�l��}?��g�Ti�c#��sG��D����4]7��]���Ϻ�<��1��w�l���t��9�0m��+4�Y�u��-�2%3�� �`g�L�+!�}x9��2l�T m���)��ɱ���crp;�OUe�ӏ�&W���~̓Ɔ����|o,u�12�B3��]���zuVn�`:J��|J
E7�������`�H�?`�)�3��]�	O�L�}���s�?�蟥P��BLS �˙S懐�િ���e���)q�q�����@��:dtĸ]����=���c�+�E�#� �q��$�o��ķ�J*�8o���8Ҝg�m������++���|c����������x�����~������������?���h���Er�*o8����㙛W�w����G����_����D���θu���ӟ��W��������d��W��������J�iO���t��e�,ۆs��|�oi!N�ᄢS8e��mpRA�}����[��;��3N�6ǭ;�����}pk�����g�팇�Z�i�mIv<>"������>�Aqkce|���o	�o���ȋ��[|�������?����q��Eyk���'_�.�0�+���G��ҭa�\/��h�ט�L �_(�0��pa�(��ƆFfN�Ǯ��X���{����Ӽ��{"
N`�=CL���[�>�tgC�w�4p����2!k���ԟ4ʘ8��r�)���Pi�����o{�{�_���)Pƕr4��i�mr�i<xfS��ѱ]�@����x)o�d�����f�������I��r��b� �0����\�0��ڋ���~m������<��~�eF��?��ON���,'�C�,�Y�8�N�(	�7q�͇p/mic�F��<d~WN�CM�]3��z�0q8���MB����	e3��A
�W�W#�[�Jpث.����,�ތ
�y�@ra�%��4/����!��<q5�<Af�b#��*ܫ͞:ȶ�m5d&|��\!�[	{�>��F̔c,�<	_��eR�L|L��vF}��=Q��d"x���i�4�#�g9J�E�1����"=)4!~IH�l��d@(�Z���C�h�B_-�4ɕ�sȞ��?�	����U&`EI���%�+\���c�i��Xz�8ۑRD�"��Be�S3��0�\rƨ�ACw��J6<;Z@XNL���<t�c;�p����!ݗi�F��R�F H͑4Y���g���F�ls� W��[�����8��b>��Ƃ�v���#��pL�S�^��}�c�r��#g�WT�l��6���3w����4�m��.�(mT��1R��g�ěKdCȇ��'e��RC�v�(���(g���q�)��������7�o�����ס�G�Pg;�@9:%���qE�K��rl]�� ��N|�׿9�Ʃ �L�Ƨ:�N��z��7,s���[\�5WG����Y�E�6����m螙3����s.m�l-������!��
�V�#�:s6�?N��P0�
�v:�N)NS��DhdO�g+,��Sd�r����6W�p��p)� �jh�K'[r�֘�F�"�-���8�ǎ������{����ƛ_�z���x������Q��ߏ�������}�!'Z�9�,2�����;�ys�ɟ�������'��ŋcI{��w?�x��?�q�����Gչ괷�]|Rf�N��#Z/���gIp���{w?�?�5>�{�N�o[W?{��/�9��.���/�4~��p����흃��{����O>�'��ָ}{o�x<����"W����\}eZ���������+_o�{����`����(����������*?Җ���7~�P�FR���Fc!�MJ=�)����*c��B��C�+���V$�b�Z3C�jO��)̮��#R6����[��!�8�ޗ�b��
��1t���@?G�3�A�^�������,,x��xc�8vR�B2nK̥E�j}E��Z�4��rP�FG^ɔg�RJB�>�	 %�,��V;^�G!�.��M��,���P����SQ~.Vٻ�X�&{�̩���*��.z�����׿����7�d}�u_պ��4�����w���O�[��{4��gXZY�^�_3�憷q3�6>ǚ,\v�
���N�|��?���ܕ��30�\�BAc�3uv^A��d�f��V�N ��g(t��?(�FT���_ymk}K����k��?�h����=��꿎y��PA�
}6�J�m�D�v$]�-�ܺ���<Q��C0�?�6���ӆ���y�W[�"C8�-��?}$b@�Wm����w�j�XS�sh]�ܰ�i��7��O�:~jdA}G�WYG����Jg���R&#�M"yމ���N���7>̇t�S"�jJ�v�c͑#-�G�㫔��yݮ뎎���9^^H�����x�b��r����W=��G;�¯xLzH^t�?�c>��<�j�+�j��\uJ�r�=�y; W����9�}��]�݇۾m��|>���x�}wܿ�� ��)����{>�}p���w��P$=��;�iR��F��~��}�]m&8��Y\�L�Y(6_���$M-z(��<V.sL�"Rc�0�5����s���1�Pi���ܹv)�����98��p��t�r�E�E42��/'-�u���u^9�Tm	UN����ǘ��ei�:R�R6�F��3���l�F�rh%g[�R�
'�r���#���N�i���)-7�z�&�_�a�ݤd���k��iW�S����Ut>NDʂϼ�D�-����;����*'D�:��B�c�b��3I�0?~rtS�TL1|�e�>Ǧ�އڤ�\]�)��c�B.i�=��w�N���7��׿��x�����^�:67Y�W�ݻ�ǭ[��'�|:>� +@Կ���Ƞ�n��8�u�����k��W�:^{�U�	�e��~���~��9���eOwl?y�*χk`>��(��Q|���G���g�*�]扷�m�+W�������o�g^xa�����n�˩�����/���@g�������c��?��x����s�<+�rݷb�/�?�\x�*v{<�]��#䶢�%�Q���XR�ž��WI�v���Č��.w��GT"8u<���{J*8��u�� ����'����zUO��}Q���Ix)�<��/�����0x`%��
m��hX��2N�T��C��E��||H��U^Y���,;����Ѡ�8���)��3�a�E�/3��Cn�>��ۉ��T[��?�R�7DÏ��������l�s�\7��C��z��������[����~p��%B��I�R)����5q��|b�4���Yx֑K������-�͸���ۑ���Nc
	x��V��+�M�,;f��߯(F �H;2~e��&2�ja�G�|+��
�p��Dg����P�(�����gM�����^��Ue�p����[��z��z^X����������L�W�pQ�H+2�2(�:*P_��٥mצ<Η┊Y�8.O�(��*5z�����q	�-i�,��]�p���m�)x����I�d��!��j#��ʪ<|H�����E�Ѱ'��㊜�t:9cj�0q�䡨X��R�S�(-�K�U�2�si�4E��o���Iy#�p8�B�s�Qh���%mF�Sћ�w��p��U.�L�#9]8h8_�y;b���sV�YI�#m6p�p���ړ��w��v������p�t�C�3u��~d��g}��?�p�ә<�-�VC���X����`/�ͪ�����;(O���:��_�l� s�"��ؼ�ӛx�JS�q�a+
�y՟ȅh�.��J9)����W�y�3�����"�:�]�;�P��S�Bo�d�H˟qW�:��V�V�:&Bc~�2�
��˨+\���{o��k���4�:�ł�����c�\��s�����`vꓒ��HI?Ƃ[�Yo���(A
��*���׆5<����,�W�aҮ/�3��U\�W��~~L;�:?����y�_�.c _ȴp�f]�#�
�ٕ܀�@|ś+Y8e���W�eS�y��x�o�����x��KڿȬ��ݻ� ��-�~���@x�G7_�����W�y���������۟�[~0>��C���}��ʕxnu���q���.���l�)}7 g�y`�o{l?#���:$��uq\�vc<��K�7�16.]�~~o|����}��g�����ng�,�������@9Y��@�7o��k�9���\�s�����l��Wɛ�Z�� �7�^� �������֡�1�ʐ΢�~~l�P�ˢa�MC��ׄ*���뢏�ӟ`��ʒדb;Y�	�cXc����ĩ��$�']̝��x����+McO��%�n?�)���'%��"��6��s6s�<9O��}������/�����_��}}���D¶�ƴmk9�M��rqK���x���㺜��u�i����r�>�����d1��neM�,IwD����r|%�����ɽ��@�Z�l�c�I168h�}�׍��x�.Q��Ò��$�Ac�Ž���^[��F���@�4���Pq�
��g]�b��sJ�jG���D.�Ҟ�A�Q��8@b�gbxU� �޼�6�⏾l^زc���TW�C^DW��'�&�,�3�1��=���>h��/"y>R|Q�pSm�)r�]q~��`'�9�$i����)�$�#Iô�`U�YI^4P����hG��8WU_Qrp�w�#t*�m��F��a'e����s��0��2E;rn�\��wE����vғ��0�K
N���<+|�F�E����:�-<�E����rťB���i�C-�+��X�<p.xݶ�p���U��8��&��ǲ�;;G��Q�Ô�w�2ƕ;_ɣ�+l�㘶�~�b��K�Z��fR�c6rl�Pk�R�lf\�-����}#s� χɠ�B���M\��$a:e��q���X�t,��&:�~:&?�i�?��ʫ]b��6��<��t��<�a�X����eѷ^�b�NJG�c>Ň�o6ݧ��ߔ�C����>dM`A�,2_��?�G߶�_e�/=��f�M}�m���.Wt��~�BW)�xp9�g�Qk��W��C�ځ,:��r�߷�?%�� c�|6�u\t��$t���"�Pj�*�`�[�;��Lmt0ј��-�ٱ����t�����_�<.p�Ob�Uu|ں*�b��N������&9��f�l�VY��h�2�K/�0���o�J֍��^��]9%�}zg|�ٝq[N�����:��ۦEwS���_x~�*'������|\����'r�x��%���]햳�����CE�wqG���T;|���G�I�Nu�g��~�%�1ٺtu\�~s\��̸��s�H�8W��a���{*��?��5���C�Kƭ}k��r�K��oYT�._��������fo��~�ݾ7>�����-��O��{^u��S���w��Y�&��8����8Eۏ�b�(�{�	qE�1X�
g�(5�_�>L�u�1�tG��H(�E?�8֢���h��i$I^)]��L�=���'�'� ?�_�S���j|��?3����ձWvW!��)�r�#���;�U,l��8�s�W��nb}F��dT�ޝ�U^�C���nz��
�uٖ�7��k8Y�ƍ�ߋg?��o�W��r��J�&���#F���>c�Ȱ���IRg�ŦvĀ`�0���=W_068M�P��^�8��ɧ^�i:������Ç�y�bO\F��ǯb���M����{��W;o9��J�3��M��&��
B���X!D��9N��W�r;#o-��S m�if�S;�g���3�A�����i�N$|`���c�<��d��=t���yj�F&<Ȇ��Oi�MY�P�N0��v���/������?â<�69�@�t�<�cDߌ�a�8������4��P���.�ב����d���Y$ox�3vb�B�4�v<
?u:�[����������Ù2�q@#�M�N�_�-�9��E�b^�|nkL;ә��OE����j��U��'��6J��j�c�N�#ǌwh���A����H7�ƥ?��#�J�9��W�H�9K����oKK��?����bx����[�1�".�̛7��fqZ88�杘�da+|ؕ���e)w4OIS�x{�&��`�qPzC�x�E�Mf�8M�;��j�����N��q�š�,�nu6��c���>�Z�(�᳣6�s"�u�W�"R���۹r�ĕUmX96o�ڤM�(q���q�����7^�cZ�������Y��7m�W_�}�.������8;^�
�/�q�\w&��>��N��zx��Y��C��V�GܮF*�:f<�w�+������ [r�^o���񕯾4.]ٴ�r�����\m��w���ܦ�ǒ1������즜��{^����������y��w�]>�,���/'k�P�k?{�-�������켍O�9]XCNC�@4�����t��˾Z��qA{"N4k/��	�+���+7���kc��%���@���DW[�����p�d<��̀�!�O����U,��~���k�<g�ɭ��/]���A��<˫�?�W�����=S������cBTl^c'm�L��R�Me��R��_Ŵ@cg�m�4V��K(3��ʪܑPy��_x�����|lb��i�<t��`��i,��W.E�+<&G?c���_�����~#�.�Z�uZ���0<a��|!{pʒ�<'%S�v������7)e�%��?�{��.NN��o�C���yA�p�S�Y����u%�g���r�.��?N������>�#'���~��]p��Q�:�#d0�7$�$s�W.�l�����ߊF
#�v�xX]���r6>��NWH�<�����U�8=��j�\'�����=g�1�j��I�T�3$v�����I8DM
�v�d�<^�A#�zd�����w�2I��A���dÈs��ӜY�,�y�Gں�y�	���;��1�V�ř��ZG{hE�E;��d�7���)C�͟Zgq�������u�ꗲy��bh��<���vS��M'���S�&������-��י�8n���U]����5���8Z���L����"8��<�GxH�'P5�%͂q����/�w�m'�<���رyZ�8�9����q{�S�y1}H?�"ƹ�_q�&ٸL��I�Q�Ҷt�b�XtՆ��З��z�b�u$L�;x��#�:�n��B��l���|�?��|�P~���b���p���w���5h��7�[D�*�y|ڹN�q�jQ��/�E<�Z�%16f��0�rljl/6.rQգ:�����r9 �tڐ�q%�"���(���y�Y�u�mn�u3J��7�0`�<|��WڃG0�3���Y�'���0���Ь��IQ6?Nì�"Kt����,2,�9_�N��A������	�)��Y]>+3��:��|���In_iO�l:ڹT
��.��}�K�8c��Ǖ!�yI{��M�k��!����=��9.ƫ�~m���k�矗ӳ�7�����?�}zo|�����;�kM?G�rL�Q��I�6T�F���t��Ҹ���q���q��{c��?q{Ҳ��#�4Y�ѥ�7��+�(m��i��7�]ϫ�ƺ�����H~}�#߾��±��>�����cCp+j$Cʕ+m�#>�s�:�w�ƃ����}^�~��oH�'�l��8Y��l!��\��u��u�&h��pogܻ_�j�ƞ����n�܇���ۉɸz�!��)uެ+%�f��x��3�0J��D_Ф=y�A{N���ʈ�#����p.�>(q��S��R� �m�'�O������F`�����_�s������w[�5m�M?��BdI42���'U��s6꿒�;��u��ylVթ��:%�o^��8�r����i��:N��r�$��d���.{N ��.�+�.�gn^/<w}<{Csm���d�/�w��%�q_���O���q��Ir�Ea��A6K<3��q��� $����,P4�L���+RJq��>�1��2�\����զ8>83\��w;�����١_�$�f��o-;���@=����3�<�o�r=�iq�Ou��b
���k[iý��XX�a��^\Tt4���W�^��:AC������nޔr&�Es��)�]��2���������@B�|����W�/z]�Y���e���a��5�Sc��q��?D�S(�8S�����_�9ж�e�l�V������ܩ&�<rΦ@��KE���?�/AS�jчÂוU׿�8�꼉����F��󳲂K[A���$�
�M�>6&Ĕ6J�����_�r����qsLQ0}ˈ�-Ʌ�\��ڻ	��&ѷM�����,��-�>It.�2��_�����t0�:��#Q��G�/�K3�/��:P�)p�e>!���l
NL�%�=/:�,Y8�|��\�ˍX`s�3'%Ԋq��-h�aR	�f�H*�\�Ne���1�wƈ�㠔@}`:�ʢ/�~S��Ѿں̠3y�@�'�AU	%7B�q"�h�s��~a�Ya�qLQ㥌���:�n� �7"U��8��)2�3e���}\���x��Y���DQV�ٶO�otʹ�-��� ���o��s?z�z&�6�krX�V�da����3M+��ߦvJ/���xᅯ��7n�x�o <�^�����>����g�V@ru��v���.��[�4���r��ޕ�u�פsg��D'<����)8Q[������E�6�OZ��sx�>��Z^�k�Ɩ�7`�P��_���h�N��_�|]N��q��u�]k���;��(|'C�:^�Ӈ�ŕ�ñϛ�%�%�n*#b)j^�v���/ظ~���)��yϴs� ����F{�Yh'�͟��/�� ��l]R�2�O��Xp�S�ǉ�G���"'!H'{	>yh�K�Ug>9.��7��_R���h��#�6[O���~Lx*��;��/��!m�c5M��*��rSp��Om;��;�|ɬ��|ް�|"�����t���=b����e�7�>����N��]�'wV�f�_��d����^�) n�iN�q���+���\/>��o��i�7�7�d}��9YG�h����iC1D:��n�)<O�_�A�Y	�q���8�!f�q;x���4�`q[�#��"�.��\�C��>��
u|��x%��
��8+�!×3�Y�p �Pd��ߩ�����-�8�^E�B�&����[(���ge �@[��
<J�ӖM�� �>s�14q��Ně�ƕ�\Ii>z�q[D�ڻ�qx*&J���	����҃�oj��q���:(#�2�ɉ	L"ʻ�x8���bp�C��q�Ć� у��9��z�9N�S�E�"�L����,Iո�'���-=ݦ�<f�L'1�h�f�����f }�c�}<4��hByڠgԇ:�{��ϱu�ʽ��9��'�"?�g� O���ɃG��vD�s������x]U���Ŭ�-i>�8Ƭ���i�<��c��)��!Y�x�M��V>�]����[�?�+�X�~�x_�㟶?v6i�e)벘K�缃` T�S�rJ|�a�?��EYs"���,T��[zzb�m�o��Ġǰ�:�\�Bꊮ�+�̙c��ү�q{EW�4�Mj8�"熤=y�V��U��0I�aB��*p�j��g�v�|Cy��0��@;/Z�@�\R��"yW��DA�|PTQ�&	W	�T7��3Ǆ\i~<L=�]�x�h����=��uSze����+(��|s �TQ��y�w���.�K���"�����k󒜫��g��}�fMľ�"�r��޿�����-?��w�����\�V`l��9X��n�Ϲ��}<x���F�^��w��*U9TK�|xE��1��OƮ���;��]����Y<7/���-<�6��]�Q��@���Nߦ�[���틧}h�1��X{'~d��L������d��� �,$��y��3r���y��0$0�w������d�8���8nZ,h�MÁ�1NN\����E�܆�0c?�&��<��D�@�`�����z�S�0��I䘺�:�8��=�����"p�M�r��,_ǿY���yjˠV�z�o�IS߲v^�����5ߦ����٫��L兿�z��8}>��&�4/\��8]M+�n�����k�/��E�G:f��M����W=Z �&)/��~��x��n�go^Q�q2V����+'������x���v9Y||N���_��Aӂ��y�6�~1�����#�i�͋��*�"�D�?B@������b�8;���Q�.6ikt&���7$��Țr�v<,�+Q��kV�sx�ӓ�^jl���Ɨ�팁�ʨ���sū��@��"�J0fM}��:ޔ��f��V}hq�2D��J4����&�yE�`ӸTR
/S�R�Q�nꬤn.V}GÀT�ɸ��)�T0v���?����HV� O����ܖq->������˺/a;��Y���tbߚ�f� �
��c��gB�(��T��D���.7�����eg���,?�i������U.2������h��:P\s�?�dD��G�t�S�@j�h��� ih�`�E["�x�6�J��7����	��ױ��O��[����k�%�����r��1I9�V�)g�8�/2��d��"4���<���͘P���9�	�*��,lw��嬷FHc}�$'�:����g�M�J�7��1�z��o�:N�Y豢�6�"5)`��2va#0��J|�<�%d�O���o���n�L��S~�+2����~�~N|9���@�ᄁT2�����\�&���S�^�Ge���$@I�i�/���A�bo��+?;���TC�+X8X,����!��A�c��YVm�����q�*�?��m]��:�U�%9Y���r����,��8��ǘ���݇{c�������m>�.'K��������}�Ev�U�7�������rXv��.�*�xB9f|�W^�ڎ�rL�9e�l�绸:F�/:8O;{8Q���Pq��!�:��E�g���s����X2C%V�L<���5IJ����֖�Лr�nz��>���p����{�s$1/$�����!{B�*��g��NSI�u��D�;���c#ud]�����A��9.P�iꦴ�IÓ���h�w�Q�\Ĵ�E~g����]NY
���e���Ƞ��8y�U]S���SG:�a>&5nD���	�������pMx:Vy�J{E�W�����Wo��<~��Č�۾p%����U{����d�a��|���r���:.�i���,����O����t�����Ƿw���8Y�'�W4)�,B"��-�,t�o�����+G�&�$�2���"���a�4Õ.om��W�	c'�q�\�����l	�GF��;G�1ΐ��Z����o������ܴ3�t�H�,�G�Rʨ��"�����/��[ҟ:&�J ah�2�2+0c���v����M<�2L6+�8߄j��7$r�#����P��b�
.3.Q(�%��"�� J�R����]�����Gd��J-o��O�V�c5�\X��Nїt��(X�yd
�&���]�0��s܆2u���gA�N�4)xʴ! h�M!gk�@���d�S��p����4��`���w�w8�����q�"t܍e{�ܭ9NY��A�_��vq��mV
݇%�3�컩N��O�#����|�@���ei�<s� �SP�ǝ*�Ê��4�*���,j�:&��9?T�J�,`��1m��ץ��/�_�d�_w����Y�$�GY��*w3`ט��ukj]�����y�\�v�<�.P���x֧d2�?vz�AM��z�q^>.��av�Y�]��0����2���ՕR涴R���FP�Sp5PT��N��%���g��|�	�!kCZ�^���D��+M&|�a�o����`{5�%yb@﻾q}p{S>/���^��s�<;�xt|0���u�Ɍ���x�m�D!Ĭ����=�c/�/9�����\o������x�o��_z��`_Nʻ?������{��g��+9@�����ߨ��e���I�>}��T�8��O+޴f������رgI��ƈ��#�T�{�:F�,e��h�9�99r,U�]�p��cOsuWΑ�EH���}ߺ_H��GR��.n��.�����͛�7�o~�[���~��@x�<�}����~���?x����timS�-�0�M��я��ny=0������gC䒚\Rd��NC[�c��¥\�dNJyo��"m-��$���R�C�|�Y��.s9U�r;�KY�,�j�:l�*�|��� _��Z.����WiX��ǎ��/���`�������*ؖ�,��4�pP@��JC��$�� Sxt��S������Q�x9�v��	�04�WD4�W�kz��`\�G���ώ�������_��������XU�ʿ�w����Ƿ����p�D� $�V�$ZM~�Mw�X䪍2rX�&s&��H���,[q���,Q0��|)$1�ШY S��a՞��(���
]^9� ����=l%u�R�(y  5t���� 댂�-��ƫ@�?>R�φ�n��+z�K����W������p�5q'�d`b`�lG"�2��F�\�AV�`n~8����v�:/��10��s(;���L��c�{Z�CM�Q4Uny���͋�������y\L��w޴�y[D�Fp�>�mH#�E_R>ɴe_JZn��'OG�}�o&G�sOe.�6�g~�l����A�se�{Ӗ�fE/�B�1�/�#��'}e�/I)3��N�zn�_U �Q�W~
��s1� '���[�C��n+xEڧ����δ	3�+v�|�5�.VX�#6� ��d�~�SJ6i�_}>Ï �~(�]�%1�nK��7��筮������t�:�g�F�~^ޱ�����F�
՟��`f�Rn���4�ɘ&��+ɧ<2��Tb�u�6��^�_�g��7tE�	�Y��.��n�X�l�R�d�w�g�N�k���[4+����S`������8��^y���30�S*�~�����Z_\_崩c��r%*��e��N)�L3|dC����3C���X]W��nl��_zn���W�׾�Ҹ~���<���f��������g�����nmx}���|��z��ߖ��2�	�9�X�3 {�~*'+k|[��]�s��U?�=�3.���tx�cXK�&��G���y�0�.�qL{�+��?0^�K��Kg����0.*^�xi\ں8����(���`� Y\�ta<������ύu���%]�ap�޽���k���I^�!��!��i[��k	��L���(��>j�E�T��kY��<%P���|�!X�M��GƂu���i ����M8��:�*&�u���R�Y�'���6�
�+�+�:g���o���L�U[���С�k��\���94��o:W^�&ڳ�.;�_��t�:��>���}��c+��=��.����V˸t����ѿ�a�9� ��7$o����W/���6�����̍+c��CK������O��'�'��l|t{<<�S[�p��.�d=�� �P��K�|�x���GJ��%�T"��3g�UM<΀JY8����3�Rh9��7�	�׬f"`%�C}�M5�c�����\]��C>��vn)��r���%
��HВ��Ư~!�� J��_��y]5g�08(�ԛ��^/"ŷ�1��?��9�E0����S��x�Q0>��M�~.�mO ��P�5ȗ�[�/���$�Wa����U��>�s�tfe�|IV�>��Lْ��I���tN5� S����r����W���KNK@
g�)��nG:����ժa�#D��}���	�v�VY�Tm'�Nܼx�?;�.���՟���~t�L�u@���ӊ�)
���&����V[_�(�&|���l�XJ��'�y�	�I��ւO������������W0c��%���ᰒ����VO��</���Ο���@x�7/n������e��4���w� t��%�ll� �y ��y�	<����[[���y�}����C�YxIJ8ߖ@=�z}�1v����=��v8՛|cH�&�n�9��Ō�4na����������8��wl8V��,�S8?^��́R�E��hH#�hZg���w_����+�Ú��9i	&ڠo�v\���$���Y¾P,�T׏���d��w����W/�w~����?���w�;��q�]���O��������x�������������B�9j�r>�������/���v���LV�~�4�ֱn�풜��/���Ȃoimo�w����xr�����2���-G䆃���ф��Mˉ�Jw��l?ؑ�v�� XN�l�Y�#G���5�r�x�aw�����HV�����x����կ}m�����¥���8�l��~4~����O>��d=Z���,�0x,��)�E��q��>=����A�r��jۤ��z�,*T�?�u�n�0��zk�JȤ��� ��/~&L�'�� �&���ڠH��G2���5�N:�Ƅ��ph��� ���2	��a�y��g:�ӯQ��qҴ;�ȟ��Ep��ߢ��m}�1u��0�,)�zd��5�D����ӕ�Ib�v�+�k��[�P����q�����W���֫��}}|�ǵ�G������O�ǿ������;{r��tYN��OΖ��j���揎ʉ��r�gCe�����k��`9�N�ϊ�VA& f��z���%��c��K��r�Q 󒆔��E�B'h^1�����ЄFxAb;g����d`3��y��h~Ń���	F���D�)�rW��ړK�����?�B��W�J��S���b������T�z�3=6�0�$�DBpѧ:�4����ݜH;�����64����8���x�<?�s	���`a���)'��b�~U�S�8sL�����I����O����j�q��鋿�5)1�i��u>h*�e���&���x�b4����7�dq����"$��su	�ש�r;�7�O
FR�H��Kvq���XҒ?�F�{�	+�h�o��w"4��Z��8h�L�g�g�8�;t~ކ�m9J��Xp���'�.��00����꧅�je�flR�fA6x��q���	{ز���oل�!6�wT�y�</mL�z0K�?/�J��r����N�6��T�6�-i�!8A��D�Ҝ<�f�Q�ƌ����}��֡��S��鹤�ՠa�Jְ,2.�Ԇ� ��S��n�1<�GE��|�_�^����p��M>}\:�����|"�1(~��m�*��������'�z(p�&ѳҸ\G�i�r2Tq��j���u�+g�Ѹq���� '���;�k<��E񠽕����[�xK���ag簾	�8��ձ%kkK΋�<������;�u�:�|����J�8H�.]��dў��c��ѹ'�osݗ������i����lh>�9IE����������4x���(yi���憜A�%9V����Z�c��>�;�����`W<.�k[��Ƶ���͛���u��?������d������ؖ�w�NV�e��ǉ���.Vd&$��ӂ��I�2���?v�(C�(���`=h50Lڷ>ц��XZJäm���h�����`�U��^�R���9.W��m
�������ǆ��;� ]�����>��s6���|�ڀ3Z17syp���E���)/�*�J�\��
����8�ha����,���)�i���@~N����s�]�^o�����~:V�,����'���??~��������PH�/���gƱ�c+&W���(n���D�Ï\����UL7w*gk���5�o���9��YLa���� ��k�*���A�&������TQӱyPF�q8PX�\)�%���4���p�*GFv�2�VV�隠�	a��IQ&�ӁSI�`	�&�YGa@]%<�ПT����	R�ΓN�Z����R)|�Q���u�T���3��;���T�Z<�Q��w��/��
_21�
�>�f��CF^��7O���+Y��ߓ�pLhʙ-ޝ&ÿ)բ�|��*d�`Z6��|?-t��s�`ն[��c��5�;��6��~�!�؛wGMe^Β�l0�^T�AE��p�` 
Z���|�����yȼK޺R��O)]�]��yY,�$�D�a�w��Np�s�_�]�ɌF|�,��b�ua�|R��}�q#��Y��eay�1�fD��,�p��!9����� ��6��3p|����=S�����"h^斾�A�:��E�����R���X��Q�_�n�O8�※0�=�s=�2of���;oJN�x�;�擂93jd��BIp�:fy�n^��}X��)u.�g�K��Q4���Ē*ɷ�9�H7\Grb1 �D�K�Ӟ�����v��Q�F
>)I{�LΓ?u�g̹�;u��ܶ漜��e9!\��S~�g��>~�����o���[�g����f������#9+�Q���P�Y����������exӞI��-�@��4G|ƅ+sq�p�p�p��^�0��(�~��q5���EPm;�1���c����������} ��y!Gi.�j��"+��o�>U�=_�;�y|���qq��w���4�f�_��}4~���`}_�ት��q"��5������#�%_ډ���7PY�*��-���ᬙ�+�E0���n�s��r��9�1��T�c_9Kl��2.��+O��n�_�T�C�p �y�m\��
j�6�Q Ge;�[�χ9��kJS�xT��o��E�a��sMSѿ"�2��P�#�G��)~���p3AuI����r�ێӞ���<lr�[k?����v�5���<;���W�d�6�|5W�xnk������r�>�|w���ZZ���z�N��� ��,,1aG�\)bF��:����J��, ;���7�X t�����,�
t�"��.I��q�=��r	���%��
�g���Ф̡`:����" :$ �/&0b��1f�Y�&by)����-�=u�2�N>�Y�?���ɫ�,sH94jVF��>��:����І�؆�N�x�����O���nB�*�\84���H��-T���QB�N�O����R'�B��/�n|,,-�Ç�2�3�j}9K�I��/�U[~jj�$c����ڌ��҂q��EL�>v�S�x��Z��eF _�l\��8�3���}�<���0�-Hΰs���cڳH��P4��� �,�Ei���#�*�?��\\�t�Ϯ�f]���k|8Yѭ����ŏ�$�O
�+[�fi� o�S����ҼЈvӱC^�p>�9~签(,����\��8TfEylL�X�_�SF�teB�Ŗ�$��co	����"'�sޑ��}}�?��7@��}D�OA�U-�܈�� 8c ���5/}(�E�H3!�M7��:�-	^�M��͂�:� �p��JH݉�����g�k]"L��VkA#�i��ȭU��:�8�oo��r�sۮ�?��#s�k�?�_�@g�?��8��or��g(2��*p5�I���Y���٧}9+���\}o������^���9('�`�R!Om�xC1o�;�i?�ŭ{p5��P�?��Z����se�6��|�!|^�m�~��7��1�x�#p�������(�8�8nȁor�����}9W8��ŧ/|�^�}����X����#Ϛ���u���͊8X�G�����͡�s"�@���9tD�Ï>�����;��Ԩ-���*�� 42�o�d�m��c�w�?�-8(�`ֽ'���RyX���uv,g,ㄞ�S��y# &:|ȱ���@�|�_��B�J��6(]ßch�@{����g	�"�3dυ�y&�?l��vfe��vm�s�mB���d:�]�oR��OL�G����K"�|�=�4G4L���lh����6<kG�L�I�S�����`/&=?���6�ƫ/>3�����;��J���-�/.F�_�d�������O�㕱�vq�+".'KʳY�7��a�+n��L����Q����1�Գ��:�y�|C��de����S��pX)svC��N�����럅�&զ�����5,����f�<�wy�ɤ1n��F�E��;��&[Ǔ�����uB��g��pz=��xz3 ���lb����ma,&j�&����6��A^Ԟ`��I4=�T���z��d� �YtL^?�h�p�(h2�eZ�u�	T��r�P̗�O563�օ�`#ڡ����q�Xw֨�7�BwF[��1i�_�0m�+͘S���z��~+�-�)o�b�Vc��� �@ӏ>&=���I�*�/(��8�?p9�,61�g���UI��}.�����"�QX
ɻ.�:߸�{�+�B���p��J��o���k�Y��]������9o-�N�d9[t���ِU�I5n�@�D��[h[�f����x��kوA3W
b?�!�m$P�}��#h��n5?�tXY��l�!����=�ѣѴ�<m�� �4�X��Am&{�*St{�9������fcΊG�b��޲�L�ڡ�:P����馋`8@��J�6;O��6;�ڐ!��	��/�~�sA��'���a=���w��>�mk�R�Zx���݆d�h��y��n�<6n���bK�.�����ñ�iMA;�(<c�(�Ӿ�Fb�J���-�K��o|}���������_�S�����K��d������|ȉҚ���q��%����\}:::�		���;�a�,�Y,�G幢%�Ģ?Ec�
���y$���r��絶��;��\ܒ�'5@��Hy�g��M��[<��}��꺯�mml�59Y�Y��C�	�q��+l48������i�g���>�@�=T�{�O>�t|$G���ñ_/U;=�x�U��x�Ы\_2�э���_Nxg|cĪA9�#=j6(�*XK])Nk� �̅�N����n� X�c�(Be�K��,��O�q�MY@esq��ϖ��=G.�Pl�f[[��Ͳ9vP��F�Ce*_,(,�p���`l�9\b�����,6� f����y�8��|껦Y��:��s�nl��L�9M�:*E��U�u9Yk\땽:��ue}e�����7�d}[N��/��g���?��O������{'+ce�:yQfɯ���,���@ib�y��|y��6Xl>r[!p��C�
U�\@$Y���c����1��˙�ꨢ�o�*L���lX�(��Br��*��ˠ�,1� a�V:_8�Ҧ���|������Z
�ȫ_9�ę�-Z�=���h��+�EV-��p(@C�����t2�_���
U�)�g�ܼ��N��C?�R��T<d�h�O�JXxj��PL�]���j�h�pQ�>2�4Ѧ̓�&#44l�ou�|Ne��c�̢�%�Z�C��~��L�Z&Ф��,s.���p�1���,��3�:8��z��8+t_����T�'C�����۬觛ў���q�,��`��*��,�e��q��)����+O)���&���Τ`����Ŝ~4�y�I۶$�, ��:G��&}'�qE�:�`�8[4<-x'|q���>��<��1�T�n�dq�J6����ɮ���ݩ<؇�Y�� :U��9������$���
�d�}d���x&[�H]3�<R�i�C��
���9&��Rvn_lHi�F������w6��|��A�k�� ��b�����#o�[���и��/����~��RJ�s�Y�i|{v�8<�4��ۺ�-�u��Ј'�JT%p�~J��6T;Y�?'rOlWi^x����ko�����x��Ab����ʜ��Ϸ��=�e���ڵk㒜,���+�#��9�axQf,��S�����g@_��|�����abADV��ɺ�+���U�܊�k�=.�[����q�����-�����AP�Ct�/�0qb�����};~���NR�A�Ǻ��������{��x��5D>����4���ɂ��P�t�����ֽi��EV�~
�u˺RP�SPc\m��~F!�_R����رZ�b�ȉ'z0T����#�|�R��a�ź����Xh��âl>?�_������	��o��3�ٱ[wm+5��W(�x���K�5�8m�B��n���(�a�K�q��qΞ��}�����"Rdg'_����ԺI�<�=������8�ߓ��:���M����o�6������UY�������������s9Y�+cu��0]�$�Kc*���Y��'�I��M�o&5qb�)�	�V��.�q�,�M��7�RN�[��D�X:�N�g�i�0H�UQxH���@>2��J�x, ٢�A��Ԋt._r6l6�.����(�p�~?��D�T|�B�r}͞'���>��� tx�+F�+l�hac���I;����S��j��5����Ə <��g�X���OƏ&�ar8��\�?S@�}�(��X?��3�=��k�2�TѼ�ld��Zf]��y���r�Ò��U���1n��ٿ�\94�5�l��tI�,�'������ ����^6o��^ ��mY�BA<�[-�#��q��V[�W0�dI�q��l�73g������۷�I���DY��AӬH���Y���'�l>4=�� {��2���%�!)�穊�b�mXl��O����/�pN!������E�+|�S�8��ۥ�$�bAv��?�K�x1,��k�UD$�b����x��@����<�q7���q��GM�)�E�
R&=�gp�@�\U]R���0��V�FhA�o���Mt���v�D;aj羹�
���H�*���u�p?��;`<b�����	Gl-��g��_h��Ww�Q�4�<���]��R�#��B�U��t]9�Xm䴬��}�d���Y�8����x���^׺�한�&�̡������k�'��X�p·�	��>ɛ���~p��W�4�p��_W�^�qaqp�ձ\�y�#E��3��է59iu���8by����"&
�V�P?%��|�¥q��󱦹͉&�"�/�@^����[n)�Ϸi�5>��cU�/K��^���߱��D��Z��rVx����0�9o�����S�w w�u�E5m�?5b]��J<Ԟ�rNئ�!Z[��~m�y��g���z`(\���s�@4O��ʩ\��20! 3k��?�+٠+9�C�i�O�����b'��!��"s�?7�7~��_u�E3����g�%�R�Z=�KK�t���E�Ts��~�KDuTr��P ]�`���a�Q��gR;Y�hU):a�Dr�F`GT��Hi��S͵+�k����z���o�j'뙫�¡������d�ݏ�?��������,����藅"N��2V&6lB�p�&�9dn("k�#�ߜ[(p�xY'ؘ��u"���f�1�*Vd"��J�(MPDq�c2*� 4���dBؖ���\����̸���
�c=)4�]px2) ��|�����H���M���-�~�N1�9c���!<B�G9�L�_>f�$�x�+pV��<�C��1��׶L�u��oU�&iz(Ppk��#/��@g�B<��\��"WI�TnG��?�b���Pc
����������hw0��0w��w�/����1��p���!x��J������eB��̝�i�`���(/Z�9lH#�f+u�&�D��:.^�ݦq�K}�q�*��풂����aI�t\F�Ap�v;؞�̓���xe��1/����_����>� +M���X�OB���C����2��m��(��q��϶Kݖ4�Ŀ�E�US6=x��3�7��)�y���ͅp�2~S�a*p���)/��%/6��dX}�" ������ly�e\l�8���q����E#7�1��-|zs/�V���s�w���v9[�>e�\l&;��W��P�?6��5߉���H��)�U��͏6¶�с�z��ϡx��Wl�uЁ�mv� �T:��¥t�[�Y�E���-�P����k������9���&r�w�]銊eB�ˉ�y:�6!��3���o=����1�2���z�v0����Ɛ����E���� ���u�M*Ư_�L+��]z��ċabY��ƕ������x���͍r�����>�D�)[Ӝ]����Uy
����?l|�qN8A�[���/�`��G��9���؃�|o�H9d��5������5?R ]pB�s�1���ǀ����g�$.�_���.�q[n�?�3�s�7�<�'K;BH�s%�X�Wyջ��v�CsE��Ǽ��[~�U�#��1Y��b0�rzdoJt�	!����Z�3��]C��`�ԮK=�s�u&%�VnF��������g������"7�<�A`:�y�ߝ7~殁5H���8����6��{)�y߅�h�����������P$� �}����	�S랢(����H�q�8.`���f��u�s�Ɵ���J�d/�m��"��c�e_��H;��2�v�����G����5�ln����1���K��xu���W�s�������7�7�����_�?>�uo��=҄X�k�`��U����R&/.(x��M�#���� ��a!ӄđXՄף�185��N�
 �fӂ $T+q"��bL�C����Y�	\�8Szx˙$�C��z�w#E�%X�C�o�6	k���S9C~��R_���t�n?њ�Ù��2y�^@�6#S66�ڸ���mB��MI�67�u���%�\�cx1|��	����+q��m��!�u}B��g��U�@
�2@����&��������t/`��3z�TS�0=N�C��x��C��;�3#C��	�����o��hA��/A����p�g��xbr3qe��e6��/�n�W�)���*t��'�I���V7_��<U\^=�7�s��.��D��?!d
��a�Yass�MЩ���s��Ն�f��$�.dlX�b+̫R�j�u�nL!u	�5p��1�Fʠ�Q,��d�}�vt;4B�2����|�>�l��|�p��و���1��z�kd�2[���'�.��-��HAl:��Ycs�G�)K���}~�A�\B��ܙ%4b��vExS�����q~f�|L{�VK�1B������g��_�BJ�ЖR�����D^a�:�_�i�7O�<<������~�h��D�7e�Mx�-�r�)'��~{#���1��~g��/��n�3��释���;$�ol��$����ĳ�^ѺUo�֥�
Ӹɷ�H{G�B<�c�Y��P��y9_�9}V>�@�a�QRh#��+R��C��|5��W���p,'��ŞH�8���N�Ud<�r"'z��(1�����?�8#�n������#~��oo��v�
.��\��!�],�ϼ"�Ex���q\CwU�*���@w������L�]�_ߔ�m(�aU�z��%�����5�ٕ>��|�0:n�XS�7��#�]� ��[���$����F?�=���(���������?��w���tJt�Kn�S%x�s��H6������τo1>��3�#�y��		�s��?��D���	�ٷ�<vD���|W_�[��8d1M��:�Z��e��t!��o��M��<<��!�x���L��ot���ux��� ���?�)>�pj��`:&|��Z�;�S�����`A'Q�V��.H�1���j�5N2��_\_/ܼ:^�����^/�xs<{ucl�����?�������{���>�7���㥱�h˛3^�cH�0JQ��ґJ1��o�l�M��)�>�%E�[1% /:?��N��F`Q
el��<�x�5�MQ`x��#
��7���az�%�3!�QD·�0��<�&@U���^DTJ�äk���u�O��G����
�0�G�)�Q<���_<�+�R�@�H>t%'�A��|��˾e�/�3)�e�3j����;~O?�O��MF�������/] ж��̏�:��t;��3��7S�d6��Ld�GK�􏤫�G~E�y;E�EV���
@z�6+֟�w�ll���Ɓ��lv��U%
�۰��3�S�a�1'� -c�[/b�}&Q`C ��Շ�����'�q��46mx����!˪ٌ�uP16���x.�Ԯn]�!�ȡI<���λ-�v��q1�=�7��вlZ�u�yD친gQM[@n�cCc��_��*�=E��N�|��i$�18V9��I���ޘDƑ5,�1-ٵ��?���������gr�aL��R¢�Ƙ�:�h��%>��ƥ|�h�&��c�Yi���3�Kt����6��^���e@T��y/����$��'��_�hQ�:�72B�}�-�pS���aݩ���5ڭ���lxl��h*�.�w��A~���\m ��"*��38�дY؆.+Z^ү�L?����T�9ɉO�%�5��>Rh�K�٠
��-Ap�-o~YQ}1�n?ۘ��͛"8O�/�9V�4��9,^&I�~N�I>p�:�5n����.�c3�W	���Țg���[�pQ6j�����> <��R5����F ��-�!z���-ݾ�g�Pp炯�s[���z�b�0���+��ˑ�a!�:>���LmV4~k��^�2���|$������܁�r";�D�e����֘�#`�S�sR5�W��M�ãmH�+2���[q,}{ج,2D��2"o~�!F����;n�n�<p�E�1��m�A�l�K��/d�1��$*����M^���C�r���+��b�>V�g�u�ՁW�U'�4�q�|x�V�3�Up����<�`$'�,�R�ܯ�jn��/�`Ψ>��|b�ɾ��I��Q�s��s���R�M0����5��Yk��G�4�����+.m��GG��0�J��-�y��x���/=;��yyܸ�66W��/������?�7>��ḿ�Q��M�rE,��@�N�s�'߁K���8rݛ��<�D�yC�y��jE���6�^�l�
N�8R�KK`I�;?�a��4��
�G)��IcV]��x������G�\DB�D6��j�����V*6�
�OT�5�=�S�!}��u-���j�G���	����q��%��-;�㒜,����u-VG'kg�y&�DO���D=�=��Ȩy���o�2�=Z'T��};�9#�K�,ڒ{�e�3��7|qLy�H�&zo��3�J�@������.�G?*_��ֵ)h�}�<k���M�$��`YFo���[���I��
�wѲ�R���1b�<��.՜�|@G��F�t����­!1���Z�k�
+ڔ�(�}�쉞l�8�'.{<�x,/�]�xQ����ih�~�����em9+u>s;����4z��^H�/��2B����?g������j�z�1:e��b,�&�B��-�fht�����l}3O�H0�·�ʷs�8��#��=r %4ݖ��JW��ȼ���w�5��ʢSyxA'��I��8�������~����k3��۶�	�bƒ���jX��m6���K���[��_Dt��%��]��:��.�)F�i 5�f,Jv�!��=���z̩����`����<�c"�A��=���e��DB�gB�V�L��}mjx�_�lZ��L��3�>,��z"���m��b\�3�/�7r�':}i|ޠPVcO=|2n�,�	���ho�} ���9�[{d�*o����<�6=q�v���hɛJ6���=�v�-���v�_��v_TB�q�o�d\y]��˽��U�8�-sR�q�D�ވ�=��4ߤ�����N{,��T��7B�3W�ދ�g�Kp.�=O����1~��//kܴN�zD�-������"��(S���X�m;q��C0�vΥ�*�VNk�t��PD/\���k����q2�-���ïB�%����z:rl�E���'� �z�M2�:Yfy�_�H̉w:�ȑ �ÿړ���h���%؋��J��̯��xe^Ԝ�~�S�>��!�ܐ��=��=~�:8�)�/J>s:����=4�d��Dh�y�5>�]�����O�1��[JȨ��/�+R��z�;�����ɘf>J>J9�<с8���7��Q���|�A�[�|�bNֺ`.m���W��ͫ��K�����؀仟}xzo�`�{x0����=���q0.�156�C9-�Z��;@X�1���#P�t��a�N��)�p�'��erB�3������$U�h>E������h&(g���i��{�$V61M��i�>��r�W��a/J�gO���(�eC;E���r�<T֯T%�#}<�#�	,9d�Daul�+l�~\�{�c��zFh�93�(������M�<Μݬ�h�.x�a<0���(g�x w�Y�k�2��hY(�1F ���1���1����O�[B�1���Sqc�1��Go�C��?&�#�o�ɥ}��M}�y�d��R2t�����q ���3/�G��=ϕn/z��u��;c��I/�'�d����J�NV�ܑ/Y)89���,�Ȉ�|<���d"��-S����W4,����_��#�w��7�>b#�f��|��[<���"{�'|����*��`,2Ф��+x�Y:�>�|!��m����x���2��%OZ��/�����~���]��\ߚday E��i���ѯu>	ֻ��������&�2<�7��t�I wd >�b,��D����!W
�p��E���k�M��с>�~��:�m�f0F�������f��xG��U^x ���%:�.t7��?ƂE���9f�� �ś݈�0�#�Q��mgl,}C2����9C�^5���ec}�gc�pk���%.��?t����'��[�43_�l(�&�tK�<���E��Ilz���m�h{��'dLh��޷��X@÷�-RƆ6�c���/dxĖ�V�7���	p�)�fV8���7S�!��n^Ӧȫ�@�r;�|�_��3��;r�k��'����c���1�h�l��6���o�k!N���_���6��/N�`g���|C
G|��3�'�{+�*G_������6�|��N��`yhM<<GX��9�V	��Q8,��?l#��Oe���t�l�_S���Sƃ����2.Y��"��UPt�)�x����e�o\Yct���?x�sU��#����D��Ӳ�`���� �xaM����2λN�#c����.`�$�10����h}4rS?-Ҷ�*��Gx�e�mmm���u���p�|[��\y�f�׼�b�}'L�aۆ�M�_��'}���n����~�]�l��B�s"/�2{��ƈ]���<�o2��?�g=�ßS�	��G�&;����Oe�xp_듈\UL�G�M$2����5q p7�z${�^�9>�9N֪�p��r��Ƴ�����,ۙ��>?=R��&x(�s|"ú�����",f�YXt��8bR��XJr� DAGK
�((�Ĥ �IfC���T6��'bXr�R��"(Z�X�y3O���*�R4@{ԽY� ,6Kve,��k����Rf���^���8� � n/�2�8Ub�ƾi�P ;��`�B��bSJ�C�D��_%Z=��<d��l9+��/��d�C�3�����������#�}�E�V>�K���&)Hy�I�9년6����d�/�i��:(Rs�t�Xx�$!��3m��x3�%*Oh���jh�@;'��2�al����+}��?��h!W�|��m�i(�g��Ȋ͆���]�d��W���\�f�� �!anyc'��1�h�:l#C�_����K�f:���仯�\���hxs��"?�@�n��1�N1b�ਟ_< ��_/oҒ��^���x����6��Y���7��@6H譮e�8�8���#޼8����~U�:����$O�����+N�O�2^w�h�	�����G7�#6]��C�l&cK�|A&ՖH@��d0�S2�E�|���D>��f�1��|�#㢟��/�t��g��f��S�\e��$|�r�ƃ��Ц7�Z�LD��l��DJ[6<�F�o�p볯@�~á3Ȏy��h,�3��]��������6�骊tS�c�/l^l^Z@�?o��g����Ϟ�$Q��Fg�ɤ��`��m�� u���U�ԛ�I�Ad�8/6U����g-��?r�զ��U<�2�L_���#o���l����,t� mZ#�x�I~�A?��y��c�z5r�ʱ��A��tr�uF{�5�)yd
�5;C�$" t��H:L{������,2᭚G�8���獃}+�y�56���-���P�[�'��6`v�v}�����~��H�5��� �,i��/6�I[h���_��-鎃:O̕i-+�|Z�+[G%_e�gFQ�RҺI?�'��N��g�f=S�]�ߞ{�>Zч.o��:
owG��=O�u�l�p[�Dt�X�>: l�@�r��|�;���{�^/��#A��3<�qꜼV{ᇿ�����k���z��u��J�E�Ӯ�ĮfMk���p���iú���i�s�H���ʩ�1�>���h�]�v�ት`a/���^�g�&���.v�k(z >x>"G��V��I�D��>S�L�]���������S���܉�˻��࡞�1P�8��3mlHҟ5pwoS?��_�ck��؀��Gw�[r��d�p5gC~���6�i{>��heP�p�D0�Y0�%H�&�Z�,���|�:-0pt�1�|��������g(<�8+�����Z���$^%<O�V�Pƀ���!CĈd���tg��`a������қ��M��&(^�;&X���˞�aR6��ń<}�B3��ո:G�2���svWN�6�0�� x�
Oh��q�H";��X+���7<�9�/�q�L�qoX�EM�,�(���H��n��/��u%��>+/���<�	���j9����T9�����������_4(�`�#��2 �M�?]�(ﾐ"��7O�?��IAo�o�K����hdQ�dU򥝆�|^muh^�WE��*�cK
������.�������6(v6��w�$Ѓ�y�`�v���"|�+�*zary�[���q(���s��o2��od�F�i)�e�O_����� �:/X .��n�#2���G��5�lBX`ៀ�����G[���Sc�g=��1�C�����V���	2~�"�h9�/���R1��ȀL��$�Tx�z�I[p���"����3���Ûa��H[���c�`�	�3�L+AN&1�ឹ{b;kܢ����'r�
��;��aiC{����sA��/����3����考�Φz��1�Ǒ�[vD �6���4ԩ����~��dS;��g��	x�чvn-���l � �6�hF���^w%#�����ӫغ���X��y�]N��?�t;t_�w�+�X�Wu�Z��e�y�(�	�1%E'|r�lx���y꓍�	���o�Ѽ)B�qaް��ae��|<9�dj�e���J?�Wx5[�gA�'|�Y��ʨ��*v���__���ʖ��F�#��C=�'|���ᾭh̵3�n�#�K-�G����^x.��h�)����"��~c�ʢ��Q��?��Y�u�e~�Ŷz��q���ؾCJQ�_Y��S�iz�Euk�]�I����q�q3H"�bzя�k�[7���m_l��[4���{8���ڻ��S|���'o��=�~1cI9|g>A����ʨkg�ˉ��o3���1ԽG���̏�"R����h''z�o����>�$�Z�8GE+VU�2G����d?���K����>Pc�.L'(�?��¥1��xE�<��@O��x|�_���?��z�5�aEy@��+h�.�2{5�r�͂o^h'Y��p��)�v�^il���X�X���$��B�F=g$�7��Xi�1�劏䜘����xMe�X��4A#&��`&t+o�y�yy�V��c�oew��D�i��(��`������:��gA"t����u�n@��DGȽD�PS;E��wN���q�R���L>W+��x������>0��yk���9���>�C�gC�������;�.qF��2��1Ƙ���@�����ч��G�o�Df�B���]�O�aA��}���6���1"х�,��	,]�l��i��j�e�_@&=A��Lq%��7>��O�U�š�3MN��?��1o�8��.��=��	��c�a
��VDuo�k�M������-���xY桎m�X�述��[�	L9Y��U㧎�����
��O����z�uMd��#/�I��<�O����`��/�*��k�p��^��?	R�7"V"��:����zAt����9�l�zB9a�W./-�0V`��q66:�s���:���r! 繆K��	��w6��B��f�ZR��Xpk~���а���`K�Lڵ��ג�e�|ϸLSsv�d#� k���ቡ=s҅r�C�Н�.������ +'��G Ȥm���Y�M���O�Jz�E�H"|��~�Z�y�B��#g~5���F���F��׭y=|3G�!�~ۜ�HĲ��2d���o@9Y�s�� ��y#��8>�x�cR�-d��."3_W�7g"�lZ����	�W�	v�xF�.��0��c�e��)�6�Q����DU]Im1.���<��tF����iJ�^���=�:�(]�O٘FN8!�EPi^X�%��M�dg�P�X[3�oP�9yz���-��1��͜b�!�^�?�f�t���[�C�Y�4��c�d~�>p'WX6��nH.~����x���n�'���P�ŋx�!�c����P2�=!֔e;W�ŕ-�&6�u��wd��S�e�5r�p(���M)��l`�;+z�zB�����_�{$�W�w�.y�:d'|��K=�k�n�u���#�H�9/h k�������f��C�[6D�CY�Il�i�.]���R�X�]��v�ē ��W�cYrq�<��6�f�:���j&�����c����n�4}˜�����}��c�۟��qa�H�2��zV<�-���"~�re�h�����5P0�I�}ʽ�=�;i@�K�eٙ����=��q|�A����G~f0&MJ���󆎜R�M)�R��	��Aah"k2�d�+>��Q��Z@��=a袨fL����BǄC��ݦ2�eR-Bpo��"���B�].�,��4�F�����u	�C� D�bؘ��Qt"Jτ̙�����}�ǹ| ��E;a&i�T�/Y&/�(�ό')9t�K�>�����D�Y�F$L8�G���LƌQx�.�Xɡ��~�c�D����{��d�.�̆e�,�#gj�-df���2a,s��t,������
�3�����X�:U��<!MJ�W)r/|�l��]�;+~a-4~����[b��*�ت����F ��}6T���F���Ü�r��yQ����\�g����/"��S��Ǥ�iƔ��U;�Sδ�_�$X�@���[���/�����4�p��z����+����4���}��]G>|Eg����n�g�lg1��������Kd�}�6K��4���r!�&8��ӷ,�#��:��^���%׾z���/��E\�g��`!���hz#Y8�A�����w��y��}�U��z2A?3��G�YF	�w�1�*�:���kF����~Ϻ�J6)�Ml,<Z�>�>�ZM���|Qr��&K������qd���p��D{���}�^�|�ʃR�p`��́�MY.z��!��64{�P��+�m}�6póu��g���P{���mb���k{�d��rx�J6�cPz
m�^^4LG�e�Q�9��w黢�V���"�M3�@���żP�^2���ʟ��1�Zȱ#�U:�&�q����M����GK�������1�x�_s��%=cC$<�����i^`SԿ�m�г!M�����.2ˍ3=Q�`���Ⱦ��v[�Oi ~�q�67�^6�`p[�96-����Ehp���5O��`�-���}%�W�X�V��
�'>���͵R���2�?k�u_��y�X��qA3�F�Di��ل}"x�=�ڢˌ�u�h>Яs����rX��m�ײҙ�(�XOgv��hV����C?�/Nʱ�s�a�'��e�x"�bH�e�ɑu;������_�r�ǌ/�l���
`��K�
���P���R��Ƞu�z��?d���ۛ��1��B�% �N�Gp��:�車J���}����m��1�k�V�,|D���8�Δ~��xְ�
Dȝ	�a�s��{,���@���7��?8�BEG�<3p`�L�c�C�B�SQy/K;W��5,&\��,�,0ìrf�Ǜ����P�/�Ջ ���|UX[���M$����Ai%���`�r�t,�s�����I
�����K��z=��^/b( �8�q�Ͱ�[
`Y���~({�<�zQ���^;�3gR>��$)y�ՆA<�Hl�� �ᣃ����&:�����3\����4�c):=x��#�'�M�V��b�4p��A˭ld{C�$�����`���@��J��2!��	�mZ���z;�d�����?�<_j������T��)4<��p���Һ�E�3rDn�#bX�;�2�3�韣��,^6x�d!���<����6�2�4���[���d���I_"�INȡƋ[B�ǖq!*���Op�����mz1 �cxQ�q?䗫�-����Y��LQ
N��Qn��L��"�����*bl3�fX����J�}��>�'^����f�k�c�x��gy�\D�K5�q��u?���E&/�,��//�]���K��MX�*6�4������qm'�cpz�;�@��ü]/�����c;Y���%�:��ʌC��/�r||�s��E`�T"��n�[�v�85������C;�-�fZ��/�y_���8Pf=����ӗ9?�D�<t�������:p�ò�� 3�ןC�E.��͸��t���cH�eAJdnK��;����n}?��ž�C(��q�WxFo��85�7N�1�^�Kv�#�f�辥��'+W�Q��9�`9ÏR�0M`�O�<d��7B܊n���Z�6��6�)��6��:�G��>9ya�m����d	?�D@il'��8Y�6V���O�&c�]��2�Q��q�S�j��C��ɷ�����H�3����NlYO���t�l鱟}}Ʉ��8�~)���P�����"�*���L�#���zƦl�ʭ�e��n<��S�U`���.{����k����ں?�?��86�x]�u��,�5��	�tQ�Vd�]��~ ��6W��[�	8�Ƽ "W��=�v�j�ã�������y��u��L�CtT�:~;Y�	���uxs�ڪ���B�ս�,S�'m�)��x��3'�Iଯ��0�W[��'B�,�
���*�b�Y덎�����bl�j^@�2a�(���ef}G��+��.�>2nk���^d'Z�q�V�H�h�����άM�\�U����^h�2�O�]�w�s�7����T1FX� �O0ņ�20����-�Zp*sG�P�D��~���D*\O*t6��g�<�_�FV�ތZ�)���D�"���"Y	2&�.�3����>�i0p�Fv�~��eW8&$)�en�Fa߼&��E}�1ƅ &��������y�z�YD͟S��?��_���8�Z�\���,ڤ��/��O�Ӯ�h��n�Z^�piC�Vds`<5���?1rF�\ue�	g�5u���	�&�=ᠥ<���#9۹��F��n^��_�GEdV�u�w��?���hb�S43�16ԓxr:2N�
8�{�(=dl=�l(��\�C��@h����@Gx&+�Sp}`"-xW�'l·e�s@��������z.�>������C�Ey��l|��i�N��{/��π�7�O��Ǡc�R_8D�:gy������S��)�z�Ү�|⇇ѱ�C��[���#�d��%9Y����:�����^��1����l�1���'`T�~����/���y�Y��V�k���\�k]�?�cSo���U<���d��':�cp�?��sܲV�w�=l4�ɡۺ��S��u$dӅn�L0='�G>\�eN�Ɋ��1m�ˆ~7_t�Ǆ�
�҆�;ˉ�5/��6,é-p�����qS�폾y�Q�ˏ~�SeYN���z����/���9��4�f��r��A�+Ս�r������"���Z�6��w�
>�2�*5M�o���Ɵ��v��{�����v^���t��t�e�U�;h`3h����J��<���v��	*� �>��� �R�='�p�9�o��9�K��X���͠��<�:L�o+e��x.�#�/|���ǝ��Lֶ�:����_�����E���#��^���JoJr�E��w�[������c�5[�&d��D?W���\E�J�2���3~��X��_l�ꡩ@�x�"�Gh�;���D��0��� �`SP>���=&��[<ڑ��F�@!�D�����o��X�,|�]3EN�S����qWq V#ɢ�K����"#�tG9 coBg���C[r��
����z䱠�l��2���`��U!:�9��f����_Nj��+F��yބ7p�V��8�ZeS=Ǫ��������)q8]V�uK*��q_�`�3��LΌ4{6�#*">������0��w�    IEND�B`�PK   �X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   ��X�@M��  2�  /   images/a63ead14-3837-408c-8d99-db2ce98ab1ac.png�y8�o�7|[�H�"di����Ki��-ɾe�)E�%d/bb�%����c�Qvb�c�����<���{�<|GG�q���������u^t����� A�ʵ+���h��w�'<L��{��q� =%���׊� (gP��%M��߽�����I�f�rͨ�����6G�0.��3��g_P8v��l�����+��8���O�':�ٳL#��/Kc_��\�U���wu~�4�@{\�{c�
��=j<]����˯�U;vj܃H�d�k��ghe���,�UJ������/84��!���Ϳ�˂���xiSSӊUL�G�����4q��w�ou4����7�:V���So������!u�ݻa�^�n��I�Oed��A���h�5�P`��[uG6������7بݠя�Ү����d�2��W~mcy��ˣ�a}�%DE����"+���G�'vmu�<Ƞ!���O:�G�'r����P[�<f��ׁ�'����Ms�V��iE0�?G��!��|�P7O&+]�:���h�K|DC�.��Z�,#z|{��#���u�E�O��Ĵ�H��WU�+����n�/Xo�pgC�J�8K$���b��m��
Y61X��e�_�ɫM���J�����S�>\؄=�~�޽ӏG���͉��D�t"!񕄮,+��E���h?�����"�w�ޚ�x�#�b�H��h�u ����u�K,�%��c�4�_Uuכ��Hӌ,o�f���:�T�[�����b�1~�G�/�ǟ>}b�7�e�w�Q�j�F�wO�x�ެ�_����u��d}�gL)�,XPY�R�K���<�h�)O�-��c����S$j��pHV�0'��"��}d�m��n6M���^�N�v�poi�c��m���\���Ϻ��u���Kh�{�\Y��B�����֥�~�q������K�y{���l9׶�?~|ȥ����(��얰�����}b�}����X<<��zm卑��;ʉj���S�I�@�3,X,���̳{I��O�un���Ȫ�EG�<'XK΅��Tr��j��f�}���6T3l�\��I}k��~Z@y��.����;S�PM}@;߯� �lH�IvBؖV,���1x�y�FR��ԁ�t�A<~x���.k`�̱��l�P�]k���+S��e��ꎿ�?�Bl3%a���/����=�H�i��O,H��V��z`����%�� `��`�%>V�ANZ���i�51��.=4Uvv�::E����?FXS���ZX����99] Z�OI�=w�-��}y�����ə��Hq���bȡ�<Y��>�U���*<��q�Ϯ9���o5aެ����8�@�x]�K+ 	��%#�`����iy��y�B�o��R���'�X�y��d���$���v�Tݛ?ћ��=�xps��g���ʐ�w�1�\Q�呣w*H��j��g��d\���9���t7�����J�/���{���L�G[��bL���3��27��x�v�}G룆�\�/p���Ő1������ N�#���f� ���Y#�$� �˒t�S�s��LX:���,�(�5��OHl�c�u��;��������GF�y��G;�]��x�bf�}�bځ����g%Lnn��s��ߨH<�@p<��%^���΀������^�~L��v�U���y566�M�	����G���qX�� P�j'�9�v��6�W���Ivy%��,7����aڟK�l��X�(H�Y*��L��1�S���CP�8D<}�`��|k����A+ڴ���T��Փ�6Ω�b��>�Lק�����V�K{�̐����RܫнHc��K]]�xtJ��;�,���4p���#K�+�����W�O��|1k=Ǚ(�Z+�f�x��)))�XHĆ�a�w���t�^s񈏒J[����0Jl���\��{+�\��Y�[A�+��8Ų�J6ES�j`sK�ðڗ/_L����v�`��OgɊ�c�i�s����[���ߘ�##�����RZ�X�����c����������Ą4�~���2�{qq�E
6YYJL��Hl��`L�pp���w�ڦ�J��ϱ8�SM�5^ͮ�G٣�.��u��0�X(����ٴ>��:�Y��)���EH�����>k3uh�UYx�a��I*^�=����(š��������ރ�>>>�
��Պg�E�Y� .ZI�N��\B�}�p'ҿVMIb���j�]�!��9+ǵcb!K~y0��b���:��o���fQ�nn7펲�\�e��c�l������������3a�+���s�%e�9,j�ֱD{{�'{��5Үē$���<K�#�;�eH�vwrr��_�Ԕ�⯽.�F5eU�(���H=v����e�Lo%���k�����/8�<�%�����[�s8�WR^m#���R4T��&u�	�����xx�
OW.Wlt���'o���󣛾k��}�n����>�m�Ԑ�4�&�k	�Hi��*2�_���1I�s��D:�L�N6�Yc���5VRW8���Ȫ�������N�sl^ ��Fc&������z�q���g��	��4nw�$���sMiU2:��z8)��$��D���;����y�Z�zlr��mps1��
j�Y���#���4�Y۾.e�{D詁�I�Z���H��GH�������ĢJ�e~�)��c-����)��7攔F..F�� ���$�Of_7=_5�,� �ߢ�r��iI�W/�������n �R_/^�7������o�8���<�.���RF��W>	�>�x�=�(_����E��O��M�pMs��/s����N��0�1�vDBJ*�._�5/�|���ي/�U�I^��HkOsKKCM͕��{��{O��/w*$nR��d�ͦ	���A�n"���t�$��>OTߺ�5'�[�lI����&b[L�F�A�<�ҧO����K����%�ɱ z6[��8�y�Q�V��`�f1raK4ɏJ�8�DwQ����Uz_�Dvk�Dh�.s�Hd��|^�Hx����(��!*��/_:����GP�ٷ��b[���!B6�E!&''�E]�v��}� ��I�DD�ڎ�S��?FGGp�t�te>nС�q� ?�8g�&�k4c��p��#��F,��EN��;=HW�>q��������K�����Q���Z�X��]�e;ƌ�y�z6��y��Zx1	L�)��j�>�����ז8�npkgV��	,�m���Z����I�"`�TD2!6=@�A(��v�n��ZZ�O^p"�\U\�P���@��[}��[\�|¨��e�u���=3�Т��XZ?�0�����[e�f�ܮ5�,�y{��ي �Vvs`����k:&ff;��F I�����LD������?~�uf�b���?��֦]�����w�`������Z�N�S�V�v��y�wA�Ǒ� W}o��H�L�PA�Qcc�<V�|�`,�}��y?]�b(
�W����N�مL���略E��ظV���n` ��Պ��5e��;�Ji�s��4Q������������O�����B<:�+Hao����@���hg���z�d����A�#�@�N]	��� �.�9�<t,���(��I��F������A�Lٙ���#��n��x�~G������/��s056���r>��2�;d��K�SE����s��CYIR�S�wOq�YAv�j��ާ^��D�4�)rs�Y���L���R�i�o�ؘ�lB���VK�*���(5�;,gb�v����$���떺�H�}n�{gL�v�Jp��PR��!g�O2s����` .}��!؄�4S��i��*X�!�=s_�=��W���� >����ֺt��_K�%��h���~�5\Ʒ=�ЀΩ��l��脄ȴ��9�!��3tVx�~q���;���C�Fک���{������ i�cɝՂDjȡ+(�5�]i � g"��K���nF�>Ȭ���Xk^tČ�8'Ѿ{c�c��ĜhF�`��7	w�ݿI�{.�"�R����A`ҶAG����8��g���&���5I%;V2���[�291��S���ɬ/��Zeڷ����kڕ�8�E��)�J!�H���zʫ�|�`�m/��U&���[������La��U�օ�>�i��8Aߞ�<�(�l�׋��I���BCB�So��B�Q�&I~�7��}Z���1�Pj?V�p��V�* {���`�n:�c"��s��n=����&1��~Z23�[6,L�X@���JFFF� *H��V���@#/^�x�3�(�<F��9sR�gy���p�O3�s�hR0l��Ҥ����뢓���]~�ctf0�xק�555��V�c/��N�홲�&2� +��g�{x�<��s)�v5�U��^�{o[���ii.���V��i� �q7��"�AU��t�A��� [�G!	���'�z߿�l$~}�2����?{�[{V�W!���I�(�"�� /���<��d�������V�}�����t�~2ٍ������ܜ_|��w%���{��D�(�K|ͦ���4m#��ͪG��|��C�B~���Ƞ�=u���)xy�N�u�Kf��p����f�V��oF$U�G
�(hj��BV�Y�W.Vԁ�l�#S���&cC��Q��oe8�x��*�������y��I###��El��	�勥7��׎�w��S�`bb����8�Է�\��l��"�Z�	����ݓ_�|@Hu���j�(~�~z��I��)|~��@�q�~�MzUr�>�-;TG	J�=��o�&��$%
�#W�����7sss�b�]���݁�� ���fJ*6`j``��t�i!�R�M%����]�yy�l"�������nڧ��m&~�њ���Z��-�����-4�Ikv�����;(�����z�(3U��6���A�@Dn�3/K5���߹���Ձ��\9S+,���	C�,�=ǽ�}�r�Vtpy$1lJ �EA�*!ː�W��,5$R���S���z�
�[F��������z�x֓�FTގ��$/e��^�w�����̒qA���&F~��`�iy�gs��5�l5��M����.�R��C�I�	la��(dD�[uݗ?�{�J�+�)��ӯ���Ӗq�
ٿ"�����ˣc�y��5$�����ﳂOl���;�7��K��]���Z��L���S�����ח�F�EC�m�f���C
���񊊊SO\k?���p,a�n��W����p}��{�+(��Ⱦ�r}��!�rm��I�]�!e\;�4�*��aC]����ÄӤu����ULMMzlY�Qq�фn�����`�ɳ�2+}�s������--��q�=8FG���D�m,�E�.,6��ܖ���2�)���'�9�k캡��o]�܇Ji�	j��s�*��D��{���ߟ_<�{θy;�gǲd�.d�R�\��nƍO�>7GuA�y��V��b���4������������i��)A�f�����bוui0�D3�)�:O���V�c������˯v���S^���R��	�޽;
�W����xuy�nC�D��|+{=�p�X���9GG�Y
��жbٔ�/?I�Goۘe�h������x�H]~�})e �J�Fl�W]�_�WG�Z�|/�[�4i��N\�(�Dǫ7�(����!`���a���ȕ��C&�35��r�H�Xb�:��!�V.�>�f��h�O��F�|b�Oj(�mZ�2�J,���'��K}�Q	D�	����-��Ve�������أ��٨檱H���e�<��˵���Q��������G�
 �\z���v&�v0M+W�L�۠�t�5��=~v/9����x�ƍ3+s��Nx�ʜ1�6c�2���׻�Y-`�P=6%`W�3 ���w_���a�u��zwj7���������I)�>zZ]F���硍c�~t�W�.6a1���ዓY ׃7Z~8�}9�ĵ�8O��j<�TE9�g��X��t]���MIV����}Kŋ?���S��l�]�+��/˫tؙ�׃,O(�ȸ��;�4�|@����6¥�WI�VV��9B���H�[<
����m�E�������[�����<��l٪έX�2��M�'n|��8Z�2�;0he�ڝ�)�g��PI�(e0X�b	|�XXy��ץ'��
��3ÂZ�d������)�P� ��>�-=�^�\L�]�/\yk�}kk����'��b_afSU���Uc��w���Y��Y���SK��Rd�����L�h�s׃�� ��3�,�U].�]-Ԧ�!���8�Y�%l�Ĺ����e(��6���1��l�B�dB�I�CE��`�W��b��N<����p��Tk2�,��{=6�$o�g��������}�C����y�����APra���w��YM�U����[��U�},Rr���9�@��ZldL�2Bz͵�����Nא�}6Yq����e�/� -\wJn/�������h��ĕ$)��|Refb��ా<�lW�9�T����`��b'x��}elLu^DvH�4��HՓ�����B]Y�����ò�~��?�z����O�o�d�'�d��(�R"q��AxG�d�#e����U.��i�r�j�_D����,!Sh�6cB�����Ǯ��+4ؓ"���kVsIY 0��}�g��=T�6�7�&��ey�@c��t�*2�����d�0����P�>�ȶ�)�Wa����S{S�,��_��a�?X�Ļ�����O�M�k㊑�\�yf3A�I���仱:$d���W2km�4�U?����c
7I�,����
���F�X~M�,�=��{M�ϯ.��_�W�b.<٘	�&n���j�X@O�88^�K�J����o��'���av��\A.��s1�6��'�s��Qe�jO��K23ղ�+Io5���Hhoui��W�%���j��m)Q��+�~��]3��F�-�����vo���E��mo��T^�0����R_s�U�.�̘���.j{4���9�J�$�O��U=j��|���=����&&��Ls�qzo]������ole�Z�ck��/g�����8�g�H՘�W��E�X���G9\*$���Mb�o;���g5!?����x@�(�Ñ	����L<���4���p���ㄡ���j������g�p���t������#=��g������e?w#��Ka�y�5'���WN��4w��32PL;�֫n���|ã���KҴz�0e�E�IH��ڠqa�^�P�$K�}-���^;q Qm�ʧ4�G&����p�ƽ{�~�	�����Ync��Zs2��c���LoK=M�M�<��k��ﱚ�L���tL�s�S=���Ǖ0��G�����C���0���u��j�዆~��.J
�Z��ү~��QƧ��,�w>�P�+�]��H~cm�u�W���݂�S��zK����*a�ONu�����ui������'�e6^N+���z��d#~���1��^�}nf`v�~݉�{��i�ML�Q�L��ӗ]��Jr��}pP�Dֶ�׭.E1BP̾�:�Cvə���`��w�j�t���n~�����%��i��dTOx��:�V�k���XE�3f�W�U�Xm�I�uNZ�޽�C���V�	��6R�F�ʂ�V�0?� �+ԠQ5e!#�sڠ܀�3�4un����S��@�a��-�w��Q4Bu6��˧!\wD�{�T'̾)F��~�P�ǖ�j��)��)��dg�5�
�+��<SP�g���尟J���%^Z�c������5_'bo,��@#CW��|��'1ʌ������@H5��p��4rxF�^$H��T^S���D��ҥ��W&�M�a���[\��]55%.w�ܗ��,?�أ�؞�u�v��v�wi`�'��1��&)*0i�ʳ�t���	������x������ܧ��-lm�D���^�<t'�S�0��q�J��l"�С��!٧�@�B��i��^um���|^԰t&���n:�߿���Ʋ���q���܌ׇWן��a��b��Ģ����>NY�_i����J8BG�����O�r�ј�/�i,�jxX�쵅�޾L`��PXn���K,^_�|~��xD�-[c���Ox�)����+�>�Ś�^���]�"^���}��5�� �Y߾�U����� V�jh==~�[�DCNK;-�H�&�C�?W�g�:�Ww�+�~]�%k�XEKll�����LK��]ŉ�a��Yd��_��O�JH���:%��'p��մ�@r%�v}¥��P)"U�&�|�/��Q���ø�:�������ZQe�����ӑf����訇�랏��n!�[����Լ���GZ��?̦����' ��
�Y��νZ�s+7k	 ��K(���b��&d���V3�N_<�Y2c�4cKe�kv�b9ܟn�y����sÍ�Do��ʖ¬
]���Ҭ#��XR�n�������iu��'k��k��������]��P*~�s��<��T�9a�i����w���T2lZY�}��Gqs�,4sL��P���#�<7�KO�� \\��Kcm�������D���j�:��^?�5T���~*�1N��Mş|]�\����m�B�">[׏~+tP�~10�����ݫ�p|x��G�y��N9�i��ӵ.88=L�X}Z���\e�M욵�Ϋ�) ��$$�����{ս�H�%ֿ<����ңA�V:*��|)y��$��c������y�.��ERT�{|�(�����j�~����L�܏?�7�c����*k�|�~|����E֬,|�uFr]Ϸ\�マ���WO ��9s#f�lb�?H�����n��9���A�p��E�����ʩ����@<�'�o�W�M�RT�F&^z��N�T��~��O�K!x�~L�M]��x঳φ���~��w_�j������
9K�k���0'�3*�Q��`��p9It�@Q$7\`G�h�1mM$�r5q�'s˜�A�zp�9�M�b�]i�r]��R�Q��;���}�aF�UK=Kӷ��LgaQW�C)�򓳔A��`J�|=Z7�!��d=`��Um!(��v�<[%+��t�f�w�Na����WeE�E}'�Y�W}ks�&�J6=T?���+�U%�[b��EC_|�'\���r��< ��T\�j�!�\�"QOEjrl�bߣ�RT������I ��QG�ˎ� �H�.�u>��/����1�Y:�x<����3��\v��r��4��"/̷�@�Kʟ��璴}�[ꪌ'��.^�ny�>6λ��}���SQ���:��TG�.��I���=������d��K��7�J&���ȕ�c�����N�+���BϾ��a�T�GZo��n��
��e�܇�����>XP1�Th�WB�+S3�
-=F��F���<�}Ƌ<�8d��$�;�� \�}��Tԃ��3�L�WX�F�߹۸��j&tvv�|��^�Ƶ2��t�@r����g�V6����,X[oMvhՈ��W���{V��H�N�>��M��n�vT�2�H��z�A�x�AhO���?�&�-�ŧv0˃k��s oB�ƭ�Y[�gk�%w������f�12��	-:	�1	o���ݡ��Tb���� ����b<������a2�� rk`q���Z ����a�T�éOQ�)��x񚝍M�I�h�F���<�q�fϧ6n	I{��%�ߊ������ɂ#��^3W?��=Aw4û��FC'��5�ܤ(S�����m�2Dz��u�?�)�e�zx|`���g�#���$i}%/�
�WI]r��t̾M��	��N!�s/����񉉹��&b����>cs��4O�63L���gq�3��~�<;$
wF��6o@���{]���'r�����}CR���/��Y

sR9��KV�d�z����"�p�P�HDK��'Y��H�ƭ�b4������s����[J�)�9M�D�?y�c���,��7�t|�:v��O$�����b|���n�gu`��Q	��b��4Z9�f!�@s�Ҋh�X��Z�q/c���xo,��K]L����*��~�w�����T@�.Ү�-�du%#֣�q�F�o�6����H����-����sL8B5!�$��93�9u!K%ޅ��!����ϯ����?�ʱ����[��'��#Ezm�;7���vp}�Ϡc�y�'f�9V���p�ḫ�7�*=�lNm(mi�Q����6Oi�z��O.�m�iT�*[ed��1�Y��w�p��}2�ߒz�Ӊ��P�a��}�Hz���@�8`kkR�}���/B����M�'#+JΒ	%LAe!^����샴ӑ@�Ŧ���W�9�?��b�J�p��_�R�����p݆�ۨ��̓�(~�Z���B7�>ĥ�0���]:��n�{����ٱ���I��E�?��>z���lg��L9r$��͊�d��Vq�&�f�K��*Aa.�2�2��
���[r�������>����٨�E��)����0�ơ�ڧ�auڵ�9+z��C{QT^a\<<rY��D;�y;60$�X�*���!b�F���M�P-W��U�����>��o��%$�~��[̘vK�ya�=A��?<I�=�5��E�j���Ɯ�G�Y����w0�����䢋������x�����f�БdIS�3A+@��Rڴ^�<�`N�k�8t��v"o�WK��aA�c�,��Τ��~E�����z��j��! ����������1�|4�SD5]�v���m!�n���{��*�P������?J�0�]FFF���{�������S0��G��o�_��贲�r@Wz@�;�c�<a�G��
/XP�66Ff�Ú~�-��5��vsJ�L�X��;���T|G�UĮ/mm|�
�:؜x��G9��g2��y�~8���ҫ�E<5��
|ܕ�)M�'�6I[0"��N�E�T7h����oq��u�~H��;�}�X��gx�$���j�h5%.,�8#P-/BB������J����[�,⑀��;Ԑ�3d�<��c�Ζ�}E*EvQK|��*¬=�Zj�k�=�Yj5�����[��U�/I�%���M3���wI��q�ԅ5��=}�~~@bF&+�'�l#$e*�^�]dɞ�G���H� �;�$�@�x�
����ٚ�S�2ngc�wY��Y	���q�9M�uV\k�]���l�t�h�1�-b��I� ��O�e�ӟa�nO�z�Ɠ_�M���Sҕ�!�r�#��4����q�%����%��j��T�ii�M��	��'�%$�U�N�L�O�|5椫����E��ˋ$;�.�D|������M���ˏ����1Qݳid�Ш[�{�d�u:�Q%
��\�*dfM���1�z��ߕM?�"8~�!�����>�9���80�����lUy�ؘc���oi�Qڧ����B Aj޺�� �<_�a���?�^L�Tl�\���Y����(�K��)I$Kï��_[)	X���`�ّ߿�*���m��}��C���w�b=��૮�1Jp����*��Cg+� �T�P�l��>.ƃ��%�.����]���7I��a�����ؿ��37}7�;���
H�|�����z�}S���2��8���W��c��洹44B,U��_�^����� P����b����[�	'�z� c��x
��H,�V��R���5���+��wQ� 9�U����}`�P9���Z�i�p�	g&�8^��)h�'B#�ԋ�Z�+�x�� D���*T֗!�H�%A�ǥMO'D�Ơ8���z�q}�M�3>tR��d���vV�V��j�(d}�e�d�Z��=�|�f|ֆ�A���{~�}�����@l�C��R�G�s�i�0j�_U��H��d�x����
v5N�..�9  ]A�mC>����l ����ۤ�Z�ѕ��ڡ�|5�x�x�s/}*��7CaiL�x̛_H;`�u���Z��3����P�h�������/�<�5v�v�����dL ]��
h���+Ԯ�1��fE���� fm����]evw�}4�zoү��*a"TO�x�xW��l�7MS0.��f�ڀ�z��c¢�̱�g�Z%��*��ޠ+I�DbbːrDzs�r�&�P���!�����5\�v2���q�p-���	!'CQl\��q����IUWi������v��3[G���fe��9u�MD�e�g����g���80�_���tP�MOO�O���]�;N�&��XS}f����\��f��4�v�J��rr�P\J)w��nDw��+��G��&<���zW�<d)�|��)��+髧ix��f�S?W����� ��j�����jp���h5�"o/{�Je/��4��;���>X!p`��h7�®c���D+�>��U��5 [��=���7C��h<����E[SS����=n����h��Y�v�;B����ǿW3�[��6&mװ"��#�۾R�Cx��zo�8���!�lY?}��^�^hr^^�����R����
?U�Μd�h5�/q�/��n�r �F�2q"�1�?��cW@ +7˽C�ob�mgdH��w�P��6/��#�D�|�ؕۤ?�\�M��h��ߍ���R(��s2L}��^}��-�q��Q.�g�bR�Sy���� ���~:��^r4�ۍ��+5~Ǐi�թ�VN����/~��j��	���/���4g����"|�,����ڴ8���n�guq�?6�����Pl���"��+Q�I�~�^��A�E�6ϕ�5��o7�z��e��l�ף:��S}�:R5%�!���u-�z����N1!0�h`r8����?5^Q�����ԣ\������J�z��xC�0� E��߿3��%C�@vӺu8�����T�˾��k�BnվT!�0n)?��9��K���zHX_��a;����*��۽{�U��"�{����Y���^~�bS�
r/Y��Պ�:���*�?B����N��b����t�Wy�
R<��}��� ���5tt���Y;�I��tl�T�/˭R�|�˱�:X�IQ}�t��d�ӧ�z�4����&)c��J����[K��b�Ch�����~��H_�)�\vc�D.�BIs��XP�K�Y���3ͥ6z�u�H���|uuY	����9|��h���
r33�Z��%��v�*]<0o@L�͚nmC����j�4���F���*�I���f	��ق?����8��{�ȏ����Cn��{C��Y�Ə9�v�y;E<F�O` �6�ƍH&�÷��w��AnW�e�nP�|ޟbZ����b
QNg���Jئvn���_JѨv(��*�(�. ��5��ojL��pa>��~1�q��ߋ�����G$tAB�J�h�Gp�F��&�~�<�7}w|/��Z�f&�e� ��2�)20V��iOs�o��wpJ�*�;�����R=�(���&�ݓ,���t~w"��*[��%�vZQQ��h[(oe0J��dTV��������G����u[�fꗪ���w�O:����0a���v,���KC4
s�@� C�)��Q�N'Vo�V&5�G���w���|�������\;Z�@u��k��Mcu͟P[����S������pᇿm_�}�!���iȣ�kZ��w�E���Mc���J���q�}�f�
��������Jf��ع�8��^��A�����9iq{+�4��F����l�K��� Uޯ]79��Ḣ�3�Y|(+ �w��6�f��u''~���t�/�ݲ����_ׂ��Pr~��~d�V4�B��l ]���ֆ��D5n|*˖��9�}���j��p#��饉�������'�L(g���.�0��~::�,@�Wep�?W%��D@�7VB�?@��S*��7n	�ӎ*ۓ�5Ҝ�t�X��������2�H��2B_�Y��)�SC�ɱ��?����eڻW��iP`ŗX�,�I\OѸ5��}�֯��P��e˻n���$�H�ʳ"�#~J�t�1�> ,9��F�t�����(�s!�Wh�U�[�F+�~9((:�#:..��Ai+���8�^ �js��_.)
�P�Ɖ9��ޛ�Zb���v1��K��>�]#{��0� �/w�RMAnɺ���%j[|�y��N�����Z}�m(�����m@AȌ��?�h.���u k�����A��S���n�{��#蝻5�=�1���[��E�T���qT��!��v�g6�� ?�y�'���ύ�o��ǝ�n5�P׉T$��X��y�L��v>nyy����;�TMA��������`���Ӧ1���No=�3�"�˺�W�@.��G߿}�w��//o�q���ڙHUL[	6>�܁�>b ���Wm�D�a3$X͍#s E���K7�Y�����Ի���U���^_�8�y��]^O�Wk��NA[XX����}�`R3
��=�N�:�[��&�����ML�����ѝ	����b/�g���>4[ �};2�(�,���?b�+�P���
��Ǿ�xG@$�C�v|�&11LЬ{��3sGU�?�A8�9(I궃|�_�亜����/o��HzpwjH��Έ�I�g�-��>8�P�d��D��[b{���~_"��C��@�:'k�����`rٖ;��G����B��K�Ɉ2��w�옝��1�;<	�N�H���y+TԶ�u۟8x����95T�g��1 O�'��T��ظV�䏺+O�>�&�>���Y�s��~��w����G�>~�� �3;ʹ�y��X�_a4���&�
�\�1�shn�|��I���
F�AT��Rxa1�������y��P]�%�����/�\��rJrH�H���=�����ii�<\i�A�-xGP�&��"��훦���)d�ó=���n�!�����!��[�֍�.-5�p��[��U��d�F�wF݇��UTUl;�B�BPh4�6��C��׆뀫|��ԙ7��w�&���a�6��&�$')c1 �"�m}TQ�#��PO8ؓ������ u������u<�~]A,�w7�q(V�	�G&�_���C��%��A�'�*bJu��6�B~BX欼����]ʬ���]�D������[���&��jz�N���;�6R��Z��*e�n���/��ǵ�|W��*��Y뵴ҥn����.[�Wb;|7��T���t^�ء:���5��r�~nt�-uP�I�ۯ�菞x�M.Q_�s���t5N��E�V�h�{@�%�V�n��$u[^K[����Mo�%C�B�F��t%�3/.h����J��R�8����|�8�����J����3CR�a�ҝ�Y0��_�D���t[(k�J�����L�Ȼ(�l���w�U��<k [�S��]�4ӛ��b��,��t���/8i����S?��ڳi��&+�c��|`3�|�ji���.��v��<����j��	����ͣXMC��7��6�X(�B�wf9j�R10a��!�缵]��&��!yZ��j�zl>t2�s�X��H:��O!8�6:�%���P% S�^�L�?qq�\���v_v�df��F�pI�`ie/��ΘA�n��Sa�%f��5�zz��}.���W��|?J#f����9�|����(1Ӄ��V�Q��y���+��V�C:�ĭqî\�pj��p���2�t@2�8���$q.��8^]^�hX�ѧ��W�F�����]�-�θ�k����z����Y��4�~C����)��ު�-\�G�F��r�AȦW@���[�G̈́����X�8Χѷ%�4��d��m�p	���=!���^�^�,�oE(X��_V7	���2-9v*�����{�o'�㨾�¹�[Ӽ�a�e;��?�}������
<���:��>��ޯ�:,�8�D� ��b��u»;�b��W,�;u?״Y^�wB.Nnu�Q���l^�ZA�33mҹ���C�k��ZA���֝��xȷ�{�߃�����_���!q�Ǯһ�'ۘt5���S���]�� �4|	�j�*� �>õ����8?h����Be�b��Vp��eg��Y��_��3�R929T*�:��	�c)db�$C�T��:\����R�g�r�m�/ɋ�0�,	S���g�K����aÊ2�������*?)֪B���;C�$w��@x	��x��%�R̋W�J��P��H�v�{]����>�?v���͵%R~�56K�������o��W�K矐�Wg� e�t��m��Ʌz��������]:����x*�;L~�LiU�Q���C���6�c�L�o����6���� ���#>_8��}�Y��ȡ��ag���T~%,U��Qz�E��`�xT?��,�-�v��Y�x�MZ��5��T�	�M��+@��y�]6���Ҿ��[1�6���ݽX���x�:,G�.��x ��P�Sn�9����Yt�>�`�yăW���|XO���.�����o��g�b�1��,wm��y�|�C_�Xj,�ʋ'K�۴-����l��񭝫xJ����t��v"�g;��G���DE����Z�0K����"���� A�=��_�zWT���o�u`�jC~?��_��=����{�߃���� �MK��i"w�ʝ����ɷԺS���N���8�0mzs˥י�q(�n䙂Τ�8D�Z�6ð�"�Nn�����'�rv�y��-5n��XQ6Oʸ�x�WM��<Z����
�[ا�໾\�x���(d�3{=��k�k(�s��&�2�Ѥ��Q�!Lk����o����`(���C��KW��ޏ>.�Z��X���W(��~3��;�]f��ϲ�?�`���	ʚ���>������`�Z=xD�4YN�+UK���{S��=ie(���n֕}O��3�幑��5��|�:�2�����F�J=��g���a�(��~fU�I$ ��]��r|�e�t�()�o�d��e�|m���ú��s�m�rNi�����fR���WH��b�����Bf��(�Y��C�[�z�N�}~�%�.Rj��G��6A�RY�Ae�N��¥� .�S�M�什~�?pa��&�7�I�̥;ϻ�l��d���]��/vc�K'�3W��~7	CJO^8�[�ላ(%U�z-7�Z�Q���9^Ct�����Y�:�Js%���܌O�\��v�s����Åǩ�/V���Syq���d<�yN��[�_OfЪ�*s���vU������(�µ[��S��~E�!~�ɒt�����:^�2A�gbL\W�VZw}�������3������]
��7&`sO�Q"E��o	��Fh�yO�m��k ��D�J�����<�+��rK�����+���$3�M�Q��w۶l�K6 c�H,��+9gk�Q1��v�(�M4d�᯷�p�>'���P��Z�i;��&;7�.W�wc��b�C�$3C���|��	�v�(Cw��h������i�Z=�ɝ(��L�l4��T��h�]�+p�$W<z<�*$�:2�/P^~&/��
n�/Z�0<\��/��?˼1ͬ������ J�T)ɀMX���bʩaB�@�����H���hY�E�J	�
�EW�x�FJV��m�~8��h�=�1�J=*=u��R��p��\.N���._��[���IPS9G�{��O��h��q}�0P����V;U������{�5���� 8��6�� EA��X(J��� ҋt$��Rt����P�I*����W�% - ��I��s������ˋd��S�羟��vg����+Y�����F=��!^t�ߖ3��A��S3~�FFد65~,r�)�O��O	1Đ��q%+�U~���G��ǻ&i)��²,�+rX\�{���oTX�\~U~g�M�3�lM���r�At�{�7{��wDȄA���G��GђS~�S���]���mq;�]H9�A�8v	f9^I�1�WO^RZ�<�bs��\���\��?e���� ��:b�S�YB���wO�k�◉=�)0���n�K�Q��S��̉�J"��YI��C-S��6�Q��D��z'���Y�������,6*EN@m�g"����N�os�N1�]w��yY��օ��ܯ{1�a`YR��d!�]�R����	�~�V�ｇd-���_uLl��+1��A�x?P���E7�kװe������g����w�k]�A^���)˻a]�����h�fo�Ж}���&����h���W��-eT�rN��0+ߟ9^#��1r���vCo�B�]���T���&����:�f���K��ߨ�����K�~2G��>�"w\�~��㕡���ܨ���G�$�t�7?��g#%r/��+-G1j�=��f1��B7��E���#�Eϴv�&_ύ���XHm;�/T�čs_s>�1 MkTt�l�-��y�lta�\��\ ��q28�1Ja^��V���l��c-��1AoB��9�9��{���I ��.��q/�ιj3��Fol�|�)�y.B���P�է��.!p��xSc�ZĘ�¯�g0k�J�����n����[�Sw��<�Tk��f�W��y;"l#'���h �W���$�J��nƐb�S;��H��DSBɯ�_��C!J+˞�W��:�E����	���*r:���<k�༦&�w�y���Ǯ+�!�O�%�m��U��k4)�D�.�1
�b��3��ϵ�'}Zλ��I��c�&?�t%M���bD�3�2�}%{2��ʰjsi��y��S��eՊ�Q-�<����Q���a�X����>�O�]���..V��� �������m�A�9߅��,f�}Km\%ѵL��'�"���z1bw��ظ�둟n�uO��d�!	�7�[���۴3��������핪�ɫ�T�=�ZQ�G�kU�a�غ�ۃ�לB�J�l������:�M�JsH������<!��5$ka�<vc}�k}iBU��U���:��Q: �O��);%�k���a^ZŲ�'ri���}g��=M:�d|���~��	�G��q%���!�N�m���e�4ks}�LVRS��jֵ�F�x%zfﰖw�p��}�Ő8�!x�8z9�C���)��H���<,�N5_���}�U���Z�{f�1_��Y=��Kм�(�Ŝ�؏���"!��~_��9�`ۃ�;���z>�K�J�v���~�UFEԅ�Y+v��Z�e�X�;����4��$�/�ߝ��1���`{���E���Ыv��~���&Ԍ�4*m�?�pBz)����
M�*$�!���0����/-H�tۛߋ3j����ƞ�Zۦ�5���ݧa������?x߆��ٿ7"Y#�t�WZ �TFX��������;\f��mB�i��ά�}eg�}1�?�L�>��P{x��n7��M�#K:5f�qB��m����xr"� &8{g�L��i�e���{�u@0宁���jGƐD���֧'T��'ϴ�J�?�=�{9LJ�jԀ�a�T�> ��g�C�L�WN�;^ñ0��J���L��ĸU&�W�K�Q�ta�
)�Z�s�C��3[�G{�9�9#R�6lZ���~��s��ٵ��c��{�T���W9C8����ɛ��z���bo�(I$c h�,��YmS .�90�d����9>g��j�k�3�N�^�N������ʩ;���٣&m�F��t�G���j�6���'���n�U�G���q���'rșLǶ��"��O���;la�j�b��F4��An��Թ��p8�poq���e`����}�Op��*q#�?�6���wP6ZOJN�Yj`��L�V��H��6�����˞8v|y٬�>'��p��ed�i����f�P��Y0�:��¸⎠�3�����ϗ=����J:�
��a��w���eh�������aʲv)e�3Y�Nt�]y'�ʩK�\�rىB�tC=�4r:O_hUY�)�xJ(pE&Pj��8�U�z'b0��V �C����p��%��~@��l�Q�]1�o|u�1�?��j{>(�@�D����e������|��ayT����/z���U����zc�L�L����F]<�;X���xt��a������"3]y"|*-��%Cr����'p0�H��MkiP��%А���"���y���\ۊ���U�/�.��|=���5��J�CS��j���q�]�q�k>m��%i�<L~^�ȼ����/��L��w�'z4��r21@�lMV�w����#s�}����:R3�D���*�ڵ��ڱm��N�1�on��~��.Rv7��)�;�[<���r��D�	�+s%ش�_�&r2"��H j��d��\���^"y���Q�8�b���F�ԟ��[�y���˾=\8R(��AvM!MU
���K#�5��K���9YiE함�tf�}�K��,�F�@���O�Y
�R���T	�4�Ijs�	�u~�)<i[k�^\���P�������n�2���a���.
Q��V�Z�Yk^gč�M����C���N���p[]y7���}N�_���������b[-��\qK}��2Q����s�]���<����yW�[�es ��i7�GM��i��@�'��(O_�CN�n���K��T�Y<�����}��]Ŷ�<�=�&�R�"w�4�,�c��wN>9���40+��S��WY�m���٧V�5?�ޢ�0��.��₞+Gc��Y���V���*s[ɥӬ����X�&�^�1�J ,<}@�Y����П��&>�u^�5�G�zo�<�]8ϩV^�4���`^�aEP7������mR�����M��������[OM74�V�eq�q�w��3PI�[���l�~k�m��p��+v��͸�ɹS����������ͬ�A���@��n/?��=O��ݣ��A����K�����Xk�F��/�I�=V9���.���p/��y���7.�)Ё��u8�3��Jf`��������_����C$��1T�3/����0�\C� j��u�}���p�	>�w(�"}��&'f-��H�`�*�\�_�|�?񽁒�W�y�d��*&6��?�!��#�d��f��έ�h�Տ��\�����=�ִ��1��Y�X��C&F�U��&�>�/���x�	\z�o���U֑��u�'���O2��^�yo*�W�FP{<mz�n��͘2&Þ������������}�{y�?�{�n?�u����2���x�zU̿oV/��(�#W@������Z.���k�xPp���&ɸ�ԡ��`b`�~��Z\�f��G�9_�����ư³�R&�*��iκE�6��JY�D�\J/�-���o�)W�Ǉ�~㱳F(_�?S�8.qi�a���É/�K�=�6�x0����m=��}�|�T���(&<��N$8�/�"��{�!�7�BI�
��_m�h�N�s�0����J��ª��*$x#I��2��~�T��s������n������2�g�,�œ�I�C�b�TVK	�b���fL��A��/�s�Od"}A��A.W�9�)=l���_9@��P�8���^s��C~�sF)��ԽC���ϧKg��5��<=yɰ�����9E����[�%Uo�︜���Nt�?�v�<'�m����+J��웤!�|{ƌ+z=�\R�`�=�mʫy���}]�rȑ�����F� ����ض&��q��GXg�y���
���N�0p����t��9�X��E������'�9tx<P�}1*�7���S���]uٹ��4H�p�����]�N�Jr��Gm�D��&�J�bn|�@�c�ɾ=������Ơ3f���%�!f�E�%�i����xM ��z7�f�k������R-�
{��XP�*��dnO8Y�$B���}��?E0����f�"N���&�?���XX}�[3L���v.�k`�lND^�nL�B�V��-�:������u-Ruو�f �J,1ї�ced`�������{6�,ّ�%��P>�P�G���;�b׾���&�@#Ha���(�.L�xzۛg|"�fn3G��=���h��| ��V����%3E˹�I�$'a23��;�w���󂣖ɥri,��}�T�ln���J�[�BY׵�=�+�ϷD���y�в�5��G]Gy��X�ȱ�����w���E�vW����Զ�
??�����}@P��=��C�e���]&Et ���]��an�ݓ�Aq��:c.r"C���b��P��w�d��٢���.g�]�RV�+�
�{�黍g��6�8��7�j�D��-N�c�+��9��>q�2�:�ߝ�7A��Y�|7��s�^����˵�l�����IY�@�.� {��Kr�������`�{�+F��M�{�>��'}�+�Pàn`�f`�h�
(����77=��$���'\���*�D�����M�ۡ�u��G�H��(͌���r���LL�rHa��o�w�l�;ڦ����mj��v��^�k�	=��=&�b�IS��S��h��~�ș��J�?���mH�Wu�U��~���gp3h/�����a?6�Fk牳����{Z鈳i0 �����H�9����-�n�u���7��`���R4�ٍvQ4ٻԲ�Nw<!T�_o�P9Հk;���l0���۵<>�71�R��P�� [��BD���ͳ[-�u��7�)���Ώ6	�	�S�2�W��2��o~Uk�ho=V��?Fd�0ݥ�;_���� l�Wa�vzX!��\�����"�A��n�̤�:�-�s`��/'��'��\N��'pJX(����w�t�;�'X���M�,���*.�1=iUn~n�Z��?)X}a�|s+��i|}�1[,Ho	�
����-������"QR��Ak�W��a�s�{1�e+�)�p�g�mC�[C}Axt��$8K��V2p�Y�������a6���0��}�9�V��t)?#rl��ն�V����Qe�T� ��G� �_9͘�M��g�Wٶ$ήR��Е�LJ�Z&�l��	\���SW%���= p���~8߆�aaPس��4N̴��g�@���h$ȡ'w��8Ə.<;jwT�BK��|a[��H	׌dK��J|�c�ů�Ծ��+i��u����I��Z�e`H \_x�4|�k^���.>b�S��-����|��W�Ƒ��0���LÝ,�J��5C���u�\n��s�T����=��h4��Z�Y���Ч��}<쳪�ֶ7W0#����?�ڟz�b&�,���&�ڗ/_�
��<P:5�%��i�O��?�(��lK��ox
�/��t)S��@�U4mj���ާ�P`�8�Z����g���ÿ������+�^�Y�\ؘ7��Qf��"c��=���O����v���]a����N�~]���n�l^�Bk��Pdd
�#���qU�99��M�#.��̯�|�z��+�}���R���D��&^�Ŗ�9LU���L��X��5u��|� �����H�AW��"�ԩS�)Ĺ9�USl����_�i�P�iFGG'U� (k����gt�RR�J�EQ�mmmZ�V�\`�Z�lyg`�l����7��yF~��d������ΘĮ�������b]jj`����v�l�_o��]YU�gddt��_/>t\�����']`��Q���M�=�L��oD4_���p'W�} �W����m1^E�B?�����_�F6��c/�2�/KKg�U�<�[\��6��Hn�@��s�\r~})�w)ʯ�L�]���������ݵ��x�l��
�ui��)��K�o��T��^xD�M%���r��602/u���*@�� �[ifv>>>Q���L6}�c���}�h�N��R4>榩8sKG~5�9\ Bq�,�2���шZޚ+�!��f�5p��G�W��^��Z��e����]�=Z���oB�=����Q�S,�F�7-����G�.p����Iex�I�;,���@{"�NM�	�Ƈ�L�f������d�$vga�XwZ���i5����gCCC�ee�sz-��1f$&%��/�9�h:���(9ݏ���!ʤۮ �0��kdA���������T��,&RN���lf�+%��Б�2�����mu�[+P���b�_�>�e�f�{m�c�pb�J���Jt���[��/A��T�­+�=v�T2��o�`�\Y7�� �v��@�Sݏ�����,�[s��9}�a܎��>%��q��C-�kR���yӶ��X��J�Dm �<�	�e�����[Ri�ߣ�KyF5y~����E"�g�R%y�'�o�A��Y`���� �0���۲���������<+�Sݪ�uK��I(�KKA���l���*��ќ�2�� H��C��!'. �z}�S)����h�v6�5kWf�۳�g��� 5�
zB��7�O.҈�k��<��T�^�s����O]5#h��|���>4]'
�4	�iA���9 p���h�����q�'\��Û,����}��X�,ɡ:�,/��F��Gi��Zp��]Se"���Y�)]�ņ5���>w{��p��w$�D��ޜhn���G���`�f�f?%_���۰]1�����?�r˩?Vɛ���lW�;/��5X�A:�r�L��˨��Jk��|��ڍo�5�%�s̖2�R�n���'cM]��*�B��[�H�wzJ���͔@9,�>Q��ͨf�3�z�a��u��w%�I~W���Sc�6��~8h����� ��`�*/��t����=f ���c��M�~�}������x�����һQ�n<����[O�L�n�	�ǒ�?���vU�4g�b��K�)�\2��ތR�$3w����=>�D=��J�D���iM�-�iv7C�%�fU�e���v��?�.���-��������҅.�hw�s�:c@uE�E��RGGF<k^W�Ǹ�`�� //�B�5�!���۪��H���P��pS��gо���Q(�83�[E$/)+F'_ߍ��7n�஌�*����w~��� ��p���)B���j��R�+��k�.% L�<�Q),eN]�uD��-�kR�Vc8`h2�?r�.��&�0�9��D!EQ����t���5��"ŏ�Y����%�������M���;��	H؜�'l�P������l%n�	g�:$�=�Sd �kg���B�Tm<r*M D�y,�Y#����>ϥ���%�0��
�ݥg�Y�������sa2j�J��U.�@�ֹ�cz�s�S������m<z�T�ұ�3��u������-�E��h�Oc
�j��X?�1�|�.�� ��$v��ڙw��(	vHT/}��,6��Ʉ"}��-ݚ�ҪP�W���lF(�x\ڋ o�{��k�$��-��5uxX�{T��o}��L)�]A��Y���;G�G��(�Ӈ�w�?4�����͆w�^:m1j��������K-�Εԍjo��F�f���t@���F��?gW7^�E�s��D8(�=:U��[I�}���G"��#@�ν+n�CP���μ�z~�jW����ڭ��=S�s������gE]�6��q�����T�������쮈�Zl�qqI_��;�)�J�Վ�������2C� ����݉�����	�{���M*)�*y�M�[?�)��[��E@-�7wŨ��5�:�]���%�QC�V����ms��� e
e���Q�;~|c��O�y�9o:b�A7�'9�A@�6a��S *�ox4�<�'��mʾT;v����5܉��7��פ����ռ3695�5>>.���J"�o�n��qRq#{��V�q��*u�N��Z�XDH׬�u���+	x3�ت|�L~�`������/'U�EsH%�VW�����@/��I�J;8��~�Ў0x�-b| ��:Ǯ���	@�*ǔ��H�$n�j��{Fyi�3KjQY)��ȏ?n.s�D�Me��������ڝ-�i��%Ƚ�������Q�8
�IB�72x�+ng}5��:3���cW�-V�W����ȋ�yȴ/6%� �ِ?9�<��ߨhۻ�hX����6�|Z�R�2nW������0��i%D����O��L&��s���������.�Cp���WZ�О�2��h�ll�n|+��i��E�'�Y�Y5��\T^�m�zK���*��n�B����;�&���p�G�f�
��ᨆ�S�#�f]�M=�{��O��k��4�,^TTL��ai��*cr�ߕO�X�eɊ[�C*�n6"���l<v�a�v��c����~o�]��Լ
�zp�ޡ��~g,3C�����R=�7��
��k>Ԭ����Oi�h�F׬R��3y��_�n�Ta?�5f #��L	��Y��GCFF�
����	���F��bT�z�^�� 
�BJˡB�*紂�.�F\��UJ]�?�`��[���`��GO�
�\Qjj<��9�}e���f ��G�`�B���\}��l�\TTt<.'_0�jv�{Cv삙��a�Fnt����Z�;�i����U�B��\���VӅ�KQ	Pפb�.�a��gv���l��:���zi&�'��]��4�t��m�܁�\�
��{��;����\��sEQ(g����K��{�(!?��И}V ��0�Z;0s&�j5�������v{��+�@�{�W�䝕@�h���opD/��I�wft: ]7�kdǍ�W��-!�)�.�&�wĔ�G�ݜ� @���jݡ}Sl����ޛJ�S�6xr� 8B]u�P���������i`�ܩ_]9/��:�t(!j��9/Be�/�6g::�������5/�+b.]W�,��T�?pojLRf�Ϻ/${걺�$����=�ӡy�� ?A��e��z��W�ה��8!,d�]�A��,u�2R>yM���#��P���0HL��K�Ml��S���wܱѭ;��ԩ4x���f�-yH�r�3�n����+=m9w�x?@�JGgPP~���n蟥>w�-�+&yQ<��$����s�z�_�PfX�z2�N\�kg�1�WD��Eyq�T��!7Y��`��
��ܣ����
¯i5�<lJ�G|�UH��	�&*�n�(� j��ChK5�_�5]����VWB��Q�ą��/���o�[�A�����%ƩD!;3ڡ���E_�Wb�tn`�]��Ǐ�>�###�8;+�.Ι��������·[� �j��S�=!�U@���_�f������V+��8��j}Q;��T�cP��)י]�S�	+��,�@� 7&; *�
ei���9v�
���j꣔g�;���ęJ�H�R�\Ks�1�ąM`�Dhʽ)+� ��F&�;lƿ�|�o�
%ˎM�ߧ|���t����W��w���3�jˢ�g~F��<;�5����|�� :,^�7�~\���F�5��p�&���.{���f�3�a�-Qqs+
�H�d��5�j��
�>��`c��m�+o_�0	ʨ��ni�K/S�?sE ����:7UͺƳjj����y1)���V�,��Y��٨�RRR{�ϨE�{PAz�?�<��P���D�X�#�(��q��;QMI���v�� �X�ڂv��� -��j��w�-�җ?���K����rF�sY���_i��n�\�ڷ���u7�w?��I��[�~���t��1���݅�v�V;��P�?�_�ԹT����M&�(�E,�"y��w��E��U6�� 4�ȱk�{0k8Q����V#�����WεE�5Z��W3R��ڛ��_�^�
7n:u�/ �R>2"lj|k��쨤h���b� ؜QSb?�v5 ��>��;&����x�~A;ِ	�S�~4�}�C���@�sG;��э�PcGǝ���35�]-����ӻg��я��a�;��{����ƚ7�<� �#��m��fo��tDTTvEE�PHbé�����h�C�e��掑���;���2��ўZX�2�7����ٳ@�NL�q�6��rU5���c]x�~�2�'���l�b��镋ўk9�M<2-5�bMr��e���Jƛ�>������˒���y�J����9O�Y��ȞW`��!��Q����Z��_��;�ʁ4/�S5L����{�1mȷu�8��]�"�S


/���%����>��m?G��5�}o��Js�H�SƮ���:���?��ey��̦�.0~���I\�����ɩ�����78b����hk+����F"��*��cV���HRRa���?���%�� ���t��h���$�:��H�������Z$9wWJ/��\{�G�+j	v�d�� ���*g�غv鞿j��*�h����V�@�8Ea*ٳ�gu��?6�n�O�O�;::�f�e��w7��6b
�Y-��G���C��	��v����x��K�n��UU�vɯoN$����kG��~� A� �Ĕ1;[[�;��;�T��ʤn��'����ʺr�F�X׫:���x���tΟd�������.��~�{l��l�=��$�����ҿ]I�U���&�̉~��V�9���^������`R1uS\�����x����fff�Ǯ���L���"18y��4"��.M������%���ˁ����)f�X_�ߪ���9PZR���<?����[���YS�4
o���;;?���q�M�8�̧׋T�y$;8:�?;̫���P��h�ԥ5�F������|��w{?��������՚)9�\������Lܕ���EFR��/��z�鎂"v�H�����z{{��mm'��2.;ű�D?���TSS�a��ID�FNrh���0��_&�3�)�����9�[T��\~�~e�A�������ճ�6�<�X\�� ��������~��+++*�^�S����k����b���]����[���dx{{g����`�����/_ڧ��E��ʿ211�E���}�c������"��! m��;����&��I�Y\��ot\eP�����\Gg�+��x�G;x06�aø������Zz&_�&V�Ԩ���H�;��S�H������1���%�����]�Ȉ岴����h��c��ס�\���Y��㳓!�Ԩ1�����f�/jd��>��N pE�NqswX�O���.LMoz�|,v$�	m�A��"v ��YI�P薔�f֨��M��I�!�
���Y�m}�"'�$���������ynq���ak�Q�_���p��WLe�����hhh4�s�u�UL�NPH����O�P��ˠ6v���FS� �;������I
�K�`���x���mY�hSɃj7m��7o�\��R<��;���NO�`�LC��
����e _�D��S��h�-��Q�y�NIRA!�}��*RSS���j��aB|��3g�8��9!*?�1�C����F`��Й �9�:9P���|�PҠ���.�2�� z���O���p&�u	�o��k�������������
�-�@�ONN�Y����cgg�+b��5�u�1��\���������;��AR�	�A���ZZZ��`�F0>���5%9�Bw�a0�\�⨧בI��_������`��~� ���x�,�XzJ��";�\jw�P���!z��ӕ�(��"oaA�X�򢉟��'ii4��8=Y��f>{���&sy�%KG{����>د-�~��TQK8�2ޟ�VqE�.�m�&t�(�߳5����_U�$��` �%��Ɋ�8A�5t���S����z��������;0��a��f��pC��a��� ��l5�F�>�3/�� ��,A�D?��S�W� �����H8V��<��� ��CI�U�������YM	mO�'����ǐi������[��qq,�9�۟�Ė��e�(��k�7<����Q�,g���|�+Ն�����{����ERJJ�_d<���秅@S�r�T��1�2�&45��&4A^���i��qE|���#P"/_��*++��b___T�$7�`���6-��� ��(b�Q+�JK�, �c�F��cK���2����;r�K��F��B�_��'6_���� R����I�UU�����EA�ei�ȭ|4����Y�봋���tZr� P�M�<�&�r.l~&�"���)���&&�v�/��Y��3�
���_�x߿�1=�0!M	��������|�xh]�Ǳ�.�x�v�'qtO?mJ�-�|rH����9�RuQ��)�!�+PM=�����1���h�kl��4��uS� ��#�\\���q�c�y:�Yԡv9����B����e��`0��JO�|�Q�����+���k H��O�@�h5܄�+��Ç0�?��NHK���jS9Li��)�Oq��Y���w�q|a���p��R�{sNP�i����� �g|���:�CE�\Md�g��]���0{Q���V��)�s�da���vU���u'� �XF=?5%�����+�侥�A� ��MZ����
:k�=�i���!t���H�R

��5qo<� a|��4 &n�@$J��w�Ґ7莰ބ&����ؒ��� \�;���6�6����X���ل������ƺ���'$$X��j'�=�#k�_���*y0�cZ�ӧO�����D��uv�~q*�Y�-ѡ��$J��sss�-���;�yM�Q2�BM�FFF�>���q��b��u�-���n	xp;(�M榦�� ����~��3!���.>,�ԧNA��b��=��W�X��'< ȫ-����a�!�
�
�"���Է�xyy_��l���䢣���> � @귾�Zd_��/x�˩�j����vJJqN����mG���~b�X}��R{o��ϸHuk㧮���r��B&�i�����(�4:#���=ҺR������~'����3l��b1H l`�b��c�^��s�:Н¾���ﻎ��TF��^��Q����m͚r@�@����<��h�eē����.����*�~�aB@A��EM�4����p��*9ɀ���D�Sp�83�A�r�Y:v�lo\�s.�ڲ��7.���Z�V��IP�='�6!*�ӕ���M��*s@8�W%@��Y������\d)�5d=��jVu���ŋK+�����\�j�(B��^__�z�uĊ��|��['}B�����w:`���
��Q �\��L a_�-�*��]bR�ޤ�� ݀Y���QO04^�V�z����XZ�������K������P��O#�?��%4%�~�ɼ� \㯱NɣBw
��~��v����X���m����F��m���;�Φq����� ��K�ݤ���oV
.�z�-%�߯^�� �.J�ռ߮OVi�n5��j\��J�,���&�ӪDB���}�	�d�U;!~�3�x�E�#q�kk���� {�}��fT� Tt�N����g�DMZ�ݞW��ߋ��M�6�]��
�P���њ�[��6`��K�ѿEoU�QŔ�]�c(�b�iaT������{[EM��iS���^�����U0�ʗ�Z �`;�N?�����^��ɓ�j=�su� lTy�ed��靉p��ē���e���L�Nk�DW�ŷ�j&�Љ�3�)Obo���N%{�F|������I$��N�WC����-ܐ��)��^0�o���MP]�6�s�hR��4��-j �`��4���;FO�N�n�3����(�3��D���53�wjJ���۫*�AhAEɚK��-Pb���Ф��"�������!@DjHLLL\���~I*�(IK�@b �D���iy��^�]:���A�T~UUUN򷻥&;f��+D�u1����qj��/	������"ٳU�@�N�T�vV W���PB����<�;�Trg�����?�3/]���qF���o_�|9I�� Ǟ��@_6-iJ���Mk��;��L"�5��(Oh��m��\9;� �.@�hKx<�Uմ�V\��j����<t�P���\��Gy��#��}kft�+'�������
D-+v���uc�9(�s�,O߇���2����f=G���.0&
��� �����_gń�%�=��D�^�<CήM��t�h)Խ\����G��<H<��������"k0�#��T�޼݁�����x`�̼��E��#=Ӓ����k�Y�6 �@-��ń�j�T�	vw��8%ew�ƹ�dPO���N������K�Ɛ)�mN@�UH`x�����zx�^)���4G_��X1%Ya�	��ۜ��C�L�R�a.7��)�T�����P����u�D*,�|QUQQa��	um�X�?��C�n�z
���z-e����H��P����T��({�z�MW.<��}i�2@�3�-�3c�Ы �Z�"�}��y:/����#��ʊ
���t��мV����������ԫ�F�[�	>=m�R�7�����sL!z�{k`J)�T��p��X �R�����������;���`s�a�E�^�+�]䕽������L����1)g����I���k�j��Ih@'E.�ZZ�Z�+��x���1�.)]9�.���?�LRڨ�OP�HyG�+�w�~C��@ *Gh0��
d{2	�Y�HV���t�N��V�|�^A֪��K��G&����W�̀��|�v��{����44rY7�a(x߉q�~���O�)�?�T2I�����.{TH�S�x����[[�&��XGʯUg<��)b�� *şj�.*�4a?Z��/���ʙ*�������������m�
dP�����p��y>"2�!�ѱ��r�l i�~��y`HEU��6�������]�}��vJp8�������#��3� ZЦMD�&1�NY����d�~k�Q��t�v���U��k!�A��x���nB*rR��xd��
���s"��V��Տp�f�>����D�u�� ������J����67�}�U�e��)gbV�l��(�M/ٖ66g#��C� ��c���x���n���9���ꛌ�>�q��G�vvh/+I$c.����

�}�:C��0;� �n�	��?��m��SKM���y� �[W�׳ �zu&�PX��r���`N"�詩��..��zZဏ$i덅n���ɨx�(Z��x2E�s֚I^�h�&�I;#����ј�Ud/M����͍��)�E�^�F���K�GKS�r.`wKY���Q�z�h{��?ۛ�@&��줜Q�ܖ��D+¯���fg�
�}*SRZ� �"1M	<wK���~v�6�7u������џ}U���СL@_U�iv�/<���j�|Dp�-j<]�>s {(
6@e��)R(�

�*��@�����B���j�,0ߡ��H`y������)(�v\||�:|���R�� �R �6�=ڴ9�y�����'$X�]�j5�	���јN��2]��Ӫ�s*pp=���8
i��H z⛣�iK���?���hV������<8i*
���Ot��ݤ/�	�m��d�FT�7�|#�ٙ�@�`v��Y9�	Í=��oۻrѢ&O�h	\���tM]������NHS�42-9Y��ԅO��C��D"N�єf	K@ ��T��0l�����mq�ͥJ�t�A��	TolG+(���q�`��p�Q��=.	���&� ^.��vJi-��@�����u՜n�K���ъ���J���c��U��q������c���Rv���?��ݸd�M�\Ԣ��vŦ9�⊻�[d2.>��f�׮M��F�ܧ�n津���鎶��v	�s.�*(�*�oo|~Ɔ�	�5�-�U�I�z$M-�<)1 ��W)2VѴn]Yh��4��������u�pÿ�h���	����n��'�	E�)-��{i��m��<9�]�->ƭM�0�@]�򰵷?�Xw7��A�����wT^����A�L@��j�٢��y��6X���{Y�8;���2h9�����	P־>���;�w#T
�"�%遦��xW�S��x6�?�{w2�l�w4�V����H�=JBE����3��S$���S���כ�ii:r�4�*e�&bC��u�"v��U�Ϛ���]coӢ���q�ߝ�)c9p�+:\�?z�YC���z� J��e߼����|��0�v�3)�O�PO#����[Z&p��P�SR�kH��?L�h=�Z�ftr�"�������V��:m"���x<W�a���n�QO�ɹ"/��+)�
j�����PC�s�zfN����f��x&u)��<��	%vo)�������H<�
]��q���ǿq���&Q��l R)���������\��Y��K��)�A(A�}��Q�����ed����B��=��a�� �K�P�m���!j��=���#��_+C�!oB�����If�٠��6֐[UUU]W������T67��m����$��߄�E�qvIU�MO��0h��b�@͡/���:����w0	[�4����~Aql)u��\��_�
hh�H������P�9;kV�b2b�i�%I�m%K�([U1��쫮V����^8�hB�l3�E=��!0���K��A�4�����D!����c�T#���kk;D�Bm:�*g����Q�VI�<U`�ڔnӺ�d+;�aN.��Ɔi�~g���l�'�f�;U"��{�G�);3�i�������E5�.@Y�ZF�!����+>�Ua���\!�����.�t���n�:�#w�`�U[�T�5�J�
���y�0��
y����w���#n��׷�sS���(C��Wa�k
w,��x"Q0C$R������e}��a��t�U��a��0)���r3A=���p� ���������3%���ǽ��r �����
�Hs�f�����j���{V��F��&{}��1+pG�%���)j���i�f󈊛������hhf�'�î(���Kç��j͟�'����D|ᬋu���JjJp,�/Z2�#6�u|��u�>� ����3!B|�s�R���o
���:�4� �ՋG�-*�����ҩ�ɵM�P�Vx�E��=�ǖ5::��������tZGzד�_���f�ץ?\����KEc�3���>���t���~?�@]�gG�% {�ڄL(G�����ͩ�/S�>J��B�P?�(����g����>���*����H ��K5�eZH.TRCI<��?� es�6�T�h=x��O=-`���P�$;���"�ZGh& Vq>:krr�3����4�5%�`��漦�r����E����r%�gX_��Bo>�	�[����utosD ��=r�E�����8��l���O05M�UK�!���� )IH������@\}�Dгo���W�Sk�5DP��̅�&[�8�X������f?�< �x�~�ኴt��t� ��/g����:�䰣�s�O�$��h���BB�fP��� a��s���>�7����9��Ik�J���A�9��Ki0:gڞ� ��)�C�����u�c���/����`�w,ꯆ�އ��a���8|�.C��\{�ਛR|#�Ro�fNP�MZ�?��FYk\�:����p,�=�ʹx����|ؘ��qK�Ԉr�bŮ�(���'���u�o]b_����g�� �8�%�/r0Q+�p���i�����غY�?��\�L���a��������Y�{���o�kE�����.؈��rZ�!#�DV^^��0�$a�7�[���F�d�$ K�;$N:B�R�Vοn���PK   �X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   ��X�Rr5�  5 /   images/d5704fd0-3deb-4692-9952-d29401de32f9.png�gXSY�6@���c!��cE&�;l���ҕ�*EzO�(�t,�����
J�*5Ajh	5��Cq�yH��~|��o�./=g��ֺ�{����g�_����)�	����9}Bc��`�>q������ ��f��W]`0�S�o���a�=�3'�/yƎ�pe�00ٿ�ڴ��E�=��͏;����1SV6�[��`���9��w~�K�*�%�6׈�Ǚ#Q#�˿�Mi~?���u�Y}��!�+�~"|P���%�1[�ߊ{��}�z�|�/�?�X�~W�@z�3f����jC�?m����q�9���?h�lĻ�;x{/��YBS�"f�uF����C�<���p_�y'7|ÝWj��x���3M��#t�R��s����W&�j�0�pKb`��/{\y�T������;�g^u/��*Z�~��n��M��JH �h{�;*"�t9d
9\�fMϚ�ċ��#��.�]'o�&&E�F���MܓꝨ������8�➣�ϟ��X�g>�1��W"b�������9��p��ut"���xx�+w���ȳ��!S�|��r,�����ʫ��Fp&���B���R���!F�$�}��K���!��N�����ӷ�U�$^f*�=;�	��n�X�w��r�ܟ�@ԅ�kW��O�ީA9���D'ԋ/����W�}�H]���ǉ�3�P"n���t��j8��ܕ�l���eȔ�ћ����=��L�6b�E�h%9���Þ��3w{������1�I-�v��,?�+&Fp�g��؊z
?|��AT���{v���!�*%����زkAf��ΛsK�f��*���-��O=�BRO���'�^�Iy�y��_�1K�/�6����`nkk��1�	���Έ�8��8		��U$�1�hk��v6�M���9׆�<TI�歈4���ѹnNZRQQ�v��V�k}�T�ӥ����،����y��+��:B�JO4�4d
]\PX~m��v���ޗ�W<2w��@ʯ��E�3tJ]b��3 <BnDv�L���QVA�*?��mV��oߜ�ܤ��7iL֗��bV�������O>�A� ����ۋg�����C(�����[�I-���
�a��=[��������=FVfO������l�R�e�F����2�^l|��W��\ �N��KOx+��M|�������C�Z��n�G�������-9�C`>�:ឰ[��q�a #;�233���C�s+��0���?��M�^�VV�ec�>��
)��sޥBR��.���8�Ԥ;�����魶y�9hu����<���=)�r}�ֆL��J���M�ܹ���3�����|)����3!�1�Qi&3#cpk���C�,B��`��!Khǫ�W��\�|�}=D'D���~�i���R2�H�r��"�Qc��D ��W)Y��O	�8O��$�8Drqq:C`P>싄T��c� �H���C���J�֬��zhxh�9����Ǥ��J�$Y���t��"|�]}���A����XoI�� QG*m�^'f�;�e��/V��2��у���
^(+I�|ǿ[*�\�	�)�<l"�����x%�*���,���Xߊ^�(����}�L�'o"�M�n��[1!U�����n��*>�eQ�U�o�-C�e�K�t5:Ӵ�3R��n-�.,�+�{X�ݐ����Xh��!i��-mH�G�9�q{#���s�K_���G �+��oQR� y�P<Y�4<<��<d�2��N�ݩ1rS$�wcfg]'<J�޽��q���鷅�s���(AQ���ǰ���q�X��/�ÇoR���UmV�zh�2L�6�iF
�`[��}�f�}"�d	�@w#������}w��&s�u��?E�]�����!�Jg#XU����48�Ю��o]��~m�"C�8���o�>����f��M+�#>~~�����J��n�j6H���#�hP��F����[��|<Mo~ u��;1�Z�����r�㵮�H�C��Q�J�zb�O��4\qr
b̥6���@����[�?�U���ë���[���i��S�����C�D�W�I-��]*�ADS��q-����ܛ���ɱ�3�4
�P�F@y�o��f��i���q��*�痨i���ϟ?�	���rV{�6��b�/�A�\��&����
6�J�[�)�<tOH���t_�n���t!Js��H��;AiD�*ixk�C6!y��ґ��j;�H�A���C�i�WIt�B���h;�+�W�#�#��<�;U%�^پ}�p�������KM���������l�M�gS���/���@jR��뮃tE���rvl9��Ձ�;w�<2���J�Z������} �I8�}���a���Jp�Uapz�y�S
�YgK���]Y;�I���U!�~� $��b�������$~u"��L�(�QM���@*^ �@%�|���VO�E�{q�K�&q�peUU�.1+�eH��ׯ�S[^�A����4a0��Ѷ�3Isss��I�����n�U��L��dû�O�K`
0�[~��Ͻ������Z\����3�J�C��ի߄cy^�a���5hp�v/$�һ���o1����3>~S̽4Kv�kHK��<����u�*��K{A��#U�,q�A��F�p_��/_�<b��)��yqG���l*7��!S9�|�3��M�Syyy��١�6y�Z�l�aY-p�9��(�c�Pu/P���a����o���:>�Y)5��+�����Ӭwi����{Q��7'v��:+
�`��e��I����h;���q���bR���ה8��h�8��Zx�2#;�@{VR�|L�TJ���ϰ��;�`����/�,(ƓwNӅe���.�������zw'��F�@�]����&�п�E��K��bYk�m�=o$~�v����Z���|	̙_4(l��]P�gzf(�5O��]sp�<A��_+޿`y��mb[�Ļ@�H������1?�Y��xC�T�8I�{����j���V|jii��"p�Am-����`�73�e�M�5Gr�k��)װC�(q�AZ(���IF��X?�����ڦ���ߛ�znF��|�T�jm)/݅(��oPRk�ǹR�)��-�.�m.�N[��0
����3�}�3��SS�S���sR������������Ġ��x...�q|暰|�m���b��� i�@�ZE�$��T\�}m&�յ~`�/��؎��[K��HB�����6I)O����[a� �fW�9X֥��?�K-�0��(voKB�C�fa�R�¢"�Q����X4-��/�AFs&d������Oi,N�����q0vA�[S�A7@��������p����T�Յ�'>��<�%����	�5G����@�^��簠�Ck��R�ხ{qϩ/�&��ri��A��A����o��Z��A�����e���t��U�Ty7}]"�d���%E�S$�%�� ��ڦ2{ %pC��y��d�ɓt��x�q .��L0�sw���>�I��ܥ!��2���s_�{����Z���!y
��c��d��v�TO!�(#�?~���q�ѭI�[�6�L�ي��x�[�2���fп�)�y��(|*ۼohx8�A�{k��B�H�3 ���ݢ��^>mJ-���n*�O�����!	u �&�8�ꪑQ�nkF3�Oy��bV��|���w)��]!$^W��_�ے�x�Sm�����ʈw:h[�q��-�d���4�c�ǌ+��XI>v6 s�>	��S�!��,?��B��'� 'ȴ�@W�3����?¨W�"ˎ-a3�6^��i/��+M��O ߟ�,��^��A`�&@{�d���]/��*$�����z$D<*y��Y�]ւӭH(qy#�)8'M�`&s�,��s8����ȐY�?텽�cz�@�T�'�PO?�N���da肝��Ŵ����SS]t�L���,�_u�ЏԳ����e������rM��f�!"����L�~dd�{��ٱ�լ�N- �gK�Ր�$v?|���ݔߤJmVUn�9���T�j٘	�7�n���c��~�[x=�����P���0{�g\�niS{$<�e��|Vv0~L�����Q���]^ᯥ��:�Ra�T��5��2x�"n���9�LU�cuʦ�eQR��(��?�J]ȗ8B��Q��]mZe�nVQ�F��ֺNj7�c�!��,$�4��H��ߕ�0òw�2{&�)	Ԏ�`��T�J7D��������A���(���G��HH��f�ڙ�/*DxvԘ� 7G���B`�w�^ñ#��ުQ�QȞ1S�=Ȇ��.������t�t����|���)��2��݈� ��8�8oEi!ߞ�q~c��g����:�EJl�}���~I
w{���٬����F5�E�T���ʐ:8dԬW*�c�j���j{�3��'��M�j`�cY!e`��|��L����y��ל���Z��U���VnOCc�:��p~����4hֳV�@��{��Mf��& :��h�Ε��B║a������O#x<��O�w���TZ�������p(yf�l�P�X϶��`���A�3U�I ��:NX;���W�k���f�̓��Ntip��(�/��<���S-(�
��>`�N����R\xo��US�T_���d����FPd<�-��zA������e�Dv�O�N>�/���iS����O?�aV[
�Oŗ��DY��Y�_6�1���O�<�E��ւ��ؠ2�[���4ogI�ߖW3Q4U�O�;�-�����b�t��Hp��r��Q3RQ�3
�]9虙�%Z��*p��3�B��S�
��@����!aaR�q�0K�&_��f�׳}��|!V�K��M���1�K��!�HR�VL�f��̯�(&�ίS�eJG����JFNJ�R'=x\U��M<n$�9��ms��N��N<ם��S$�Rh-aI��xb[���:�+�� �za�����ê��*���i�ղ�x-f��w��t��MX�$�`�L�Թ*?�(wJ�,R���s;$�e�qr������
Y�^�s��Y����G�=�]"���2e�]�j��������z��.��@��p�l&��SC����q�
M���V�g��I��� �^�E��jF����#[aV�*Z^�l��8��v&}�I��	�� Z&p�f��L�\��̖��7m�h^O5Ͱ�Ɨ���M�Sq�G���Ŭ� y:4�ߘ���En7�������FIkf�l�<������\�;�Bv]��[������G7|^���J`g�.	K�ӟD��8q�x���T�-��w+:��-+K̊��D �J�J�|��0�@ufP�,�?ڈO(\�,��Zȧ�c�gT��ʖ��^��[w�a�K�{dvB��u��E�Y�O�X��\Di�:�n:w�ɗ��ʞ���֖����O��H�/���
�|y�b?��J�hp��Hh�@?����,��>ګJrQ5�7;H�w����9.'S��hs��1g�"T(�q/�Ka#�e�I�֬@��@� �ݫ���n2ȇ&A%��v��]��f~�i-ٞ?�d����x˱)����G�����D�9T�i2U��l��9�Ւ��^ \3m�4�'�7=�2��\�R^���6Z�,o�*9P���1���Hq���y�^�d3_D�'Ee�kQ��㚜�.���:��v��8�M����Vh�B��R�M)���;�U�W���u�9���]�l�=g�IɎXD/�Ӽ[Xi�"�DX����5G�\�!s��K��:@�$�fޢ�Σv`��y�!rӋl�{c��o�t�c2+1m[ޑ 'I�U-�k��6���wM����iR1�гFUI�MXC��5P��N3Q �}>/U���X4K��K��	�h��&�� ��v뢀ڲ��@�]�Y8��0)��-f�Z�V�����E#i��&g�{_�]Y��Rq�z�{l"����!�d����ʈ�~c	�i���oIO��`e�Yy2�ɪ�n7n����̳_�
?O�T��5(7��?�2��X��E�ٌ�a��]���93� oS��(���ń!)�̞��u���Cm���%V
:v���&=��%7����'y `f�1�z[j��e�}FscЛ��M}�����V\��Դ������d���˚&%f�ӑ���a䲎H��b��w.�̯�F�$�q�$�yϔuQ��b(4��C��dU"��
�b��R�����sr�q��V��7��?W'���s�ϟ�'Q��Bc�bckU��fkkCV��u��wx��XA`:���Q5����gEbM)?�"�&]¼��]]��PVmE_��i&Eh�n�"a[V���'%�/zU	yD���I�CIn�\YG����Ls	�49{Gc{h�E��2��(��n����x�����!�5���.��s{/��n���p"cϪ��͐~����C��
B���<?��~�kW�x���ny=\+�r�(zxM}s�CP:�ϛ�������KK��2��b!�O9ҏ�p-�AξQ͹��|t���j�<�tF�q ?�.q����a-�sJT������kB�͟g�}��K��A��[�3���J�
H5,����M�=J��4�$N\��L����rT�w������zj��2�)�r�/u���eg7�u�1��ng��\7�`U	'|+%[#�
aD�]W�,#���K C�;09�~k^�����>Lc��H�n���ޙj�������Q��1�EV��7	y�Hl��x�W�i$�}x��՚�$����TeÊ/��M�!K�n�:ơ���"�
���Jm��#�1�~�p�@�b��cR�X�X8��._ҡ|։Y&�% ��|k������lǄ{��};Zm���疨��YV���x%`ɘ�f��BI˞r�,��/Jξ̤TӆX���e��q"T���B��u���[��o���D���Es���~V��k�ۦ@��>���Di�����	G��bl\���j�J�[픙�
�04�I�k���~��hX���x�|�i�ϒ�V	U��Ɂ`B0Y��X���Q��h���	%3��5�w�>57E9����j��B��S�cs��0T\t�P����˪|{=D�3�LҖ��c�0vZ{�߽!>i�8QLX��s�S[0�VH�����z���?knn�E��ץ�9�;��$�o�c�I����9�5��G��xצ3yx�z��������#y�Ǿ�y�n����kQr0+\������,���=�@9�z����_��r�l�6W��2?�ӻ0	W��ߪ�3}�***��y�w`|x���Ws�������hj�æo���\�:�����A!�SLm��;,BcmF�.]��!�/p>�dԚ?�#M��S��'�T���a��(O�g%{�'�S����U^���q蹅P9TsS53����ؒ���=b+�0�n�#T�$�*U�Q����Ȯv�n��ǜ)��Kh��r���P�����ٷ,��U�4n0Q,�	"=�_����&�������Z�U�a�3���-��_�og���3! �ǻQ���x���*w�?m+��=��v��҄�R�_d���Z'�2��q��T��m0ٝ�OJ�|���\�퓇"�4!�V@�-~���8ʅ*K��v�m�:�fl�7����6�PZ��|:2
G�I�.��Jrݚ�#Z�#��H��a������i�q�N-��z��e�$X�)�r_K�W�@�"�dz੎�����?�O�>W%�n��+�WL��=��q����%���Zʻ�BY��M?��ϙ�ϯ�O��m���t`J���p4��a�*�7ә�#�ݞ�<��1>�F�ULY�<�(+�� W.G��4��񚩓i�����=L�Z��287E'�Fhow/M�صkׇ=>`z4H�
A�/k�����X��i��#��b&#�,�Ͼ��-S�������~V���}6P�U�4(�w�ﺥz��֐sZs��֗��]!�%� �rrru��+P��	To[A�����\Z=�[A�D	�b�uW���(�6�O��md֋x����lմ��a�g�� $dp!r`wS$_����P*ݔ=.��?���y�w��w=�8��O
�ɩf�w�9����|��#Z#�Iw�k����m���J�I�-D�>(9M����Ip�S^��T�irz<�A�g�� <���_eJ�ٿi+�B`2��?��{����EgQR�l(�?��I_{�#VI�Xu4?P�奙	U��,���
��x,�d�<b���K�ӡ��D���1��;|ϻ�E�|����J������N��>smF�=-P�iKjvl�ó�>���G��4�q�̏S������ts2j��{Ks��N߉μ���~��
ٚ0�7"���+��o~�΋����^^���:��=��p��pyQ����^�ޢ��,�e��0Gi�]���N��� �_��M��&LG�D�;�4�`^�P�Y������h�[8���$��tx�2���YB���ԍ��f��U��<`�xt1��$ߣ?<i?�)�Xtn.~�7^c*�;N�Ñ)��Ս#�@P5~�6�X~���h�h�3b[��i����!RH�ZPB�{����lu��T�l�^C���R��9��+s��o��hYA�`�`��
:��}5��5G���C^7��J~�ی�(�ݞ^�>Ѕ%Ш���\q_/���`
9�. ��&�Wρr+Lq��o�މCS�Ķo��j�x��*#���a˥_�M��¤���/�fef!=�C��/sI��s�G{���s�s��{#���[a]?J�.��$l�a=�o��_����afg;����P>�4�1��g�Q	�]�ʳ�����F�{�8��`gg��Oȉ�,\0���Rv���wg����K�j�!D����-α��2Q��vg'!�������g�|�Iw�]w�[����7�|v��>c���\�f������h��Oފ�Ut���gNK[%(?y}ՙ�(�9aWCs�>h4-[J{�Sm�U�}N��f\{����p����	���a��L@h��j�uT��-'�W��,�y$��*���_��.S���x�lykq���d�b�X�4�V�?�'DF���|xA���c���H{�� �:�kb�"���{�[y^��;	��zXݬ�h_H�f����?�(�+vظ?��ך���Dn|��m���b��JRrE����4���S�������A�|�Ҭ��#2����T������*+�E۫f&^��
B�XVr�m\�L�*ѿ ay6%���K�bUg{�Vqn�^��QVfT�Zs&��9z�[gU�����é��c���S�J����
jw�uJ=�-Sfjt�}��~"�M�w�0�S�r��X�r�t���U����\5]�aJ��){TY��oN�n".`�+4p7e]��!$�����0���3��$���}bm��EϪtU`vF�.Wn���9ӎV��`�;{�﯅�?P��
��^]��4x��T#�>�L�U�c]��o�w&	�G*z�A�I�B�����bWt�XO8��9�,?��*WMU�Ȓ��'߾F�z�{U�N�����A����s��۸ڹW�Y@��jy��*m���d��������YXC�d�v�Bs�r7B���:b@���}��I"��?-���Mޟz��,���ݱc[q!��󷽃��A��&K�:~�^y��0��zT��cx�&�<a�i%�+qc�.�m�-e��|<	b֕�@yDAg�
X�_~OqM��p�t�N��c?���_�����!�eW����̯_�[���lpX��n��Y� +�z7E؝U�*�V�ʷk�Lh�7��:�E�&���"x+�&b��T%U�Rbx-��Br�?�p_���K��,$�|@���1�0F�=�Χlا�y�/��Q�g��5���d*�~���O�J:�ޥ�ث��S���ga���4�#���� �J�]�*	�����gj�1e~�;���e�����P-�������NE���ϟ�"8q�Z���
q��##���F�C�y��T�8��"D���Kw�����ذ��b{��O۷9|[8s,u�[۔	�P�Vib����Z;�;?um;��B!A���=#Y�*7�0c�E�2���{��d&�&գ����Y٭l��F�<C4Ԃ�!�gt9�׻|@���K�{�|�>nZ���FZ�ު�<��M����S������HN|���S:ZZ�����J��D�m�������X��%��Zh�(-��[� �$�,L��q��a�Eno�'M�A����r%�/_�Pa�����X��,���14�z�L��_	3�
GBc�9�}�2���S���؉y䠗��/0P'��YS�y�@�΋��W�����b��qc0�*>
R�3n��S�W���%?�{�o��	�p`��|dlaa��V�Ԭ�)E��t��_]��P(-hڊr��S��7.��i^�*9�:%�2��N�"nmSn�58躻����ܺ����.&�-�Țz@�e�^Nl�=vâuv6ׄ�S���	����n�;��ϲ��I�����3����O,~�r�"�#�ڮ��N`��}�I����8�*<u�L���U7�S^�j-���9a�2�A�����si�Ж�T%�jֵW��
��������֛lWf��9�T#����%�$���za��)֊OG�\�h끌n�>�r4M���W�׻5�c�l��u[���w>�}-����=(GX¤O�������W��ڜ������<�S��ڌ|���Z�����#�B#o�e������v�k��7S��|]XȂ�%�,R2H��r�@��^[���l�� T�����n���b��U�y�7����O�q�
�׷�+q��aD�w��^��C�w-�	��9�X��§4�����s6L�&v����[Aj�u0�w�eV	��ʆ�.��X0d8/FV��,�<��L��E�.w}�ڜ,f�k�!fM1�_�܃�2��Ҋ�fQ��t�5��d�ن�s2��.T�5M
4�m� �6�RP��Ջ{��llR����ŗ>n��� ��;���f���-�1��K������|�y1�(�����z�31�S���1b}��|�@�����V`���ֺ��`�KG�o�@(�X�F�I�U�Y�)F��F<��`BX�j.Xq��>�B��f��=�<��Ԋ�_@����i�L�uK��6���p�]ߝs��՛��7�x��i�!'�RjJx��%����Zg�2&��.g������VffZ���}lBB��_oaw�4�^xg�Tb��Eh�I���E�Ů&���cZ���C�i��\��+R��+��p�����h�����i�}�J�Z��C~a�D�����R�N��A�����Χ4�=,,,:������]^���1e����D�v�ι����=�α���%�����`;�=��V��5C�V�m�oo�Wi��ko�f%CW� `�P�B�r(���I�o�a�ݿ>g�"0|�s��d��Fd[W���V.m/�]�wh4Rt��R�����A��ެ�r��l�߯�U3-a	�'�B����RSS���������}��uQ�^���cc&���ס�4 .�.Y֝w�����(X�!���L�5�����Ֆنd��w]
 ��?��f���,t���R ��}=/+�Ɖ3#��I	����k/����q�Y���Vݜ�5��X�D�RN��|g����|�_�'k���1K�F0�zi)���i�ӻ����J��xv�eO��M���[ <�S���!�M�ϸ�f��)�M�����=+oy�}�$���9#���γ,^�]ap3�1�ݔQ&�t�q�_>�: 6%L%f��<#�c U���\��`#��CkA�lV�x̲8��%7������"�/��mϦ%�հ������}�.���\� 0d3����'?tp�%P�hk�=��7[K�S���,��O�R��RpO�
����� ��˥�|~9X���;;��$�����R9H���z�{@;B�\����<���P�up�O� _�,��v�Sܻ�&��5��LL�fH�n�� \#�)���y#��n�@���gIY�z1��|I_���ye�h�}(ZǾ�w����y˯#D��H#E�A�&�%z�k��''�l�2歐2�	��&���-8ǒ�Jg��Kc�~a�c5
�o1k�7���!����%��?js�*�n�����I/[āMD#��۷?]y��~Lk�D��q7Z�R��$q�׷Ma�@pM@��U�����!���xJ�~���,��;j���:�����PM��MS8k� ����ۅV��Y��x8qm��E*FN� �(d� p�h��vG4�P���J��S�Rq���yUx���UV��Y0�r�`�~�5>h�\L� �~��� �1��5H�A���h��J�P[��\����L�B��3�+4ӱg�o�+���d\hKt`I���~q�z�u55�e��-��8�J �����:V"���?ȍA&��2�v��i/6��Mh�E�pU ��_9��do�i�Un<�n��	��؈� n��*����V�L<�B�G���NǗ�=��[��v��Պ�!;���p�:�Pٟ�P(x�l��K�7<�����i�
0���:�֞�}�{���h�7G_�l�Hg��?�dE��Ç��6o;��qs�k%�Uj��Jom}~�-�]ɱ��69%ki���º��Ɵ�.z1�(�_Uç���>�F�Z�W�#��T�G�UXqa�Ǩ�����͠�r=�8FxT"YZZ
�n������?&������Y=�A��	9��던��:�ʬ��/ �:�q߰�5;ui��g���5w�����&��UI���w|�"�n�&u?|��,���)++KV��5��v��g�{+�(��a��[�M��r����I�_���CP����M��|��"�3UC!�$v�^i�5��7.v�(�SI�c<�����$���rb�A��w7Re5`hi�`|1��O��V^�pl\��Õs)�n@R���:��<��B�QD�̪K�?mt�G�k�oq���65��C�vJ6p���+�x :;8+[mr��C�3P$<B�_	��r�MD�Jha39a/C �[�b���
敞�$�*@�v�nn��bC�}�������s����8�Ř���<Z��q�R�]݃�� E��脘A��d1æ�G������8�W�U9В��vv(���Q�@RI/d�w����>m���Mp�$��֦0�_e�1�Yx�jk)=r�ު���[�J#�Bk��ur?�Ņ�Y=IT�'�`C7�s�]||U���[u�hk�T��ֆ�g�c"���Zn"���[�0`j�/2Z+_��uE8�fx�&+@H��d'��u��M�y�����8#�z�N��SM���'�L��E���0_ ��Q�3I;���Ҟ]�ګ���,���U�χ�T�V��ŋ9V7�s�W-4���w>��	���L�Nq���-�1*�k��614x�B@*z�hY�`;�j �砉�4� �Y4��U"����NtHKéu�o��i"�?v0RCr1��)q�{�ެѱ�b��.���2%U�3�0�#��f����5M.���S� �v�}�.Ũ_��_�E���B���� �W�h,͛U#;t�xW�> '���nD���V.���jj���_�EQJ>|���ʜ�
(��|\v��2H�'�2�PV�0&�f`KO3��s�K綗����A^����_CϦ�N>�Ry��>-[m��nݚ2��Qz�	��/��E|",��:T�	���}(�|q�$}��f��U����aЁ�<��	��gϞ�F���1��,d{� P�ak����B�`/�8�"��o��������:V�� h�d<Њ~���8�zl�"�ZLh0�e�Mo����{ȈW EDGE-����������>}�F��J��E0[�ѐ��w�tGH���)[K�i=��p;
J�~6���#A<Zɱ!��~��6��Br�fC����G��<Zꘓ��@�?�͐)#F�7g����S�r��� Lʒ2�r2P�	I8n�����N5�E�O�%
���D(�=#sm��%h��O���ww>!�9�Jg�h<�9�YU��Q����-����m�>pW���,M�bt2)�����T�AVV$��I"���H��y�� �����~'�NWd~\B-����A
c�.p��onbԤJ`˯�6��ʮT��`�ʊ����nm�׽ks;r�Uc�wQȝ��eQ�R�^� �a��@mZ�Ǐ22 ���f�4%�����9���s.Dg,�IjW=�498B��|gy��/gv����}�%$iuׄĻw�@Ƽc���O��#�v�*¹w|�)���O8�|�2**���^���� ��9L2	����s�'ԗb�[������L ��t���m�Ɋ[�;~S��E�h���!�}�����JY�Pk�z�/����Y[D)g8��t�0jJ���a���B�<��#9�]�~�2���q��G��U�gQN��~���I
P����V�s��=�h�b`��Z-�*��'�)�0p暫��;1��P���gc&w�����k�������p��Y9<�g��ۆ�i$ZOo%�� ٩:))	�a��(���;�Èn6~��C_m����Nw��Y��8�����!�&��]�G$$d��F>�cM�pd{��^F�W����5�zԞ�cd�>̞Ԁ�y1�e���P���Ǐ�N�ǭ՜@�3@�R(���|5r�W\96�����>��;g@�����b���z��.Z�����!�J#hR���^:1i��ō����kA$g׫H��YD6�
��p�D��=*�ZD^��N'�0�ݲ[�`�_�Ɂ����6o%wtt@ (j{�����KX�{ 1�f�V&_�hG���ȩ�m�]�~�c�0[�Mr���������Z��r��i���_��vHLc���/|!z�1��+�1!R�S�1�M�
x�`q��<�������h���j��l���uQ@+:�ʛf|Ĺs�V��������[��ϝ@U��:�YP�M�m�������P�pR	����C��*�%?�m���AKG��0N|-�;8wlHj�[8q�mm2��� 	JII�mLUKL�l�al�>6"(ʹ��M���\�`h�Q���-��C@+1̀����.f���)KM���:P;0�e � *}I2����9`��n����xP��Y�\��:r�c���	���.��<9��M�
���0��얕��cW���՝s gmሥ���6���-���� 1���V"�/�mY���_�Í@�&�w<U��ܳ�/���b�3c{"a�7n$��Crઐ����tƞ��'+��1������O�lW�v���q�P54G�CƁz�B�>��1����a�o"�m��,��
�BJ�N�Z��JS���|�T<Dֆ�:�'$<�μ�{7tl�wz\Mۅ�Nw������5cD�J�Jb�62� `�f�ՠ���J�*�2��R��m�f��Ӷ:)�2.��s�	�D�=� �OA�?PO�6ܰE�I	�O�t�f���w<F����e�e=J{�`	��2�geiY=7�V��{��V����SV��y�ӌY�_�|95���5�4���{3��x�N�6���!�#5j{@%ܭ�³!)����5u^��wE�~�+_��������C�9��9}��J�(�z�S�����q���*�j�W���\�#X�;��˿�l}w?4�}� A�nSt>5">{#Ѻz+y,�xr�����,ݏQR�KHDf�C~������n������n�-y���F�&�����ˮ%�����daR��ųsO@�	���\���_�8_4A��0L����!ن����E�����? e�=�{b#�=X������P!���ǰ��,��I�ٿ]��XT�fgg?�T�<��a�ʠ� �.}Y�r�6��R[������CI �z�^=/=�������h��$���߭첲x?�#�ːWz�lT�,���y^v��(���\���SyI��9�ak�-�4W5���G,d@����Es��'�y�ůQ��ړ��@��p�N�&w�~.-�=a��.ʊ�&`&.u�쇈f�+���(�?~��U�Y�t�@;IF�����UǾ�e��I8�L�Hܦӈ����n.55�p���oXƀZ����2�:��܌
p�=W��o���I����𫃱܁	3sm��X���IVsgY��cS�R72g���j0� �O�p�]��ҫ�]XRR�g�iQT0Fc�����Hmmm�3dee�v���+`ԓ���쾬���|O`�"�"��^ۼ�/����LJ�v1o\�����������ԕ�'|� Uo3]�¯�@��ެY�.+˥�E �lލ}w���	�[��}�&��+����/�ۀ������I�=s��K��%f���<op˵k}$��>2��+C��v�c����i�BKY��R����>��	�9����8N�F5��8�?Ź�(6Ѭ�$x ���˱�
�>�XˣtJ?|��7�����J�^)Ֆ �ĉ���G�1������CI54��	q�������������B���o%�8�,T
:�S^@�t|f���8��w(V��Q��D\my �9�R��ح������k�OX����hK5���Β?1j�l�j]&��Kr�0�����v���ZĊQ���'4��8��=t�����2�L�ؼ�ƂN�tڤ5ϫ��o�{,f}�~�LW�Z˩G�:Tol�q�w*��+��tm�ݓ�Qۛ�������Sǜ�n;������|�ϯ�"�|������5) �gP�|�C�F�ǳ�V��Ro	�pDso�L���ZaR��!�ύ��P�/�_0�=�-�'�MY{z�|h�7�
��J[v;o�b=z�n��|`僉I�^�-������$�Z��A+�g��12t:G&�ƿx�@!϶U�v23�:�e��-Ӆn�'�l�l����jR/k�� �G�Yv�uX�w��<L��[�+�j�vT;��Pw׫܀%�Lv�B %X����ɏ6�	�`۱��r�����㡉����Wr�o@NV��~޲��|9��|I�u��Kw��rͅk!؁y�@�;�D�9qO��x�]_О���ej�>��^�f��Ce�Y��uZ�Y�N�z�~ {�1��D�!�m��OT�:�0�-�O}�:��`�*+�](���
�ﾔU{�a|�t���:�w����)g�oD������U(Z�5Q�����Ui��)?��G��k�~� !`;Q���F�K��d&�YAb�Ԗ��ă8Q���_�MD�2�X�}�՗�4`6{�ܤ�{x�A� �x�fkи��K_�fW5��'�_tI�y��i?�p�J�?ҁ=wJܺi�7ϳ�[sz2P,�U	`*a�@���	�8�<�pb�e颃������+�/�й���ZS�G�^�z�vb^�t�_��`߼���eq�ѳ+�/ج6��,�@����p����}���"a>�I5/�X��W���M�;�}��Y�1I���1�Ţ�vp>�7O<�Ϧ��1�ژi0��z���?��G���������c�l�/��G�����S��vڟ�⎯����Q��������9d���D^;�J�������|������<�o�kZ&�������_�/��K7�6B)�A[�/h讠����@�P���}��g�J- �^�B�6~͜�P�X�`9C�i���q3p��'þ�	e&�xb��2�߱37�p�Qt����كI�Џh�?e�j���Mm���ل���I_<�`�3saoV�h�e{�ɼ��]-O-W�����հ�0	ߝeb���vU	_>�]�2��8YL��:Z�G�gD�w'�� �c�o<�G�`a�u�xV���n�cYhe��s��r�:ߕ�|t3�וo:���U�wa���d~o�-���.ly���gWT��z.ݷ���6%��Lɇ|o��°)*3���Gc�iP9װ��#S	�2���V&QJ���Ut��kv`�[�����2ye����
�>q�>frYn3a�7���ٵgΖ$�sjM�)��2�u�늹����bK���yE�Y�-M*��^�*-�����k�/w����G���?_\�j��W�9�+#�k^s�:��K�Ŏ������#�]o��wP�e�����x����H��H�
]��u�k�|���#(�2N3 ��0�������Ҡ�����L��{�x���oܒ�rJ%���J5e��TR)�b�(��3�E%�i�u*E*[�)�mB�uƖ���e�>�g�,Α~�����������i�������z_�}���G���)��d���$10h���|�мM��v��9A!��Q�i���(V�7�^��ϣvYN�<��mڸ	!��s��4�.�	E�\<�dA��^H8�o�%�$P;۾Џ�OP��2L_�Oh.L���DJ{��c-���m)�+��f�)l���\�/k=��&P�P�W_aV��F~��K_�N(��´P�˸7�A����&)Y����6 �(��ͫ ��H�}��
ӹm2,�Y��9��H�}M`E ?TeZ(b��h������J�s)H�������p�b��X:p1�b�S˯\8��w��"	`�&ȸ2�q˧�o��P���Q�7�!�
�jQ�B����J?��B�N���ݤ�ϖ&�����X��/D[��y����:��ꍖ� �,�҇);%��%8`�;�����g�>}I�`�'9����N�ǀT���C�|�%��i2��@2m��3�ˎ S�f���&��G�B�	]I���k���mOd���S��3>�~��b�5���oTo�^8%S-����Ya�ԫ����D(2�~�
`������7���@I�G�Y�6}��`%��V*Ӟ�h>�(�=��P�N1�	_�A�ΐ����g�,L��]`��S��s|򣊸yH�eqA ���S;��~!�a�����29��0k�Zim�Ef���S�4 ��%����%~ZP$�b��T`��~5VZ�o�O|Ԏ��*0hC   ��ڝS̾�`q��hq�{K;���~�wp~�wp�o�'i�_�|�w����������������������������������������������������{��m
���s%�k�~Y���5�?���HCW!E���p�Q^4B6��������uGV~�@Q[<kUf�4G�3��s��6��iD�O~}�B���C�VJ7�H�bx��+P6�Sc#��C9�ъ(̋�Lg�t�h��FЇײ��^�����J�ݏa��\�Ջ�I$K�������TJg8��� ��=]9rY��^��x�@��N6���2Dxh����t�bΡ��v��xy�I�"Ngxe3��z�57�ч���>V��q���_?�41.����M��o�_���DD]V�tȶ���m$R_#c��¿l}bA �Y:���,�k��5���7��S��mo��(���5J��Y�U9�yb�*JR2�͜�,�p�~����س�dϽ�L�`��;HV�)L���SD=L�)u�\z���Ǯ�La_�H��%�ӑ�TZ��|)UPĥ�6w	��wiQ2.w���f|��X���$;��^��p�z�h'�?Xjϴ���D|�	�j�~~m��pL�a>���jė>�{��d��]3� ��|�6ᐇUX�2�9������-ԑD�S.��&c�B�43��GOM��̡w9�y��.P�p_�2)v�~��rťe���1�h����S��_<�߸�B�	��zǇ�rG�́�m�Xť��TN�E��q��D�$��R;��<2������	y���]7���K+m��# ~�5Ц�����%��>��[f�[w]W��~6k�s�O��n:S0_=�����N�2;'�˲�\���a�5��Hx|6��3��;+OmN�B�s yu>X�.1'j�]^|�ΰޯ,��8�����4�<�s�c�nw��(�ۺ�t� ���H���>-�4�L�sZ�I^������m�u�v��y�4���үc��^��x�na7g�sr8��T�w���������#5U:#vS�q�v��fAL���J�	� ���#6HN���m��ə�ϫNڕ�6��<}�mO;�_�����"���W���ե��h�p��٬�i�N0K��Oy�U(^
ao��h���k�|���T��ې-Kt���r����u���M��iYa���Æ�v�����X�Y����jrS�W��7̦��<

_���_�s��D�Y͆w ͜Μ���K�&S�!��۸L�{�i�����L�a��]���;V���	sl�=��4�u�9��Qng��2�����6�X�ι6�~
9Z?��j�ŚAt*�����6"���J��0XQ�c��'����������"���c�]gƻHb��ױo5O���o�5h�I�OIh�0*�����ϡ-<�~��	��2�o7t�$�nz��P�����EȊ��Lu����S#=�a{�j����L.1x%�J�����cǸ�z�j��>���1n���>p�&�UGU�~)�s���ʄ�u�Hq��M�@8����w��7uk1Z[ʵ��818 FY彌2��s�������j.�"u[[ͦA�%.�+�G@�;�+^���)������"O��рI��3\x=,��~5u��t�*DW�ϑ�=/��t�(�]����E׳��CJ�'�׃�c}L��ȿ"��3��ׇ����<�ZVH�ͪv_HvjŎ�*����I��Tck�}�� R��H��"7�qe`��x��S-�?�$:�a�Y������橫_�X�1ӶZ�g�OA�� ���9=�b}�Ž����ӿ��8~3`L�>�[A�0��e,���렞n���4�|C`��7.c�����4gNU.����b�V@5���%��?8�!S��$�@�D����~�Z��������^[P�$���Ϗ�o�w�G�ȫ�7�\~lԥ����/3�"|E�(�����K��@=� �׆�u�����=3�3'(��BE��)�d�m�S 6$�Ћ�M)# ����v�G�	_���:3��<_	q1k�_��8��P���#���S0���z��:J�j#�P�f�]$��r�ـ���ˡܠRfTZ'�_Dz�'v_��?�+���o�o̎��9�<*�˰/�B�uʸ���t:�H�V�i�FZR~p.hi��k�d�9�[����e�EA�ňA�p*\s���ݰ5�|�V5�J��K�|�8����"��#��B�Ǜ���a�4BsGoP�����"��_J�vm�@���N^-ř������<<T��}|�*˂^�@�9���vA>��ee�r�ELtF�fN|���Q& ��:��,�ǿ�DA~S ���Q�+��iw�ŉ���9�s}Į9%	s��]<l���� �B�E��/��$��*�q�-�9��a�� �ĥ��?T�@Wd&�����-�z!����X�chҙڄz�E�5@Ĥ�}p��ȋR����@
w�b�`웒�j�e�17�S��4��p��wegHF-f����*�@��o 5��@���`�*�o˻~x�n��5d�]�/d�.���i�X��ߣ���"
���jIWM;��K�O\ ���k*�T�K�sj:�p�,�%1v0R!�\�h��c�%��!�-�(mW�o��?A_SHṞ]���)�٥�/:>G�RP����rۆ6��=:|���x�U뵽h�jʫ��d��R4��ޗ�r��w�d4����Rr�;�zqQ�h���ה���T���Y5V��g&�=���qB�)��)|�i�j��8�Z�У���I�j �G�k/��v��ig6H��`�"3J��<��s�z݂��K���Ik�Z�I-=��,����]�!�����íq���`Y��F��Y�z}�ǽ���m�8O�gX�y�k���wf٠�=�II�,?�3
X\��˹�����H��$;tȰR^�vט�7!bbF�m=����囲�x@=o�	b#f�s�/+/ۖ����YC���E�w@�-"�*D��IǍ�і�>����6���qc7���Y���}�	�m��9���)���(D�5T��ܿ��6(�sT.�yB���ΩjY��~���#ƙ��Wp_5Yb��O��x�bL�������m�v7y)�; -�E���t��=��bEE{hi�
�]hDl�c%@��
D��1p��>����;cđ�M}��H}��'OL��~���AtGp���. ��w��{�\���)��(�b�����X���t<�������4��uF���%{�M�4�4}���>�M�:I +my��L�w_]g���f(,���ݏ�KNNb4�B��zg�a	���[�KS�/�)�
,����h��o�S�����������:w�Z�Y�ET3�n�YKl@!ˇ9��/)Z�gݺ9��\���E[�����:���"B81��AS�H�CN�vD��V��gsKqN�Rȋýge�:2��N�_����9�H�*4����Zc��$���$�69[�^h��÷a(�>�dN����O�!��"�g�a�+n�,Zn$�e_Vۦ^�v�A'�o��i��_�[z]�Tq�|�O����.U�~��z���e"��-w�}E�q*�'�J�_��2Rl�ðq�B��GU�sΒ|�$���
�a�(���iU����e���A�,�L��/<��c��ayJ"��J��/3Н�i�3T��]��8ǘ1LF��]�w��3'�H����PA�@"�ɬ���51�'֥TX:v%Kq=��ڵ-�B���$;l��&U1&�2�qx�������M���"=.���p*.]�	�bw
�$�jċڧ���<%7UqtB�;��»�@�R�츽-;KQ5T�hw1��VIy�8�-�c(F��_��2H:�Ŧ¸��dp�l�$�7"�I�W���/�d�-���^wc	(���ަ�1�n-A�^���A���o��f��!9omKC0�ӆ/�a���.F3UC���\�U���i�)ͧf�U�\�iZ����I�g�p�]��Lݼ;.����ʣ�T1�������	����4�� ��!���z�9�%�5��0/$�R*Y#-�e�����F4�BP}s��~�?5jԾ��5Y�U��M�LuOdl�&�a�*��x��O���T�:m[��j�~�J�e(=K��g�i�\P���h��z��g�d&�s�&U��hH޽E���?yaQ��P���[q�-��� (ǜ�?�������n��XzME�{u�J�ؠI9��1	�����D��>���Ɏ��NB�N-�0c��x���ƒc6�*���| ���j� w������n-P6�G���
ɣ�O��8�ml�a@i��Q����ī���^B/�)�9YG[Ǹ�;Y2��m^�ɦ�'Ҫ݃�N@ �TV�l'�'"2C��uM�Y :�m�<����3���sQӂ�r�C�<�q1�`o���0l�5��{�k�VFJ��b(�5�����[�yy��< \)�v/��'�pLǆkiDnҙ���ܳ��(j� U�ޒݓ��&��jS�q�T0�<&��nq{��΋�Ĕ��W�B���e�L/F}���,	2�Xk��v���������L�9Uw"��Δ��n�J���.g��b}�|H@X�B�Nُ&����(�u���-���;�hB��iZ�9������⥖l�/`�GU������v�����e!s��*��H�H��/Fsr����T'EF0 �*�j�;���Q^qO��ф
��ײ�"6���{�K�§���������WxA�"je ,O��Ս8q����|N3�I|1�s��l�o�2�|���v����;Ыb+];�n���;��®�;�
tl���9����{u�j{s��\�397�004�p���:#r-+6{/�ŌL]V��!�^_��Q��m~���:\�2jpR�{��Qo��L[�i; ���u�@�0�g��=�.hF�?ba����P��CuQ�.J�������g�%H�yM�@��:ř��o�/!md�p8)Q�������*3�/%��yۤh!�s�y%�/���y;sNB�㬉�<`�W���-%����� �y��F�+���z�G����@�Yo"i	�.�����
Ԕ��S$�<����/";.�rކo���ګ�{j�X�Y�1)�J���g���(��+�洭�u�'b�:L#��X������Q|��h)ë�9��Ԫ��2/,K�;Կ-H��/���%px�J����w�5��:K��'W��&��X���N��g�	������N�����):)�褫d�F ��<ɸ���`�AKE&��:ܗNNm	o��}����������.���k���r�W�R��������p�A����$�p�.��\f�Z�r��|D�w�(��'����4Ru.#5�;ʤ�Y�O�|Ǌ�:n��z+��ͅ��#��]�;G�]���Q<�qɺ3㷘��a�쥕�=łt�2����?�mݝ�	y�QZ�oa�7��7!=SB�{Y�6�]��1�N��h��ӂ���dj�s�2�,F|f��ݐq��:.�~/��z�����VP�ʹ�:#�M�_�Iu�D3�4�����3�(��:D�n��f�n��)f��!��e
�����Qǯ�-���`���8jf�50����d��t�I8�b����(����ʥ9�P�)mݮ���o9��:25�P��xT����Lk�7�nÕ��`P����'�.MOs�
y���0���P���R_H1�HD������w��^�Bby�=C�����"偒���"Zշ-�����Hsu��I�@I�/$~�PV��sؠ��m ;�B�~N�W�s/^�I�����c܊���ͥT�%E�{�ݓ�	K������.m$����+�D�%ԝ�7p�(�����e*TAG�%T�B�,Q��K��ė*��>��R=��Mä�z��p}�Uw���pk��6oi!o6���t0*|�0����72�v˻P�豑��qd
)���:w�A6�Ie8
�	��d��W�?j�&DC��=���S�D	��(6��X�����̱D�,t^IM�@�&�sq�4m]vn�$q���3��>-����%��0ﺕ(<94X
Cqؚ�*^[4�1B��?_���(�,���{��Hɮ!�`�)N [�}:�o9(�~�丨�f���j���;l\sN��Ŝ�'wʍd]�utRG��W�@e�&jw��� �o�Ȓ�p�\E(��C$���X0�%���k�.(\-�°#�d�Z��W�D��L%���|p�rH�V�׺@z�9��IC=��q��R�9ւ'�w�gC� ˢ��kϱ#4��Ӏw���R	9 ���AsK��8��~��p"��^�r~��&�G�����J*�y����c�biِ�.��6.zՀl�9���L}S��zGvG��f���㨨Y=���)�=8P;Tҳi��������f��Hk�R�#<��.��8�~;+�ь{�XdC��E�bV�I��2���=���^~�E��[`�q�.�G{��Nr�>Ms7a�6�Y�=���4Ur�f�Qn<�h>��`�!������!#�92��VI�>��u�*'�_/D��m�����A`�f
����5a���힡4cƫ�0e��;-�y��{?�B�8�҉���x2��.@�\{�������~�g������>w���\�k�9\F~�E'B�:6����T�_&d*�sZ�p�t��C
����M��!?))�;���}M��	���/�Mw����ٗwiѼ��[�1Ka�6�C����{7��ן�ߧ����>ZIH[jp|�x����p�E����ҳ,�C0wh���'�c{>}Ȼ���������m����"�sE��&��R�q@�8� �gԖ]b��+����U�x�mu��K[G	0���1�A
G��"�dA)>м^��&��Rb��(�ҭ�#l�Ad8qe�j���c����='�%�h>
�y�J�5��@�f#��̡��/m��WΏ5��ug�.�o�UC��Bԉp������Yz�Y��c�/JU�����r�u�Z�����>���x7���X��ŏ��qW��P��3��E#�4���0^g8Ҏ��Ҽct��Ls�E�)�h,��j���ewe�'>�=���?���w%�*�C�'�x%ځ{�ۛ�b̧?�b��X�DV(,����<S��zW�i�46�0�M\��o��D�>�e��33�����o�y��e2�f�W�����R���q�鐎!���M�^e:wWV,�l}{�w&������գc�{�aJ�{���VH� �)0�繯�`O��_4zNZI�?N'иi ��� Z�����!>�ɰ���:L�M������ûs�x���2�����<�1��"?�C_+�"�2\���Ow�-ǹ�0��̡���0E�V[@��ǘ��ߓ5�)�|!��У���&YT�@�X�%�-��-��d/o�*lx϶p@k�l*�e��/o �Xo���B|0w&>X�Ğ��y�b�0�#	X�����v���G�NM k�i@Й�QI֘�X�O����
��4�Qݍ�\����S�x%~"2 �C��U/�<b�Rǥ-�/�7����_%{ջjX~��3'މ��*>���/���%��mg���k'|3�k��d��(qs�H��T��縨d�e��&���T S*�����6E����j�/�� ]���������?��N-���Ŏ����-&n@�U.)4ShI�w���Q�D�+O@��
���6lQk�;y?�r�QCn�ܾ�*�����ȶE*��=�߹d�t�m������$�Ћ�G��+��x��(M��8���]�Ǯ�)E����Q�Gح��#@��_2����yY�}�RL�7x��,��q��I�yH^_z�iA�eJ�e��L���D�������>��oK^�X�Y�"\x�I�5�glEwe�ͅ��)B�]U3g�%�B:s#���|���e %,����vձ�p;�0 �T�y��@EU?������3)v��V��4�C�V�@�L�	��7�I~����奬އV��ND���fe�$
��Id��M6��[v{�2]�eH=����e�L�:a"�e��qQ)p�7
卫�>����/1��1V�Ά�Z���)�ÿ?N���k�ȶ�.$S���+�i�=|�rʜ�N��ܑ�X���f��%�O�'�y���D��e�
�c�2A�E�Ih���Rs��lM�"�����RsE�!*`Lվُ"+�����c"���aA2��==�q/����U��2n�\�{U��9?�q;�����V��������ʊ���9w�_v������ʒ�~
���{�oi�?�F�z88�E҆�	� ��q�4n�36�q�h�`�10�.?��L+����~/7M����@DD��A�����Cs�KY/����2u��@��V��'����8��J����l��"=��h,��JG��#�hȂ��/�ؖAM4�a�#�#��j�(��D9RM ��1I��$�.���1�Q?M؟^$�����o"#p~���p����u��!i$K�X�O!�RX*�=�'.�)�R��#��;84�L��`�۷x��^XaSH�Ta���DT7٭Ӧ� ItD[�~�fagط�����K+5P�e��R�-�=a<���Q�D�$��	��
kl��v?y�����y�SZ�ea�;���-�ha�v��.�x����G�#�-�4�`��y��J�n0�o�H�Ⱥ+jD���[��5��(����cc�A={A���:���HKD<N8�IͿ�,�c
�L��|!;9�����C2_i3k׵u�L�B�ք�NIe]۝�2�KYk�K!�+���7��^߆b'Y����tCfdA�!9����� C��=�	i����joGp{n���<�#��솣(Z��w�a|:`���k�~�5���%���j�Q�hn�b�mD���d����DF�f�bD���>�>����`��6�2�>��!) �Aݏ�����~J�zV37>0�4�DnyOV��<�6q0��观^l=�3��v�Md�����(�f��D��<^��pi9��Lj�w�	O_��?�}��y-�^%p�ڋT���H�G�������}�q��a7���`�NH���_��
f M��Հ&|����b�p����+}6���]Z�m�,3t�{���9��&�0��ɂ1��D.� �H���`<'�N������U�Xd����s~Ặ�2�C�� egJ/),EI��.�l.4���"9��FH	����Q�=�<�
qY��H�ߩ��<���[ۭ�kW�R�o�I�r���E�������F��k���=�q���t���0��	��7��#�#�f��x`���_
��([M��ss 0�=3����q/�;;Z��~.�� XU�|Ax�?]�G�塹��f�w2�0��ć ���A�(�&h�9�H>�x�>m�JMT1���޸vM�gH�`�J����?���BY<K�ё���ĴIÜ�m��;z���泏}L\��SI�]�Ď��FD�����o?���Ə!H^i��'�^#��=�\�����V���t��V��t���*ZH���*����*e7���e0���˴�r�?z�]��!��D��Mz��V�*��<N�^�4�9Tƥ�O.aR
��*�A�hI� �=,
#� �r������m�h�n����6Hi�����w�7��|��Ț�oonn�<�E�������z�^x��-Ýek{3��޽령Rn)K��(C�Z3��N}�u���q���_ļ���2˅�L*���b�x?�̬��#�1x�z
ű�F���b��g^}ɈZ���Q�{1��Q�ⳮ�9����N؊����Q�	GG������#���%ƿ��~���[��$��p����
�09��l���A�1m�y�o@�Y��������"����;_�-e�KL���1>��ړ� `���Z�v';F������7�����kV�A��9��PdR���`�Am��ɲNN6�Nn�����Ci�L�k�a�=t�Ui����w��=�����T�֖�-lQ %���L���A��|��Kq%r	�g�sr�NB>����K�I�DSɠ'A2��/l�w���v�6�8}�y�Fy4//O�Vw}pp��Gy�k��i	EWG�����`�F۟c_�`V�54p���`8�����8����J�'V	�E�������{��@��`䜩>�=��>�Op�\WEY��qሻ�cV�z��a��~Ŭ�2��"~[p����J]�"����x�dZ�<~��Q�o!��#��f/�,�R�҉DU�,�9*)+k�s��l�p8�>���p<�������:�杔ɗB�L%���/���!-�x-����R	."9��}}?w�NK�Q.\�����䇬���j���\�����
|�E�F����脪f��2�/��W�X����5��.=_F���c� i�=���64��٩/0ht�1�������8Y�w�ߧ����
7��z��}[F�z:�C�Ο9Ӌ\"�]~��-n��,q��fgeg���<��ݚ�X��ny��gч��蟞�=qB/vGttt�c?��0�A8q�SN^�W�}��+�KVVV~o����g��}|����zj09�Y͈L ��T��<)n���׼�u��C�>��yk������uf�`j i|a��tt?��`煍����+++�h D
_���s���G�LM�������*'2MQ�����Q���&D�=��J�9���'�Ffgee�w�V�9X���>��h����4m("藰+J^�|G�L�e�P�'�_����eP�[�U5ǚh�O���W�ÿ�,����u䘋�t���&k�ȃ�� ʖ��j��/~a8~�/V�����?HJ����M3:�|�� �����lL�Dΐ��s�?i����B�����_�ߢR�`a��2�A�v¤�b�U��V]��zig�qI�n��u]
GU���s��j�ɑ���8e��3m��u��*`�Ƕ*}f�ۛ���ɕn:d�|����9��Cr���1Z�ϟ�9��9�&d��2��7W�k�����Nt@�*��Q"���p``�/t����RcS��&��C��`�B2�d����G/.my^P�����`©����쯥�p�Z�
�R�=&zIkruPgO��֦c��H�B�����d��lȉZ+����П5�	E��rY �>��/w&B��
��� Ͻ��a1�l��S�r����	��g��W=KK^�t�DC'�����/_�{�^�Vk�J9��zȌ[�⒙P�D���v��W���x�Ģv2�k����R��;�!% �nX�Ӥ�/��_�τM��M~���mt�T]<^swy$���p�e���>�2h�.�?��j�����._:���L���^��
��bu�;lY~�������*lpM�>����\���+SI.��72{&���r��4U��+l���>�M!��.���w~m�VU�H���HHpb�e�?3�溇�,n<H�Z�����L$+��q��_����Ҳ ^a}o���H}�.�+E�_C�oY
�B���P�BavC��Wk���s���UNٯ��I����_`(�h�i z������7&:��V`w@���do�H�����慨¯�3�x�#�J�v-\��4�M��oi�Ǯ0������t�[ղ����Ė9�*Şw�{%����u����gWݩ{����Y�|BR�b����"�._I������gϞ�6\UVV�績�����[�B���������`a�Zn~�Ⱥ�a1Jf?VՍ$�]�� ����nXM��tｻ�>}b���7�H�0�k��H7i[�� o��7�2�OJ�-M���O"��o6�JO�l���S��B��TH:>KM�e��z˰�"��'0+��g�u�㷡P1`��m����k�[���B|Ѕ4��O�n�"��j� � v�����.@��7e⽓�Zi� �J���jwru΀��=���aȍ?I�\kn^�g�X���g�ee�K�w�hW=Jg菒B�Q��ل����M̉��&��{�_�����{_�*�:��TU�G��:}�g�I�n;�ߴ?W@����n�YC
&~z�a�^��:g�#�[r�/@���q^{k?E�͊�M��|��n'��^�%rU^]ũ(��t���`w�z�����n>�O�5(��@�����5�:��w�#�"5��C����L��la���-j�&3�[ FA��X+U�)�s=�*6��`�%8И��U����7�J�VΨ�}K�L��;��4s`S��@�T��y���j�@κ���yU��8qv��
�S,`��+�)�J���>�t�k�+�9����v!��SRRR���x�ۧm�s��g��6r�k���h�`��[[[S�q���N���S������}O�Be#HZ1ۜ����@ྡྷ��e{;���C��1���/�����G~��|�?�\�����8�c�̳� ���747;�S(Y$8W}\�1򐼱M���Tf�MM�н���?#3�y�4-��ׯ__P��*��s������r(���������@�Bc䪩�*����� o���9��@���5b��.��1I�Z1-Wr��'��-��Ϡ������s���QC�*�Y��UG�&�a�	N����N�y��U�Ï�{��Y<ӒY�?xz��7��S����p�Tt�����@:�k�`7+Jn`�J�a�W7W�c=�U9iͣ9́Y������{�p�C>�7���`�B!����6���X��̮��!�_���I��1���������8�8;k`���a ����m���Z*�GG��b[[�m��������|��w��SO���� �9"�FLG����s*�o�����k���GH�S�sw�x<���&3:��SY��zj���@
R�b��4ȧ�-�[��bT�Y	*����o1t���@X���=UH~�k5G��^��m��� �Z��s��\s��"q�Q
/��݁����;M��bʁ$��;�KG��|����&l)��啕������;��w���c4��nQ�r=�� �a�w����TǴ��A�"fe-��Ao�������oA���<��T|j^��W����D�x�7)��i�Z�2�>i�%?㪾�~���bm2�H'-w���V�(_wj�9���]�ozNk�~���u'\6�-1p)>�K�`b-P�j�P6$=F�=�V�/��}��ԞZ���ϟ�h�S|�~��3�:�����rR�6
8��;rqs�����{gX���G9* hm�����v��BP@Ab���ޱ���f���L!�tf�	��s#�P�x^]4�n�����+gd��g�Z_��v�K�Ә@�k�;��C�ڣ�㴳�3��tO%r6�P���xk���qq"|�1N��|����/���Z)��+ŕ_�Q�Im3bK���\Yed��L6�y�!������|�7�\)�(����nG�L�}XS!�EDFTX��R����)v;gd�_�<�������nzv6e�,�@r{d>�譓g�^] �l��(.��SI`j�����e���4���7>�8O�x�?[W��g�猩�.�h�dw���O9�ŋ�<�ܡu����x^oՌ�^��[,�e�����0#�:)imu�Hў��tB�����8�Wq�JN=:%���x��K3&��r5�6�N�R��:�s�Sp���Q��L\΅����5������wl���w3rG��6(c��W�Ő��Ҡ��*�f��6w��u�b�٠KQs�:t��.m�&�Z.+N���t"�n7��ߏ=���e���L���?���1?KI�~��O /T(���qž���ԻSR��-��7����u�=>��ΈP��G�ֹ ��L����M��S�Ug������G�&�s�,��p�x��^k�@ħe3��9�yy�#��T�4�R@Eg ݞ�ǳ��P���.��i	���$��$dFH~����s�Ң�������O����ƾ��:��0����,ZY�N��ܝ�f�p,v��]Z_�rT���
�~���?̤��F~�٣�H �����2g��bc������5���c�E�g#fL�3��6���PE->�r� �*0��3b��]����J.�����-���<-9��C�ogtg�C!1����+uoQ[̐&#�f·�B�0��j��� %�6��PǈcJS�t�ڇ.��g���U�Ote�/_0[L�YY���ba���λ����U^�_�Z=�w�!P�vB��GϨ�N�=�� h�k����퇀���,$��ܤ$p ������9b�5��k��i�a�ȑ��ܝg<!�;W�X�\P�࠸����K:a�`j���Dd�B�d�G�w@�ƶ	݈��f�����3���Q���Կ�˽��6:��V��@P�O��O�&%<��g��?{�����'�o͍�+u��}���S6e��
����n>EN]&���QŠL�9�I�YaU��75Ey��ϗ�����{�7��2��㓔��%���O��$���Г��	k&f�ӵ���Q��H��;u0�*/[���Zx�5"�J�G�\
��;lr��@����8u R�TR؀Ϛa ���Ѭl#��Ġ+�A�����8�8���1]:�CRb'^;%�$�W=?��mPJ!9MM;\\R"�m��x�tS�Ё���=��;���{Bq���M��!%�1*�n%b끹zyL�k�kr2�?"�����.��d�U���$��`�q��I�+a�w���.{Ѱc~�M���b�?5̧#Q��̾G�oke�C-:�X� 2Uo <�$��$z\�C�����D9C�J���X�AR92{�R����ѡ�9"�7	�H�'�8���T���I,�r�������:w�"���L/��q��s~�� �sv���D//���Ass����5g��JY�AZ���QU�/.yo�Z�w���&o}�.H��W�	��(�`��:j�84��
zh�������~�v���ڒk�kd¸!!R�n�|�����HVeb��6����᤯41���9Z�n��hzbj����ֵ��=�B��˓P�E�~wK2Hv�;K�2�Ν;����Y�L�*hp̺6�!�3��?����w6X	I:::�[.�R�rJ����[U�`�F(G�l�P)��p�v�zn��	�z0d�g[V���>hf���چ�;`����D�}����|�,���?L��y ���	�=� w���P#O��yQl!��Ri4���f3�n0���7�RZ����x׭j�$FVǖ�"���Ƹ.�%L�>@�_j���L�m���޸���<���_�b<�����m�������~�CW���o�o̴�x/ڒ8t�ژ��y�ڿ�YRR��^)���t�͑B2��z~S$d�ſ�IheL<��͗N��;G[|6��Y�8`~�E)Dxccc��`�����W� �aP����<u][s��%7 ��IW�k��t�� ʷˣ+mX�@)�X2����}�G
tX�����B�(@R,!N��7��9
�Sx),��
��
�����G���p\�re�-����ij )���^�w���3%$���� �{m��~∣��_e��Z�ּ��t����_�#u+(3Oz�6���r��M@RC�t��}�3 �k׀��}�o�)%�`7�{�f2�@B|Lb�N����+���d@L��u�J Z�����H8ܭ�}L@}��`y{��]ףj�u�Ha��w�����B�	�j���ڵ�Z�;�c��٦`��O���R.Z��D�E&ޖ�6�:�%��͜��1�_6)�n[�7�A��Q����t���I�.���?�}c�.����%'�^�-U`L�.���2\ ���um�m�][��j���|I<���)����У��v�u�F>�W�){A�{�X	 M���f4	bȹ�����v�'>���؍�� >k6�w>d�H5ǚ���z`̪�LR�[�uSyyy{�x>t6� ��4��tE����[u��х�,uEbm���D���а���.�I�y��iruz\*t���[gee]3<�����fg�X�����Ii�ZqS�P���O<���A䵁]F���lN���dm�V��1�����AT(� �W?���=V�̗���Lr���Y��&�3���~߫�R���]�֐'�i�f_. �L��9�1%k�����WE�)���umdWN|�!wz�C�B<F�f�4��y�ھ�~S�l9L2�J�&���Wa�RT�X+�Q2p�T��q�o<@;f�X��+�cR�C��C��" [ؗ�VF�@�)���.�h��$I�r0�*Ր�#ץ��m�I����]?�#]F���:e�2�>�G�,a������w*.�,�lVY?�yXl��I��A�r���*7��L�%����<�*JJ��:*-�2�5&��jdzU���jO����33����gö�$[i\@@DԪ�����a�zVo2�~C$P'yxhBڥ�|�e�$���g��K�z�g�xi���_ _�3�T����rg�jE�WPaT�N��%$%!G���O���J��贿�"�wK��nH$,j�W4-i�Xʋao7tS�ww����O��_n�\�~��R�=�������[~e:�Z� 
�	u�����?L<f��V�I� ��y�V�ؐl�ȥ�:r�z�J]Ʋ�?�V|h#.X�L�����*cf�@Ĝ5���z@@`��������$a�=�K��O����^d]еY%�,�!Ց��`��?�-���k�cÞ]�H�p��4Q�MM�6W����a5=Ыe���ސl&�lhmݔ��w�%[�p��u�)Ӣ��2V�H�c&�v����u��06p�����um���!���@�&�|�y�bZ���x����s�+�җ��
זoh�{��f����^�аu�n݃@�\p�/��%n�>z4}�n~h[��Ͼ�j��a'[���\�%75�Ng��юYO$�`ۏ�	��$��2�)�F� �����\Ⱥ6o���l�����Z���*Q�zSӪfn^> gt�j��5mh+�t�e��hր�rؗTu!ҳ�VX�ݺ����H�v_�C<(d����-I�z������Pb1�i�wD�w���k{���)
�HLJ�oooO�ص('p�����5������݇$CK�v���܀�`$���SO���zx�f�i��\G��Kg��*�e2���4_]�B�ބ��V �߉�xJr�Xj���1G¡��� �_ޟ6k-e�iw�?0A�1������V�<� X�27�.��,��5���^��i��{�R
�-ҳ�]��}�H\	�E���!�g$�����;R���)��E_�迄5��oJc�ϖ� gJjA6T4e�����wU��n�Og��ʾ��8
H.�k�%�Tx���������{i�_}\[PSG.8�ibe"1�2�f�L%��A����`)H��%T1H�S�1�!� �(�$r��J����#��B`����n��I���y�Ӟ������'��u/X�k�jbgQHA�/{�;�����?k��·kt��GQte��b�o�j��u���m���h��p�J�.ݰF7�n�=�+Dt-,z�����Գ�Q��ϋ��<B�M�'��0��t�9Y�[�' �F���r�ɿ=��V�����~¥B�r��"u��6����%�p���x�4[�0Mۄ����F�7����B�_��G�dx!���īZG&l�A>(�5�DB��� 0t?�\�ݬ�e�_c�' "�� ��f�B�;]L���ڜ!gr���9�]{j�R_8qHHHD&L�!��FV0lf��G��ܸ+P�)E������nvE/�w�v�f+?Y�9�Qs�$O�|8�i�Qx�m,�U�����ϗ%�;�������@����N'�Sͪ��&㈮z��7�	�?�S/��1��_L�4�|�L�:%���'�ʇ�m����������$�l�\��D���.)|Mܠ��C���َw �{�y���h@��'�ۯ,KV�W�ZW�������xR��~�1���� ��2`Z%@�kX��Sخ	�V�P	���:�޾�}w��9�ьA���Bp��	Ϧ ���Qg	�KsZ��T�\�V$�-����nQ�~,&wF�rJӻ�p�䋐ƐK��Xn�k>=k���7�UGWvT��{�3��BT�*'��}�؅�Sw�߽$>_�o7����������8b%ؽ��>�][]�z���2� Tu(
\ݖb�tZ�ݾx}Y���x�T��K��V'Gmu�@ݥ�{�Auʹ�_�<�3�9�!��p�a�t�V�)v~��W�������[u�C���[�T���j���!��NA��կ�>�w��Ĳe2{���Fظ���c���PP�����k�+�܃m����C_�7�a��v�Zss�;U[��N��S�)����`���HR#0S��;Qv��U��of��C�f�jS��q[o�3W�Z�O�A{��y0lPA�q���j�����9��ּ����Tl�`�GMx3)�"�	�L���DՆ�3�7��^�n	<�CUF��Ff����G��-�w�`A�Y� ���*�D�y6d�N?й6O�T�g���\�o?�QbS����.V@����Z�o>�����<z�ǣ��fs�Q�e��lAϗyr�F"-p�qUTA�T�;z6��!+��^E�٥"�U�x�	mIq� i��Is����.~��Ħ��`)��u���'d�d�H�|�git�Fbh���"��t�?���b`�	�A!��5�~Ĩx��|���f�L�Υ@%���P�aq�D�0�=eB���2���8������QSc����d��b'W=d�Z��x"#�y5���PK   �X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   '�X����q  �%     jsons/user_defined.json�Y�n�H�A� 35����&V� ���``�}q��I)��|���~�)ٲD�Me��!��b�N������2LϦ�&���2��lzꦨJ��3�8Ӭ�vi3=�����;{���������U���ϰd�/��̷x׳i�a�r��2�R�}J ���i���T�˪����2�|�;[�����<4�.����;W/
ǒ�u�(g�#�Eˀ��B�	6"[�7p_�r{��	b�D!�"F��iun���n�Mx[��o�/���gݧ W�E������˴\�΋f���ϫ�qJ �X�v�>T��5�-�@l��.�?��T��qU`�N��j������"3 %j��Ļ]S4���SU���[�<�7�+6�:;O�����.�'��x7ħ	|��?��1����?
�����r<�	x=��o�������J��G����$�Q#�G0)���0�R�%Ԍd %�R&̐�Y��-�HL�H�))1�g*I1�����Ofy������d�'���b�Ofy�K�J��'�<9M�l���>����50\�h���I�k`8Ii����rǆs����h�3���y���c9&���,�;�#��0~��
�����	K22>$�@	��f���ȟ�9�d���0��ѫ7P�����r3��5�_�T]-C�*��ub���-�DL�/�������{�q��W����sQ݇��z����'�$$�QC�����Q�ϣ�6"u���p`��V2���e;�x���3���y��n���8BE�����8�3%�ҧ�#�s��)P�����y��z�\�&?�0�<1"[#��<�ZA'�&��L���yS���_w6�>����Og\-��^2$����n��s���Rjð	۴9:���>y޾��M.�	<��Ǜ:��D�w$��
������"r���`�{L�R�ۼ�!����K�����)�AS�G�G˙f��i�l�7+[�.��ʹ�yg�3����P��5�q�i����?U>$Yr��Z�3�E����-;g�gG
KF�TG�
�0T��.�6uo�;�/B/y�<lU5�G�Mj�.��{g���o�@L�63 .�m��Tݿ/�!�=o�h���ù:������M[�����5���Wue=��;��窧��`�
��+��19�yC���ߏ�w�b�'M(���x7��|�!*��kO��A1r('4���g�us��8Z�.(�9�l�;��O�C[v��G9�\@�l��1CF����Z����oo��L:��,��T�t-�d�:�g�ђ�8�׈��)��!�Y Cx��	��	S�S�s 6?�n��	r��W����m~MѬ���z�lI���N�BH�C�"̃�,��"��i'��6ZH˝�H򶍴��\2Ԣ�u�nK�c��75���H(��Ȳ����؀F�r�yO�\���x�}�*�j�^T�M��҅�>Qp�A���ׁ4m⶯Bݝ��`���w<k[|�D=8�����/�E���N�pPu��:=��N�l�뎺ߴ�gs�h��|�tߛw����}����ov>����Q��e�����߳$Җ��0&V����,z�Z�����ۢ,~5vn��\hm8:h��T!�	F�i��
���r��<z��9��Pd���Sc��F3n�Ē�������,t�R�~�P\H2�2��3Z9<	��]�@? �ϧh��t�	G0�(ıvH{c~N]0��R�F�)Gr�Eo^��Eo^�f����속�^1�T���%Aib�A�$�>x~ㆍ1�C��)e�"�F�x�\t����a�?�a���ӆ���a#"2��u���ib��В�of����PK
   '�X���@  H�                   cirkitFile.jsonPK
   �Xh��;�� �0 /             m  images/08e4a639-d7b6-43fd-85af-03d86c8bfac2.pngPK
   p�X��
��� � /             e� images/243a459b-a2a2-4803-9716-552aaa3859a0.pngPK
   �X��"�IY eY /             T� images/63ea08ea-b384-44c2-906e-17d581481095.pngPK
   �X ���s� �� /             � images/6c5cc51a-5517-43f0-84ba-83f8b91107c4.pngPK
   �Xd��  �   /             �� images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �X�r�44  /4  /             �� images/863c2d63-52da-45ba-83bb-7a6a6689309e.pngPK
   �X�1.:�  )  /             A images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   �X?S��� 2� /             `< images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   p�X�l����	 ��	 /             D images/9b0fa5df-c9e3-4cc5-abbc-d39b3818cb07.pngPK
   �X	��#u } /             �# images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   ��X�@M��  2�  /             �O% images/a63ead14-3837-408c-8d99-db2ce98ab1ac.pngPK
   �X$�8�l  �  /             ��% images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   ��X�Rr5�  5 /             Q�% images/d5704fd0-3deb-4692-9952-d29401de32f9.pngPK
   �X�GDU7� �� /             Ӕ& images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   '�X����q  �%               Wx) jsons/user_defined.jsonPK      �  �)   